��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U��S
��Q�$�#�̓�tk`����!/����Gʁ��C�����Ez�h�v��a0@����Ù+�*�a�t��w�E�t'�����\��i��V�
H��(�����SǊ�},�gd~�Z��VXR3!q��3s�����6��A�鬁�����V7����ԣ�j��6�n.S���G�ق�����Kq�{"J6d�Ni��QL?�^&���zW4Ao��|\�rn��
��:vഗ��ѷ�<a1�kછ�m����r�IHw����e䟃!���Q�{U@�+D��V�@�SA9�EJ�C/y�Oε�#<�f`����b�S5A�0���*)Dk��B��d��V�ӌ�2��*��,~���Zr��B�}��ᾣ��m�r���S�ɩ������B�6�q�V�u��}rw��6o�#Hj�'.�mZ�,�Y�"|]͕� ճP4�u~�,*
ی7_�E�m���w��E�����7^�+�n�'��WԎ��ii�f�Z/��(xű��Oth�kZ4�,�gUsA��t)�O���Ex٘J�8�"L?k��	�pӶ��Z`DD��e�4����?l������y̙�P�P:J`��3lq��:X�.Y����7�*�Ө<�(ܑ������U��.W|�+�{�e�Ӭ�0�{��D��*JF��n:��D�% ��n���s"�Y�o||B�La���ai�;s�A?�L�g�ZJ�~���OhwҬl��P]�����\(D��Q��<\m�^�F@�k��0;F�����M���Y�l^ �V�y��W�]��`��i|�q����v�g��§*]�y/�e�ڨ�1�j"�����q}9 Bq�2{|1B�%J|�P	N��)Q8��ę���4%(-*�P�A�u]E=ٸc��0Qo���/����3k��s� �yR��k�?'���*��$�̳D�[R�!��e��g��"��G��H�;�U72���Oן)���/Ӱ��|:3Dz���[nv���ե�z$���6�/ſn�k����ij��-g�W���\��H$j>Z|�DD�LB ��p=G��֬"�^YT��$j����������GF�/��-i�^#�a�[~��]��������������A�L����fH�ɶ�7�f���\?ђ�:1_�91/-l)$�ߣ�=B��V1������f�������V �T�Y�%>���9hW�(�m�>@��n��f�D�2_�ӺkZ���	�M(ML�|���3G��%�=$�"��^L��&�Qܚ/��`J�52�@��sԤȷ��t�I��?3(Q�С���|j����T�'�_9넑��=�-Y�����^0�v�)>)>i���b��dYFHW�l�hBz����y���i��mL)(KD��N��}��q=loJ�˵���0ʋ!?���G-�0���]!�����.G�^�r �6�d��qa�+Lz&���{bQ���P-�(�=J��՗��n���X���l��܉ohO.Tps��KC�g�9b�Z���5W�SR���V#��z����m�p��ĉn^�P���l���<gɏ�Qxk|�*_��f �X�٫��ܹ���8��:���O|��Xk�2��Lh}��/�;��R�g1#V�L���~&)�CI�@q���(hVϪr��N����)q�	���/���͞������~�j�3�b��=rC��"���D�������"��Tr���jF3}E���ߦl�Ia��Tv�.�*;+B�f�P��	R��mi��a��g�;�����.��yL�tu�9�w�cn~w$���̋�"���}�ǿЬSG����5���Z|�����N(C�Ń��&F�q`p��@�p�������G�9��Z�O"+w;��S�R0\{Cٚ¾b�
	T��i��m6��!�h�($h3~�r�����4��HT����N-s<��SW����4���� ��'�L,�uN�p�m���_*Z�t�S������^0��u�6�g�d�	BR���l�bH0>G��!>��C�N-���V4��d�:`�>��7�s�%ڎ/�q���º P\�>^��c9.T��E�Z�����Z��	��S����TBmbWC�R%.J���Mb� D��u}���FC���R<�k�����H��������U���?w]����W;8���ږ��$2mp�L�8����G����O��Os��oc��G� �����`7��vS@(q<��?Cx.�Z���rD�Ȓ��PU���(�P�kš;�/��	���P!�;�-�g=Ժ��\Q�pŝ�:6#�{6�\rg���$|F_�����]䭜U̧�����x8/|���)�?�3�L���ZpɾiC�Ox�\Ю;�WNr<��on2z���+�.��q6L�e�����#�%b�c}�7��܇��!Ȗ�R*y��&��;�������/���"q�C}T[A7h�H/�ۮ)�����tC���%)G��i ��e_X��iuMK\��� +��bO�����9N�P�M=��e�GS2���G��z���	���_�vj�+�UE�JE���T�AO��ܞs����X���6�ޥG ��D3�t�>�۝1 𩾸�)MC�1?M�=��UU�l�����}ߴ�ih�C�+�ȗw�.��G�9A�Ty��2
�*'n�[͒�TTe���1�<���7Zx=�u@�''�>z2��i���W�it���"�l8���
�cϳB�D�xl��Ma$�/tH]�1�x��+��<,��R��{u��`�0��)��{O�[C�r*W�����'�s;�t3�2K�WvUY8��-ވ�R�^�qCA�ö��M�i�r4۾\Zŀ�X�K��@����JUR�����
�+�j\(�i2x�v�`_GOK��wiz����g ��3�~Y�����kE"���so�����X�[��ɧ%���/]� �d�}���� ��Z�n�ޥr�
0�P�Hly��r+zGޝçx�D%�@#�
��5��l��S���Ql�=��>�B��7vY���hY�>pًX��7iQ:�J�~|�u��a�z����B|-@��@T׷:C��WXG�wZX����1V��% 2 ��1riH%�R:|�h��x/1��L��)�:ع����������| ��������mP8v�)m�f��%Q��'b��q7\a��Ez�Q�}��:�T����#0� ����Lo4��`�9b+,�UyZR�*c�4�)��f}�7&)�?���{��ݟ�>Μ����-g�-�� ����"��NW��Q9/�g��N��,(���<Ms�Y��y��j(�6F	����|��^�8X8��o|�մ]r��:/|M\6�nY!���5Ja���)��Yi��q"����*:R�B.6|�L������٥/�ܯ�ԁ�p21	)�]��.����G�1h(����v��z����,�B����Q�4���խ?� 뱺�n����Ǔ�9V���8��r+Qa��f�2���9�߇���Uk����\�m��G�D�����sʡ{S�έ���p��4�"�r������c�A�+d��N"�,�(�.��y�y��"�iOp7&Ly1��#�|d�o:�Yͳ�eb���S�"$�Ĥ�.]Mu�Ę�����K,�ؚ�5�e	8�9��]�d�Od �}ʦ�r�[	Ţ�Yx�1���d|���>}��Q��gP^��	�i��$���
pnHcjЋEh�o)׀�u�"C�S�_�K<%r�.{0%���w�-.���n���	W� �-7>�������T��&(#4	�Q��=�"��*"i�P%�;�3����81��X���I$��Ddmnn*M���ӯ� �M�j�"^���.�ׁ59H]�ӟ������d�l԰](m9Fu�?q3NzQ�=Ll7{��^��t-�@�vy~����%�#7�#3Φ�Ӗg�C+���b.u�q�!��(cph	L��0�((ٳ�$��]�[!sp�a4�y�<�|�hN�M?����� ���5���is7 ��$��[xs�(g����a&�B+7/ �K!���U6z�L�?�X܅:���S�uwkҳCc��sO�LUy9:y�N��+���d�*��=n$�sT�����j��=o�U�E��H!��*�Lԃn�Ě#8��5�7YX[_�����nylAE�A�u4�7J���o�bǼ��UX�|!N_5N���z����rLv�_x�$�,��>n����E��{���B!�+9����B�8_Ǫ`�1_K�	�B�Aju�ա�Im�J�j��ke���[�C��B�f%nָ0N�R�	C1x�:!ճ3��e0Q����^��fg���	��Ӑ�T�WW�\Ш���ol��1� xp��A� ����^HDH�D���xbM�>{��d��_\c}��tϙ��g&��]<{�N��A��y���-�Z6`���r�BG��`�'9�
�V)�|Vj���x���	U��.���B��=Ҕ�Bgg�8f2j�ǃ� ��Wb��a���A1u��Y�� j��L��Wu��}x��u�}��2�&�KC�֛�#��aW�A�n!D�A+e��r�;}�v#��E>J�l>&:��γ��#��i�W�߳�ׄ풘�3ݭZ�`��֦4QT���2���	��i~ڪE;i�Q�xنy�R��K�fn�E�,�/�	�8��z�i�(�"Kb���5A��h�W�b]&��Z=$TD�{�&��U�� Ҏ�bi$���V ���X�(zxg�# ���>9!{n1_̈́;w�ݷ�["���娱�3y�L~���2m(ɠ�rf��� �nsX�	��7BySv�-:�z��;W� �q�H��6��
�xh(�b�d�h����n�g ���g�[:n� ����T��f�� �b̪2�A�G/���?9k2���G�p�6�m�<iV%Q3� �Xa������ QC\��f'��D��p����Z.���h���)�6#�V���2�@)�4;�>Q�G���Dq[2�/�qw��y��Pp�Yo�>�@��P#-¡pk_���_��LX���:�{��c�=��	�0/�p����2��]|��dpTg��j�Q���|$��.����N1���v]����)�	vL�p�n�I�I���i^�bT��t�d��{\�&��9�'�wA��uq*���C�E)_�Ϩ��♜�p�+0�Zg���f'P˖GvBq���rNC?~�M�����<�������av ��+����W����)��M �ÈRI�PA0��/Մ�s'QG��Dy����
R�,˽�2TB��yQ��b�E� %�H^��:ћ�@���ǝ.��X	j�,�`��^�	�֍`�E�d�c�2��l�?��m��z9w0(�0�_����<�U����9#�?P,��[���[��ը�'���0�3&=u��o#:B���"s>��۟iF���I��ܾAO���`N��1���j����y
;��V}���2��A�+/*	�]�6i��N� u_RFSr��h��y!���##J����˶�j��Z{�Zi62DɗD�o���U���p��P�흧�%xiI˴��n�1GΈ+�Պ�.�s���16�a6�Wjb�j���<˵��õ��s:�����pM��s������W��s�R���C�_B�C�x���]�!�r�=�]�,�]�,�B���m��^�<�{]8/{��c���ί����#��kke����O����K4'N[-�Hk��L�����i�O��8���|�Ё���SK��Y�O�||if�(�[��
a��_b�'HA+�Ԋ�'?^���R%��o��V�bɃ���"�/| �T�Ԥ��oԣ�f�E'g�����8h�mg~��2ʒ�Ԅo����؜q�+�Z�E[�mV>����C�P�����)�`fP��Ƿ:�&�8��D�n�+ ����8�-0"|������+��(!��> �����V��z�F�P�3�!-�S��+�cI�9�����t����_�Z˟VMX�V���'�]F�I;K�^Yn>2`��R6C4�Pmv?���M���3��[b��G_(���{#�?a�eQw�p"�i�b������p���fX#C���V��&��YZ۴�*�K^���IHm��} ���J��<�.A�t�����=����k�8�5|�t�b& z�D�A��$9����ӱ`eo`ʖ�v{$����=���N��/"���mH�T�3�0v}�Xo �-=_�f39<w���gMv������FmX*�h�X�H'.� �b��lǋ	����TKߏ�����/�%�ִ�����a��ʻk7�q�����Q�l��A)��V��&�*a��Z�C�X��v�������-���%M!b�:��\��j���Q8R�g�j��	5����	��;�f���{�h!~\h�O19�9Yah+G�KK��xpա�tvL7'YėB�n��t���/拙U3HYl+b�űT=+k]�8� �P 0��5;��c�X�n�<�H�w��>o���c0���E��uG85��<!���Q%�MnL-��.�qm�85��D���-��P1�d�G �����X��^\�]s�˪���`��F�N�ۤm����G!lXj�	�2i�X��'����tZ1�1�uE�EǸqt߰�/�
�,G��l�_n�|�e�Zת���8��ϓkH�γD�f�RnSN8iC�_�ό��ɚ�nv.���
.����-��0���+�/�
<D��3W��m���Xq�������'M!�
��-lˈ)G������~W�;�h;�#H�ܓ���DDq��_ DIP]�6��1�G�Nk7�G�O1�s�ٚdL�c_ӂDP��h�j���um�w�ʪ����BnƬ ��d�+��a!�(Ik�U�Eͩ��lI���Ԉ�^~*��K��lќl]dy$�����Q��T`�8n�:CS��\l�{��@���>Oy�;��c��x�\	O��چ�g^۬[�GS�����$��B��>n<�>�TEX��8g�_��y;�P�H�6��s'�*�k#�����b�І�a���&��p=:�_�	��Nu����g_�U�"U���[�d�(��ֹ�9'sl��&�Jb�I�G��1䈰\��ϮZ�<M.$��(�a��Gnrf��M1f�R�#]NYvs��T-���)ԙU���SCX+�&7T�f����Wk_j��i��?Nɝk$ n���퍥����*��ou�`<��J�Z:~ļ�f��*�	�K�9�VS����Q'�/*K3Kb�.?:��&���������>� %�j_*�:�A��d��Ə7�[�����Ǟ�O��b���B9����G�;^sW���B���� ���y��ɸ��h/�<���o�)�C�	��S�iB�Rv�Gp��@�h�O2Y�ҫ�\vYP��$$��i�ɾ����<�y�>�v�bu~��w]�6�ix�����Ƕ����-�i��C��T�A&=	����5�T��=ۜ~(�(C��ժgy��z ����;�\���1�8�B�xd;ћUp���
��tbY2G���j�1m�+�+�_Ӂ�#�Z3q��A�'�Ʋ_��z�~Hs�Y����FR@��
�IMd��"&E�:�u�j��;�/�Ec�)s��0�a�8T"Ij9��R�Q�7V�O�j����V�:�G�Ĝ/�ǘ�7,R�m}hZp?P��:83)D[B'��"L��xw�tȒ�\��tҊ"�pL��
�n0_~�ִ��s��ԋ	�P58N_-��%�8���%�[�5�@l*iQ���s5 �QK]h$ k'��_1��)��l5&�e�+ˇ��>�.�ڮs�5��mN>��U1�a��qʲ�����P��ؿ(s>ӟ����n�-�@�!�Bވz��0���p�_[ߨ��j��b���P�������P����4�\K��N�눷�9	3�/�*{Z���e���@U�[��V�В)��>�u�#�.}��9�Mu/33y�E�|�^��ZZ�c�߳ �4Ŭ�*Ή{�A���ҟ6IoM�����ԏ!�R���-�4(��yӷj��EIu�h�쀞?�to���p�e{}�i�:����%��L����\E�C�B��oAS��Ȓ��W@��˶u\y���s�蔽��_���U	�E��r׀P�W�VG�b�"5D��@���u	�1ر�7Hގ���ʹB���Uj����I@�3������<�?0O��'ؓ�H�1�j�ݱR�J`䌿=5��%C�T �����$c{Ӭ{�t�Bة��J���@p�ۦr=�1��rHV�Q���N�y�A�SU�/��Xr|��lsMK6����k�6`����/d'϶���!�>dxN~]o G�~��W\|�v��-�Z��J`46I���ʢ����ajk��9�%���� V8� UI�y`�9؟fXN��7��y��ze��z�odW0c,�f:ӊ-R���~?�qmɼ���٦u�Lm���Ӊ+��Bw��giyj
{�Q0���pU6�W*���È�}���%���9��G��o�}'��X]'s��W�3R0������1� Z�<;��&M�}1�E�����dXV�iDG-\�%1��t燾���gzF��m��Ozx�́!Dص�&���k�ү%�}{�[�KK�8��B%B����8qcq칪���Ad�f,ΈiԤ~&�����t`���+p�\f{��?��GfL	g���@@2kq���(g+D�'���و�#�J؏����W����#�"^����y��:r6��q��.#-��E�l�EٌH� =�n�`�O�{5�
V�����GJ��"��I(	��+S��GcJU��lRW�t��1��a}��Q�i�Y��	���.��CS�r�C��E�(uU*G�Q9}&Pm�CTx�n����9b�6�š�ڽ�34�S�,.��H1ǔ�l��@L����*���L�&�m<�g�o����*.�I`�9�U�ɠ�\��'���=�].δM��q�W)v���M��Bɶ8�9��� r0�!U5q��<��w��K�^�/���zY���R+L�N�-�M�����	��(��p��8��zUP�h@\�9\�,H��D�A�gL�=o�q��.[>��&�$�/��Y��:m�tr�/#��viQ����XFn!�.�p4��?=LKC��~l�F��4ipY
�k��:�-s�_�ɂ}v��/��e��W��g	ъ��~W�6p��)�(��,>�f>�%$��CW_��`��1W�T�ա Ba��r���g�@~P{�H�������x@��ܴ����`H�0Z��*q X�ڷ^�����w��ƙ� ���^�ehh��q{�p	V��y /���鍌[c�=�ŝb�@�������E���&ӡ2��I�'��|�����M9d��_2�P��QѰ_�6�d�-�>�PXY��}Q�-[:@���Mo=R`��Px[d��f�3��2mh�iS�M�n(S�~#$	P���ZA�O�"�S�'�n%�)�Zʛ�
�Z{����}4��	�U�"�,{���}����x����l���o�k'WQʘ�K{ R����;�Ca"~�R��m��/g/ȑ�08�m�Q�}�B�x�˫��V��k:�{��5�DC_�ØΟq;�A�F��.���H������WMPL9q"��ܬ1�-������O��LO�4��r!���dz�Osl#��[![�7���y�"��˩3�a�-.���b_3L8�v�����Y��Fe����(�p�85��; 5���צAjbA"Ǉ&��^s}�v��xoێH��O|�b$i���%H��I5nc��3=��O�и�-�/tk"tЬO-~�\}�k,��X�:�f��2x�X�獍%s��Ȇ^*�ϵt�Ͳ�������'������F}�^̘��o����*p����A��w�"���cN��z\�&���Y�A�`���-��b��8+��őfz]��m1���f�������Z�? Î��Q].ͷ�N���y$ۄU+*��vF��i��R@��R.��󃹦�j^���"��s��^�3Kt�!��{����z�tB�En��Yd=_�O�V@C���Az\���7gnS���u�����BQ�0͉���C�X�(��^�\��q�Ӝ��V��p�~��`u��)4�X�3�#��\�<�.*;�]'�A�\A:����]�3GNZ�¢���?��E��j��	�b����c�yw85�B��k˼q, 2jz>8�y��vM?8�+����l6.hdUҜ
����D�! V<�7i��s�P!��o ك�B��g�p��bsжy~e?�)��L �'Y�Yy��s�]ψ/lb��Ip�����fQ��d'�>���Dw�p�ix̽�<�bh@� ��uƲMs��>,�!�9�).]h���&qo�b�����Z��Pc(�-��-N6\Ӎ�s�Y�ׅ�@<���e��yF�"@T��8<�O����Z�cG��9ϝs\�g��n��|�ii
�Y�}c~Kd��̘���ޜ�<ׅχV��xO��
��u�>|�g��`*->>@󣳬�_���K2��?��HB�l�Oڀ�݌G��q�0�� *�@���nA��0C(�#+U����e���u�%�C����7��|t��`Z�����#�����t�is��4����q�m�kU�cp�]�"��V9V���&*�QY�
�H
 Pİw��_b@�XhlN�;4�0Y���Wx�ܩ�g�q!�J���z���j�ۆ�Ԩ���	�fR��� �&�M��Z|��Q
P�T��p�8�q��g>�hR&����%�\R�tN=�4"����nq�)#���+�Bd�G��Xe����.�<�o�:/�Q7Dp��T�{P�CuԤ���
�Wvyp⋥s;w'�HG�� ���:����P�r��F��� ��z<H�{�����R�͠��H��Ҭ~�%��L$��¯�nqb�;=���2�ޑ�:MuY� ���ɗ�Vz�\�@7tp�UH�%�g�5������v���=�VhNw!��Ų��oP}	�"�A% !����o��ƛ�Uҳ�1��@!������B ����mvS�(��>#�	��:6����m���q�nZy%�K�0�9U�eץ�fbL/�e�0Q�[�ē'!c=D��	����i�om���XR���D?U��4y�����~fVd��kG��{pr�sN��c;�_̮�N7F{�"����uo��?t{9���#�ݗ�ȌQԛ�4�QM�A�rHCm2�ld�Z�a%�/7��As�過y�Q.ͳ�����щ������\�YԦYJ��i�S˒�e@�>�kN��,U/wW�5=7��������3ΫEۣ%�&��W<���X���ųG	�;89��&���!L����C��2���q��J�|��k	�Է��V��q"��&�*�gZR&�'��]P���B�5�3�I|�R1�Z��=Q'!�``��T�`HFǋ�_�._�f;�:�z<1��[_Hu��tl׃�5M���r6ރwS�cn��+y�g!�>{"���� � �K�Ec|�n2��<͍m)����Lx��EVG�w�DU�r<�ʷ�㨋��~8�HE./�N�@�ʜ�:�i��!�Z�Z=�C�u�<�H# ��n�Y�w88'R�(SXOL��	�� ����!+�`\��-�=iɾ���o#�J9�p?����36���j8k΋����w�-f_lcJ ��4��v�R�����pU�2"� 9<�B�&�w��Pv��L4�xN�S�qk���K�M.GӒ\
)��l�5B7�4:��!�|�Iߓ�d�܉C�\�� Vz�mP�P��{�ї��T��T	�1L3��`C�iG#��+�:��g֨B��We�ʲ��=+r�bJ�@h��w���2j�}�n�A���&s���r[/�)�H��z��^%�j��%w`����g���q5�U���
�}y3� +w� D��qa��\�n����@�(a�{7i*�'OS��e��Z��5��4��5�0�>��<&9��A�<2��2��e��6{��Ⱥ-X����ՠ7`���FT�E�K$ܫ�#
��` y�^���q+���]U�1��y o�l/�`tz}��uj��T�Se~����~����=<���Ʋu�b#��c����d���U�t��)�k�;v?O��*;�����ݻ�M�iގ՟�h<��u)�Ϭ=��	btŖr�_Dv�=��ԙ��F���[��`��E�v��&�*����\\��ft�Ki>��z<�0�LM�v�盛�I����]N@�z��:�<t��0�ʓ�m9ߔ���_QSi�5*1���hS���R����Lf�ڣy^�PU��h��ڍ�-���E�&%߱�=�3�|��T
���Ǒ��t&�0�o�N��_�7���6�+�H�]YPSu�6�F��z����<�ԁ�gԑ����~28����}��y�~�=�SU逤KMF�u�Ѿ���8���J���TGS&�TE����ax�_0�1��*D.٪�qR���̰?s'��aI����M9�j�z�;���8t-c0��
R�}�� �GZ����o��Q��
9�k��f8�Ehc�(R�!�4�E���޷��,Kf	���jՂ��b�S䞝�U�#MG�P�S��wULl�.��*�Y~�9���`��-��˼ �!��@$�Qy.cϐ;��E5����>��96�c�q4"C�QM�Q�@&�UN������)Î%����vݴz�Mv9��2���o��t"�8� ��'ٵ�C�I��]����r/�s,ŏ�	���߫w���º6�9�����s�Iu�l`�w�K��XE�����Gqj����p�=��׾I�y`@��#��{�����vgj�'�˾����*�yx!)if��ţ{s��FW�M�����*�Z@P=&�^��Ƚv��_>D���g<
30��>[(K����=�HD-<B��|��}�P���ۣ��ﶞJ�'�/���zq%���O#�.�J�V�bN�!�ߑ'M�G��u0(8	(b�?���(��1�����x�籗�?\��T�a0�2��*�ﳨ����Qֶw���u��%h�B�P�P~�NQˮ\$��Z��?���7���0_ool��ciQWG,�������.e[�M�0�(+�]r��h�����J�s���
�^�Xڼ�@���^��-��3��s�u��PIl+Ǝ��,��u<�(j��@����x��w�����ll:俬�#����W�E�F�F�H�rK�_ ��T[����K�9�X l�0L��W^��X�$��sd���N�ϖ�DIS��|ٓ��%����p�͗�����]ݡA]��'�x~R}-�b��PN�\������K/E������HѨ�ی��$
����K���4 UƩ��`e�Rb�`��{����v����	1�i.�+N�K��cc�yA_��r��&�:�_H�¨_Nx�~�eb�%��c�t�Ά˿~0��\��V�d�e�D>���H�M��|g�(w�xg�kMǓݕ��(��#���DΡ�~gm����T?�jGgc�Ak�J&����E�Sy�� ���V�b�x��EI x>�!
]�����j�V��%�Cz�2��`������"���iD�⺋:�q{z3���E��A%Ǆ�)�-��oV;m?Jdz��UA���<vު�n$H?�A��kQQ�E�ݢ\�ɚg�"`�7��'�"y5��<"0��[�k���� 5�Q�Y����R���]�1N D@k6�4��>f�5�g�]nDlpn��Q�~����n6��Uא/�Ѻ����;ɿ���B-�=C��D:%�:�g�`�y�մ������ŝ�0f@1<�&�Pg�8� Q[�ϱ�����9������_%G��ު����*YE�)E�"D���S|<$����Z���9)W�&t����2{g�r[T�]�]�N��?�!��xɥ-�(�M��m`�mR]aF�3�*:�N�H>�����{gO�G���"���/��������E7�ݟ��v�6;�6Y�*�'BcYk�A�5�_r(��7�����Z_�I`��ze�={=Y��R����'�L���μ�J�Sei��@�z��W��b�+�h��ȣ�\0�HrH�8�t�f`�Z�~����L��d���$5H�M�A����4\�E��rT�^;H���)8y�V����T��7�w?K~"��L�<�|#��|�TcF�O��}�z������C���x���x�yzݾb�Ȳ��`�=��9{L�n^������ӡu{�r�BLs��%p�x@P>��tj����mQ/[��\����R37	�0`-Y�4����5�˞e\����
7�y��,.V1a����^�|^kr�3�9S��/�چ�z����s3���6q�}Ff�3*c ��B�:��feC]U@�>�D=�b�H�D��Ta���|Ϳ�r�����+��;CW�g??�&r�7n\9x_{�j�n�,}��!0�T�d��ƪwro!�;�Q�К�l*S����b�_��O�	���
_~�A}�1��(���4�ϗ���s��KmU�F�[��ý/%|�l�g.Vi��D���'����&���1�2�ϋU�Voi�SK�"MX ��ׄ��U����Z��_�J���2$�� 6[���� ��b�\����w��M��e�<�����%_yӂ���*�Baɴ�#r4���!=J.:���|�>I�(w|��^�F"J7>TS{n��C�b�(����� �ÌO�T�hk�T����}�>�`�E��	��q�&��-5�0��*d�mZM�٨�r�kwBX�5�o�Ň*tDN��ƒ�����!)e����[�˝�,i��s�L��z��dQ��wp%UEe��ac�p�>pjn�:�T"旟{��9R<y#k:EG�&vl>' D��V�Mtd��g_��� 1t���!�Pw.X�m�8����� V\�?�����4.�P��X�=�	JJ�=Mτ]̾�UT�� ���k�PN������g9YRV��Q$�fC �'q�L����4��2��[%��+�^w��$
�z�(�S��`j����g4^!�7l{�����:h���C�5-��$ޕtN�`I=�nI<�kZ��T�CW���mե5�
v����#t_g�G!�D�Ng� �w�v��t9���%Q%�&��I��@FYK1�;@��,��;�?dh�����n	�yD9��J��2x[����)�K��)$��M�f���}�"6�}؊���>lON�G��z2�E�yJ�]A�Qo�b�;��!nm��da����Rބ�^R��7��I5��7@�C	�y�'n�#j��$�́)�^�/�נ��j}����o��ص�r���ѽ�8v,K�ҧ�����X%!$-#%���b)0��ݐ�ĦM�R�tPpGxw�,.����@��צ���?�)�cn�y�@8mʯ-�]�AMTfV}6-���^2�;��I��n�F�g�s�C��rvn^��90b���z|�f��.�ħ��������7-�S�,������F`��2Yx�WJ�uH9;�����S�0�����P����x�4R�Ҁz�B��88)����t�6��Nt�L|��䚾����_-����@�S�k~x���g���2���MF|l�N��F����V�8�nO+=:�L��s�Ą3\�c���k^��'�ƍ99�n���WђU��O�|L�g�W�	]�N�	��������[�_f?�����Ηn-*�;����ʎ'?޷P\���J
u�_J~��g
0��i��,��;-
w|8�X��U'?��k�3���$;쏀�t��C,G����c7��Ş0c�XI�:�+�]r�qc�2�DK@MKڬ�nm(�y�9#G�@���M7�pn����P��ʩҷ�@�����`�T�FU�$�6ZԘ�<%��O�R�O5�b���k]r�s{Xj��65�K�:�-mU��;ň&f�q�����=���=��T ���%)0�<pq�YT�3���s�	�{;n��Ej���P��j�c���\$TW�FV�n?yl�]u�����>�#���Pm�$�?z���>^�����Λ������� ���-�"z��T�3H�aC�mnt�먻qv�'-E=tXZ�B�$+X��9��!\������?'�2w[��ʍ��K�6�(2u�e�60�N��h�.������2�Ǆ�s"���:���p5���	9eqG��ņ#NG�F��<�Q������PjF�#���8�L��&\����L�|��&9�J��7B�iI�ٜ��'8��3�'�"��e��H�Gq)�e�C���Kt�9�(��ug!f+ݜl�x�ѧAPyd@�l��x��q�S������bS����oS9G<�*Tbi.�w���r6�^����;�"�r���2U=��,�����=ul��X��@�zc�Z$�T>��-v(f�S9�YkG�3�D�/ܬ�ON��v4[�
������b��!\�EQ9u���t�6jMx߷k~;1�N2Z芇�X���
YR��)�p�P��1#z��5�B`���EĞՕ������[��<�V�tڭ��!�<c9�)��u�ь�m�4 ~{�EDN��bŇ"��Q�q�?�e����۷�7���=��p�΁Z�lLi�_��]?V&j�:5f�-2[��~�u
�>�bا.֞!��±+����KM`E}"���~�����1�f\�(���=���C�W���Z�䰐<9��4��L�	�B�0�N��@Y/��wш�i6^��û>�Tx�q�� �Qb�O~���t��
���M?�/�����dLS">��e��ݓP}i���c��CAoY�#��Rcn<un�>1}���x���-v�Ӵ�~(�t���F����T�攫M�Flb+zD��CtP������Wx}fuf�4�����SD����JJ�s+0<�8�B�L�J�T"Ի����o���$ ����D�������{P##B:���t�=��|P��;߅����p��l%����q����T�z�! �"�X�hn��߅��߶ش����S{�FOҔ`{,Y�`�-�F���-�c�mHu�������qi�,�u�*[�����k~�C�*����N�O
���ldu���n#�s�Ê��HJ�,�ֻ��i�L�R|����w����%�=����ɫ�c)�j����t�uF��|f�$u�mH��66�p�Sj��'��$��}r#�����a��7W8+T
�?Ӊ&ty��ѧW��MQa�&E�6�Hcn"��(����P�n�b\��6��^��^`Hg7,D�X ���b%}v<Ux9r;�H:�������M�'�/�b$�X�����"!`��	������"�<@�\��F���<<�4`�4�D��Q�W���1{�1e�n���� d?*���H��a���f�c��`�S���?p���C/M�cC&��M�9��1��YY�F�C��&����/�w���ڮf]�˟�kt|"��h�F�ޕql$�{�Re�p4�6W{{ Fʋhd����|3i��7M���oR�gq��`�����E�&��]�m�f�o�$'m�˚ʨZ3
�Yq��n�(��=��&[�&����~J�W}��Q!��`l���Ճ��g���Aj��7��
�jN�'����{E9�F���f�h��� Mk�&=-<�N��u !7���M��������HZ6$��TO�y9�63u*�rZpϮaKƪ�E��� *7��%v�S5�+M:j?ڀdE���ˍ��3$�_���ѡn���y��"�۠�(��/{��@��+�j7T߷�=p����u�34Q�6�o��	���&�u�*C�b��%S.�WHU_*������Cj[u�]��Ư$Nv�/&M��}<5����Vڭ�9�s�uQ:�y��&{ ���ux�_s�Zs\��`��ij4���'�|�/;R��P�+i��$܈�Fed��gUE���'��+��DP��>)�@Լ���ΦՉ!ނ�Ɍ��R�Sa�~'��_$أQ�Ыm��13�Y1�C䁖��z꾖ϭ*&��eޞ�")5�@��L֫{V#<�V��WVkK�MԸ�h<���#��T��;�	�i9n_����G�`s,�t $<�ʇ0A�AH��u�
��py�(���u�����c���ڄ��� ���D�ھ�d�6����'h+��cqDz��F.;�:���m�[qބ��x������6��B�j:~����;�]	H\�-�l�4��~�� ~��ފ����>(rٷLL���ʯ���c�%U��O�)���?�k����*	��z��s��BZ�� ��v��JƷu�����/���m���?BmcC��NYe�kb�$�%�9�n��ր"����\*��Y¼�E����
�ذţk��x�:Nr4]��d��(�eO@�s��A�?&���8���C���_�".�-�y�;�Trҧp����}_��͈�0)�϶؏i+������T|��(>��j&z����桻��$I��mؾ��h�䭴�N�a ���-թp�0NQO7	����1ĭ���#�D�q��Bvm��	`is_r����s�a�#C��O*�
��)�Xֹݧg,A�MJ��f1�Y�l�Ы� ��~~3^Ě�]'���3c/I��9����$�'�q��N �t�ȼ��2���VXz��/�V���_�	�S��h�Dي�a�y
̅�vH0�P���c���Lj������r���ʢ^R�Sw�&��.$0v.�% &[�K7kk��-*�?��g������G���.��O��ՕK��+��8sP |�P̼�3��,�C�z���S��z0��-�	��ㅮA~��u��y5OQR�^r,��3�EܜY{D�̊0�����a���{M�}��\&3���L7���!��c�!	XX'��L8��K��;��2�w}?�YOp:����� D_t�}+y�{�m�o����D�6'��u8�=�",�f��oo��OJM	I��[4bO)L�۠�
X�k&��g=�p�k~����}8q��R�ț/�+���J�����`G+7�a~#��aB�򇂒�Bɟ�B�Qٮ�!cc��)��By�(�5ÌG��HR ��w-�\����j�ƿp�AN��᭲�'%��>��7)�m�+p|aZ��=��Q�z�/�i�Թ[9b���C����Z%���4_�֢b�����v�x�6��E���Vb��+O�$�9��'~(�N��7��	��P�h������k����k�Nq�:U�N��"j��q���i��ʱ��һ�#{�J�<-G���G�Z��t$�v��$p�K��,�c�6���^t��"g�6iQVs)^U*l-90dq�c������|�֡7�J���A�\?姖�(�p��E�kD�hf�Rb9B{~����� �Q&Y7��� _c��,@�q��)�p�a9��!�nMF�%v��l��� N>i	�s�$=(���YCH����ً4!l�`���/�d����H�<X�F}g1r�/��`y�㾡xf��j��
	�y�gA8\17.��s�y'ng����=�Pj��3u�a���h$�1��IAl�������׊Y>O��e��셈���P���Sfg�-ym�0�R�m]LV�?��4Gޱ�˝x�,����uy���*������y>%\g��^�t+���];�hJ/�IU���[�d�Ra���o1���?[���V�v쐆������Ù:�}g5����K�)wfuW�]W�1+>�����]*��9߆�n\���F~&��R���HYܩ�J7�9���ȋ���`��r�R;)�@�)��I�����>�7�����\�Z��M����P�G�#fqi`s��ln��a�G��ڮ,֗��� �<e�\N�������FJj��j��P�BZJ�^�����5.��ĜO��CR�����lR3��5}��߲S�Guv*j=t���I��W���{r�J#��� �����o�߯:�~$$�+G���oY����	jP�ё�w�pH��A;�4�ڕ��G�VeC�<�nSM�Ɯf�ņ�;;�9zk�Թ�V8�{��=��̳xӰ�?xO�¹�̢Y�L�v��!�ha ;��J�$Y/_ln5�L���V��i�"�[
�e�5�90�����<�nh���B�mOOrfS�wFg=�77eM5Q��U���+��Ɉ(w` ǹ������E����h��ˎ�(��<�}��,�f�|��a'�KK4ܬ�7�v��@'�U;��4S���U��{��mB
~��q�+9A����dx��&��B=��Jt�O\�h�e~hx]p��	�<N$�V���q�}+/�Τ
��~��?T*㴴\C�{��v� �N�>�I
�/<c�D,����m1z�HHo�	�n��v_��:�J%��@8��!��>U�dH��Ỳ����S�yEE^�%��$w]�ylYQ���y�G���p]da&$T�P=�-N,�V�ǔ��F�'j���u��k��tB2U�����	8�i�qύX3�5B-t�Dg2��h&��)���I}��D��{��ޓ�V?�>-|�Vqu&��b��X"�m|�O� ��<������z�&[P��qo�h��g������ N���ď@F(g>��&_�����y��)]���Ek�9�N+:�'�sGJ	�aw%�_.>��<S[�ru�4:4M�Vܹ�
	�m���w��1��̒+��u��Z�����妌y��2� ^�s(����w������&1~�Ua꺸�Ue�<�i�f�Z>��T63Ȏ���pY����1ٹ꯵ѶV�@��:޼�&Fo�h��~d��yy\��ߊ�8x�����0Ƨ}�㨣ҼC-��XQu���Z�����N�d���2g�|��j��`�����\�F
b�B��bR����¸7AU��.F�v�u�8c,�9n���>>_���� ��ۗ9�iq�_�5���erI�?�AD)�(fC.%�y�z'�t}�1d�8q,e�P��Ռa!nV�&,iI�
9���)���1n�V�����*�cL&���h�~������vsx��^�� ���q����>��%�G?��v���F�'���411�����L��i����H�_♗�}	/���~�"��d�f|0�8�=F�d���["���,9�1v{�*~�^'��g�9�yMb�ՠ
�����r�����W�]� w+��*|�*^I���ɼ=�_��=������G���{y5#���{��t�۷s��`Ȫ53"`��$�]=hr�u5��d���yP�W�7�ᐑCߣKTN,����F�к�
�^���[�a=L��TR���W��s��I )�m��~��0&(�=�C^��E}��C���b�C�Xz��L�[�E��	M�J��ZY܃�~E��0����R�%Z7-�f��=����4(Oj5} ,���28�5�ˬ�:}8z䦥qx�1�N�*n2_w�t��i͢�x��/�ݦS���O�{>$�<+���)�ܙF����֣����X �S�>��?1��C�j��%Z\�s�p�
� �R�?���
�Ⱥ�S����(}�С�ckp(��p�P�`2��}\������a��j��4�=�{zfa���q�Q�X�30�ɔ�vf��A�=p�kE�&w�- BqK�g:�%r��V.��`�0�24����"Z���[��B�3��:[�wa��o؏/��s
�MI2t=&�Ei�J::W�#�`?����g>ȵ��JlK pp��:F�h�91��1�6����fFA�}(]У��Eϡ �Ci9$�� �fD����e�U�I�aZ
,Æ��h�}�h��ߓU�\�j��e6�r;�}�a��k��x4��<��u���f����-�AK�@o�#�e�.H�=F�h�m�§
)��/������9�nW ��'ʛ&"�x�M�X��ǅH��ai#��u�6�`�����'2�,�`��	I�[�]>�sxuaI9�T�����ˣ��,+:^�����E�TD�y��xk`���p�&%��(/��cX��{�ﵹ]q����G����_�?�v>�� �`�ziG�cX,���= ��C��o�z��%X)P���f5K
����k���`!�����V�Dh�K�S����q֒v��V��t�`e{���B!n�xW=;� 㲼���V¾�6&�A�9��5H".u��O]O���&9?�̠�����|)J��<5�vT����5���)
 ����^���w�VX�m]w>ҚOA�2��j�&k�� ���,5gu�4̻��*�l�����K����3��m���ptRC�/zk���:�`��G��F�ɍ��-a�{C�����;��P�#� ���[��8M>�/��C���Xp��Z	xKW?���z8,��
ye"��x����K��Wz��k�ؔW�{�/c�����&�����I���y�� :�M�X=�<`��!���.ȑx�#,�����Z:���>'�����gʹ�	�m�kh����)����J��WZ�1 R*���Rh�VX���w(�0���#��o�����Ξ��gs�S����v+��D�S�XQ��I/6Z�\"�S�<��5o2���'R?�eӆ߆A����|\�w����dmw������H8��ͽ���$n[�y�|/��1���R��1�]Ir�A���K�|VW����#8�O.Ю����շ�o��|�i��x?_5�W Z�?���pe�B��t=mxW������7�cL�&�LF���?*N^��:��$�(T������hԵr���\П;��YB�����s>��:;.������$V!��&?����Ğ7���|Q;m��}-^8kn�H��zMH�L��(e��'9iy^�fQ�X�σ���
J=�W����.H�AWC���*�r�0��D�\�rO���T�{�S\��u��2vn���i^����)8��]�K|��_�B�YS^���_mMɈT�{n��[RW�����ck��"87��㲘�  ��~�t(����&����޻����׎v��b,<+K�/�