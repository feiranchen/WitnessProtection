��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�����GL9���Jd+ٵ���ξ�jm7��*����u���5Q�sl��v��s�n���:��2���tr�Y\Jn���;H�ht�C� ��g�`$:��	�Tƭ�X��prI�����zi��6��@��ΑD�g�!�@t��C��z�z��K#r�$���hF�ߍ�����)w�;M��N�t:T~���N�Xa�����LYO��@C6UB,���JbIv��<H�b��%����nu��)Ȼ��%��ͧ�f�l��#S�u�w������$5�(4uyc�CK�1�,��]���<mCι�簢nm
J캝��nz���z��n�p�n6�ۊ_��"�{peɅ3�	!���Չ+6x�D@z��EG󷛯�瓿֑��$��m����0*�w�*�K6ۿ��|8C����܋"��j_�$}�=�IQ��fi���z,POܹ�j��{��Eѷ��x�sB�W�;�Koc�'Y��������m�����-��l�3�w�|�2���.�p�W<'òh��Z���+���=�'m�Ԉ��4���:F�Ս�y
!Ԁ�,>��\t��}�"�|3Ve�����
:_)���I�?'K+�Xm��<�"�\v���ؚ��ه�r�l��!Ͽ�h�g�]wxW
`�P�������?AXJd)��B^|���j3ȺH�^R��n!K9(46{���mg��j$A`eCZp�V
�7�r�i��Vժ+�h�l��S����3׳����N��b����A.���54>�֫�6���/�a���WE��Gn��c���l���:������2���:���t������=�1m�N����*U�3�ή����,C��U��k�Vu�%)����Rf��x�0�C&�R�N'�d�A�v��\&��I�S-e��ތ��}�ϐ�?a|M�jh�CF��l
���»���͐x�7U	E����L�\b�:��\*��<��?%1Lk�����/r]�-h�"�Ŏ�m[l�
�%r����
eI1�G� ����` �^>�jyvj�"P�e��c�⓪}H��O�f"uT�/�C�xp�"�朷�ޚ>�]�����
�1�ޜ@��jvrȕ/� ��K������̧�>�hĔ_9�us@YuN=pW�ee0@#(�eL���v�~cS9��z9�N(�t����ϒ�^1P�8(S��"H�ɧt dV��+�gTéX/��5�vY�+v�I�OQ�g�hT=����{<POpG�T����7����Z<\�B��1³^6�ԋ�G��8	8V�r�e����m>v�<Q���`\�k�u��Q��77�ţ5�� �AK��$�o��W���^�ؽQ×iUGH��2��?�W\� y�H���\��j����)1K���oL�Y3�8�Β}�;�����l۱�9����-��}���%
 ?ςʟ���(�|i����O�Hhj��$b'�\٘e���I[ce��o������)����qI�j�R��y��&~�^}0X�=�J�
rU��I�g���%�_�'e��s�h�M�I��+-T�M�	�G���_1g�*�oYP����.��ݣ�b/N?GV+~؆�;�����Y�W�"^����r��|JR��1
<��RH�
]H=.�ׁ�og�"M˙�*�.6^��Ԛ��S�z#�1������5H=->�^=�87�[ś��6�A����"��v3�G��j%5�׭s������m�`z>A�Z�o@$[;� (}>TQȃ)�K@���FsY*��舺�*����|�����'&#�C}E&�'֝�������3�t��g��`����2%!�]X������,�کD
�?��'&eba�3��:���B�e@��X"~u���W��$���k{)�b�F����4�Uݒ�=N��+q�K�S�>�����O����
cn�:�������tz�I<^�?g��Q2�0���#+��t����������ԧ��{��V+
��2ğw��4g��:�;�?/��7.��9��Bciib�8֠8˱2�t��/��� 	o�X����{Rd�� ���Q?9��Sf߄tʾ�/�������q�{���uϕ����[u[�ۡ"i��ר����TM�1��H�1fǇ���b,"I[���r��Vm~ozCy��s�ao��9�K0BytnI�$s�q���6���2��s���sl�Q^~Qv����&a9�3ˢ�q��.�;���~��F�5�YշC?�%A�����	~���P�x~c�]QN%���d�w�x�K{��%'�:��-BTSCK�X�q\����Mq�W����U�#��:�rC7�n�M��tyLM�;�a,r�����z���a/�ޙߺ.\D޲����9U� �4���#B=�-�������nO�4�LzԸ�Q�u�&�t�Y=� ��ᯉ|a������V,���_�'�ὄNBif�+��ăsg�
����y�6y�X�� E�p��S�E$�A�7���쯒1���<����Ӵ�LMZ##�]= $h��O�Q���@7��>�V��NLd�}m�tFI����">�k�QQ@P]b[����J ��1l��v,��8�ʫ��B�D:���ɞ<P6Yuz
���t�鴮F�C�?�0�ek�9סM=��5�,�];G����+�����K��\{�>"f	1���8�J,��"��%%��m����c��mSH+a���p����j7�#?B��v�2����if�,��ơ��2_GݞC+8�Y������tX�#?�>�D�<�æ��
�B9�{2��yZQ�<,>j��Pmq�[��Hߩ �<�g��n��н$�K�?�ݘ�ݢ�"$��M�%���3a�Nu�*�_*6�P}	��^2� �MA���������\�f�n��[�;�����r����T��p��A������Əz�m=b7��Bsp0
-+����R���Ab�W-�#!�h��T�߫au���|NB�]��7��Ŋ|����!���JǏQ|r�/=����W�Z[i��4��sJ��U️�/�ï���J#ԭC#=�v��I���[�ԟ]�kqT�^�Gu�$"��n��F@,���B�]��c+B;tk4CR��Q�Z��4k��Ɂ��6�hO�+Nqc+�~��v�Y��ɢ='�G����C-�[��?[��_OJ��WU0*%���ues*����xtT3�M��JJ�/���f�AJ�
(�i����:;�l�^�n� *��y���x/�eEV(���Ѷ����,y��"�w��GQ�����$��`�_�Lb����(&��.��g�u���&��5D�"�pf��<	�Nz�9ln�9w=�&�7j�l�މ���zR�K�䙷�' �zS��%�Д�Ul��2f�J��o�PJ	�~g1�"�5J��O�/k03����6��J��|9��	�8N�n��?>�0,��xc�>E�u8Ԥ(��$�MHV%�`��z8�
5n�>�gn��5�e���ژ}�%ja>^��y��J�/��|3Q��Ol� $铋ug7���O�" %.21L�[1�� �
@2H�	<���-��0��wWW[0�\��c���U���W���V�`"Z���C�Ҁ�5�@7:?�g��`s����5ء�W��ئ���%%6a��p��7�5���-�g�u=���fp���P�OȈ�y B����ˉ�J��&�ۿ��i-n�F/�0�ٙĘD,�y\h�3�â��Z6��y3�G�ІKLp�G* I�q�]ª��^�5�8�ݲU�
(�^
	�-�䫣�_Q�>uW�CP��5�ܯ��4��-&���gE��]��9��x�i��GلM�lG�1=�M	w���49G��YHt�v�R>Z�༧5d����D�NC/z�]�u !��V�mӪD� �I�1��f�_��Sg������o���*�n��m�g�t�^��٦�u,�.y��͙��������aA��2��w���o3���zY�]ա���^���7 M�R0L�g�j��K�J�������A0'E�iAi �.������<d�,Y����f.��69�:�t����c��!�"/�j�)�lE��H[���-���o#����4L��*�	]������|����˥�5ȋ����yM���y'�!b����^2��(�շ�D��wQJ�$��	��(M;��B%yj�m���<�8_���伦�
����	Y�9g��?؄�o�t���_fӃ�zj6��-��4�?�������׌#q�R� �+�m+��l�=�����8	�ٿ���$܈�
�K�y�)�+C�"�!gx~��G[`\m������P\�ۀ1X<-����/[@c,h��cP�X+Y����H�J�{��]��@j2�]_�ϥV=��I�e¶;
�[j���~V#hΙ���b��6���;�=���t�ŀ#�H�?wΖ�>��P����R�'B���b ����-��+�3�c�ڲ��sSk(4� M}��~���3�
w��i�T�gz�0vK�?\d�k�����vVK�-�>^�e��p�A��y�a�m��92}�Z���B�-���b��tuO��,0����k���=f3`?��l�۠�`�=��0�k?�~���g;A�]QR/��IѹH��g����4E`��x�-_�կ�u�9Wfv��ku��[9� Y�n�_O᎟�5e<����B���sN�� ��T���kݺ�M4L����nOx�cg1f^����?�?�����Ȃ\JI��6�{2�N�3+Q�ؐ�I�#e�a�I���JN���R.6]n�^�dԲV�V8��^Gz:-}�d�4�>4��zȀ�u��۔�=��[��4d��-¡��cnW��x2��H%T�d�������
!hꕨb�/Pqg��	t��Ù?�T�=��0��j�U�΅Qzi���U���	#��
x������c�z�g���`CIš�x�p��H�l��Ğ)E�E�r�^kG�G�r��ݏ�/���`�B�/�`~��>����g �0o��-�F����B�]���֤M��C�#����$I���r��)�X5��\v��I)�]��������`�v 3�#�I0�t��&���K���i��=ëO��sJ��������΋Y*C�.���u�a�s�{R��$�����d<��ٌ�	�˃�a� �� �]��Q@&� S�TPpVEL�4�O(���x��Mc��ƶ��%#cuˮ
��&��}�Cd������̈˽1x���8?�=m�?����H��mI�N��p�1�@�q��'�&�5��]��d��6Wx!8�
2)�V�99�[��'�RF�x����v=��9Mƚ� ]��8��>~�~&�k��a�<
xsq��)�e���~{��be�ڌ@�"8��ᢐ����6�Ю��:4��e�7���/ѣ2�p4��	�7�	<h��{��&�1�}�(y�c�ϻh�LH��,�u����(�\��֪��X���@𹖞���e��:�	z�!Bmp�>� �c�䶜���y�Şz�P��=*n�yr�k���E�x�]$e��jۄg 2���m�=d��)*Sr�_,�}s�P�e��yf�>2�E��{HS���x�۔�B�RR�,�����W��_S�s�'ߧ#Ŀ?R 1���	��l�$͔z{'k2�<�:�`!�F�;,h)�K~��6�(��5@�E�sOS��>����ts�à!Ja��J����-[�q��}����%%����6V���f��/5a'M\Jq�������_ԉhG�̔�V���GAY��i��N�v0MË��B��70T�	Ԙo��	6+0���I�c;.��PIu=��q%����U���0A�ӗ��`���@�^n�op�qw����f��Jݯ:6�А���"g۲�����%�Λ���O��aҪ�װxq���َ<\b&B����t�	��]F}Ne��G���wM��ج|�����\K��h컽(����QD�����_%]ujA_$�	��!-���%*���=vov��{	�I�Xs5D,T���%��82[ېuN[@C1M����C@�}$KHZ�TM�*�Zt� ͧ�����	�3������m�U��֡ba�9ɷ>�p���7�Vٺͺ���9�����;�������H�
(DpR�mT��S����ʋ�k��lnv��|�=�]X�����`�M�z��߸�:�M�1;�F!�/�nK#l�~M��*k�f�`*�5+O��Kfk*UV]�^�
�]���j2z�tB�l�E2��S��@���ۣ��b���\y~ǞA���R�����*�6��N)qH7��z��yۥ5��4��[��L��JuΟ�����HB/3��U���'TK8�}'��?/q:Щ;Fǀ���`$�4J�!���m��R]�{3�2�u?�\[&��W�xO���QdF���*�&3��j�]�� �>�⒦��x��/
|.ցK�����7�9<�iIɩJn�J��������>�V����1����cEz��a�P2o�*�9�F
�VC�y��	̡j�\�\����9��p��S�+��v���i�'#�ۀ�d�a�s�y�+yRD�lj�.�]d�6�"/S���
ǩH:�(���uqZd�>Wd�'��?_��v9�vC�.��$�P˕��@Do�����^�M��;nYԀ�,y�.`�]�x� ���(�'DC߿��D�k(�z��p�+e䧛I�u9�m�,6�*�k�"�U�#O�}4|j!���j|d�RV ��>��J.��$Y���gMt_�0I�v�/P���lޠ@Pn� ���P3@�=�}�tۋ���D�oN��h��#���4`d?!��_���Շ��5:�z�[���7S���B����|�����(��г�)�:�ڬH��<���{����`�?�һQ�ŕ���ҷ�d�]57���VY�S���Gvj�w�oD�8��O��	9����ڔ֜���۳̟�qW� �.����a7w�1U�r���v�Xe����7��a�ߍ����FVB�:T��7h�r!�F��E�����Y�}��kP�i�f���B?��
���Rut4�1FP���O�L��鬞�����<MQQ�~48�}������P�G�i/γk�+��!B/qБ`��G��vGC�j�!:�2�
�j�ar-,��0b�gqLUµ��׍6�v�'ɀ��⹶L��p؟�=D���b��W�Z�̿���/J�v�qk~@h�8�#�[R�Ͻ�S�˲�,na�:Wu�`����eL6�nIb����gc��Yސl����]���-��=r��i�<C�\��H0���3S�~n��~��#:�_0��d�U5��P���Irs@S�&�"Ahb�{��`��%��)/yf��^�fa���(�h*48��?�]�������Nķb2C����ϳ�V3�(7"�%k%���x)>�떙ă#M!�ɖ����hяr$�������~�kqQ�w��g��B7V���mA5gQQ�s����w�f�Dz�^r7D"v�=Y��G�1�@c�z��y��SkO{��Θ�ڪN�Ե}��P���9�w��Ȍ�"���wќ:!��4��#�}g￪��Ӷ=!MA���lEW�TA�[��=O�K�g,Xx�/� �ZP����`��£�����{�(t+5	�m����t
	dP��%3Z�*G�,���֎���>�lh���WK��د�?�0�������s�	vd�x�Ա���C!)P�UHH�bF��3�Y��&?m��������!� '픝�(7��-9���歛;-\3<�X¤����R1=ri{4�ZZ���g�OT1�7�y�0�!�[0jk��<�}�C���X����^-�N���A/R%T]�B�=#1dO@A�A��^8
Ƨ��i��z؋T��L��>Γ*��K}������C����x�����n����`6LQ����Rz�>����p�n��z���Uݥ#���QzF���d,��a��?�n޸W+����e�����Jb�[V�8n���`���@9ț�FVѽGS@@�N1��0����nlOqV��h�`Ʒ�<�rO����c�&�`�ur�qc_r3�
|~�S�px(�8��Ƃ	 �Ra	���Ů�K�9#a�u�yw�S�$�9���҂rK4��QIG�N*M}�T�g��=D�R��'�*O��z5���RD7fp�Q�/Y����MZ=��=
E����{:���{�ľ�l�ĕ�d�(<J!w��<Q�E�D��D5 �:Z�i�x@Y��,�^h�F��Ϩ��$<����6��#<�#!����y%�z�x	<���(�
C�^�#�
��ry�D�4rG�2�S�:z���g���d�r���͖���s���DZ�72��	�>�;Fa���M�����"����_�'č���t�n�1��j}`!0È�A3�nJ���9G^PGl DH�u�_)�Q��z�t���`����n�)!��E�!X�ȅx��##��^o���+N��7z��;�$��)����)I��|G����-dѹ�	K��8������R=_ZC�!Bjl2�u�..�F�5I��u��61��7�A�q�<�@eq��~e���uRj;�-��ʕ��n+��� ��������K�V$y���2��h*�87��O�����o+�[;��I&J�n 6�JD+/r��������.^�n�x���w.�δ�&��1�����M{K�3w�m8�O�A����GD,?�n�r����K,�m>�hZs,��5�|;�O��z��W�� ���i���/��<�]e#�*�g(n��o>*��'�T$�j0wu��>��Y#��,1���EL|{�K��w�ԯ�*�Xd�v�������QpCa�����Q��`����&����)p3~4#�R���(Jbh�](
=^���T}�ļ�����"�jX�����6��� ޹�,��*,S��v� Q"cm��Dk��K������3�뵴�*���'x�ĸ����y����2RF�󤋯���v�
u�o�l�.�Y����?�J�/!��'�	id�^H
���F�Кv(DF�XG3(O��U�*MMy#H2
�L������0�C�^0�U!e/B�;(Ֆ`��?���'(}F Mg���%����ٿ����@K5�d�vB�f�J�:J��R�\Z+��J��)��^W>��u��`K�gҷ��>��J`+�3������lg3���$7#��@|�FC�x�2m�5�ن#���_�Ե�<��1`�L2�/[�N�S!Ա��Q#��4�c[��Rg'�Ȕ�q'U�Ô��^��yyߙ�J�ld\ �a�(\rpRd_9� E�����+��8.�;
�0�3�V1��eq)�s8O�3Q��O�[��d�<�5H�K������"��7��]0YO=�GR����P�����7��Y�1�ab��P�>�:N�^^�˫)���i��p����������=S�T&3+t��o�c\/���1(=�J^H�1�!�}AӂBUw(�9���������uuHn��UB�`��ꆁ±t�~ n�U�>�l�2��s�#�HI/~�<��3�|noA+[,�8�o���q����a�v��U��]\�ľ���~������5\FK�&�6�1}<�H�5��n	A�-�\i�]a9`����yԆ�
2�|e��̉�y�([�t�=���ͮW�ny@N@;����#u��R#�0�"�dz���f��)��Y+�.�M�g���G;@z,'�k�OG��݈Kr$�4V���-]S�-��x�̖�w;�G�7x%�w��RT�u9�6,I��1���.	t�9���m�&:��&�Ev��"s�%�4�n���d#�f�-֋�y&j���_C�^LP�'s�|�&1�7�5��Oz�W�j�͂o�i�>Us1t���ؽ���4���z�FǊas*���ڭg])��"/��p.Ͳ^YL]�C�IM*,�RvF�8���x����!����3��0�տ�иZ��������NF���,WAp�1 ?!Iq��H*�߈�۩3w��K��u߸��n{-�Pu�v��J�� ��/y�0�N���T7�`D�a� �H�	��g3g�<L�Y}�{���l��7��������&,^"��b��|��wwI}TRr(�Ww]��y�J�~�m!1E���Eg��-�1а�u!n�d7��ǧGϺ���-�r�ܮ�!xgT�>ǐt)6NA���2����o�Nn����me?`�S������P���0 1�0qD>�=��1ڙ�A���Zl��,��:x�g�j(unc�	�M����-L3"���U�.r+�
����X� �Ҷ��u>� ��>���J����6Ja�#h��*C������4����DMr��/bá�8ƙ`P�b�h��1,�_����h�ďG/���k��J3�\J��d7�T�g��H�M�������H�n�뮍ڀm��z�3OC/{Od�n^y�?���m1�p�:e
8�k�n�T������9����1(	���$1���nrzJ>�rb�O��d.S�A��y�cn\���;�YM�oV�bb�'���U..�}.�G������C�*ܛ]��;݋��B��/�-7 #5u��L��������-�ۼ�"���lq2�Z���|s�p}���Uy�sm3���L)�!��dYs�i�E�)v�ON�m'�<1� bsHp�rI�^A���@J��Uoͪ^,�*\���!��,��=g��mPbbP��8[�x߯b�W���2�q����ݢ}c���uH�Ⱥd�Q�5TQ� �C�0�dܭ�UN��rY�?K<�.�H�0�&M��A4�0@�qj�be���1,� ��̾�:2�ך�Q�rXfY`m���Ψ��{ΰow�AJ���ҤBd�����LM�,+���lu2#��ՍEJ"@�$�x����l�U;Q�zj�'�>$�q1g0y��mbq�WV6��C ������+-E�h5�x��ZT�"�4 �wG���۲z4؊�yf���vE�w�z0�A�`��3O���w�QfQ_���W@��	�J����J���u�y���'�H���SV�-�ďw�G"Z J��>}.L���.��3�^�Jz/"@��Uw��m��E��u�\��l� |��#�M�~owwa���2(��)���LK�W����v�����l�v^ީ����	�,fs+g���̋����T���%_��F�fh�Yw�DHue//�ԉ�N9X���V�O�U[��f���@au�*ļX��5�n�Ԝ�#�);=��[���S�\�4� �q��}=c͐T���`o���$l���kn ��\����O�n<����bAAϴ�5;{�L�ۖv+