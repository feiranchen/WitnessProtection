��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�g+z������b-�ݦ�e�Ow$�i�y�{/ʳ�q�c������޼������iqV�8���~�u#Q�3��hKu�Q�>���)����	B|=U�K +�������0�$3,��;g��o`�!�eb�3��Td���n��J1�:���W�0We�c��M�Ե����{ԐQ�JHR����@�����t�h?��|���� ��rEd�t�(�b�^�ވVh�tWq��y�ca���[��^�Al�t���k�qq�ةí'��Z=�;�$�Ly��r��هe��4�t�b�*Qҧ w��@�@��$��^;Գ�j6�Z����������8�7��b�lEr)K�qiD��{�ZԩC��I�0��O�[��z���e��fڏ�y&��y �����Xj�g������j�0L<pf�Q�"OB�kL�� WgA����\}�V���<,D�~',Nm�)���"!bK;��M:�"q옳;,�G[}��8W�F����FM�a�/����h*H�k��Qqpޢs2����� :5j���'qrC`���'��?��P���K�C&��n��Ϻ7ش�������RŪ�1��@:�B�Y:�Ə��8-���iu�ݝ
��S���?TE��.��Av�J2,n�fQ<��P*"S��r��K��O��_�Z� U���ԡ�^Y^�7��EyWG��պ��a �%g���5~���ʜ������1Bώ�Dx��~�P�؝����N�[%LF�w���W5�y(ѽB��ƺ�?Y�J��9�J��-�N$��Sr�\����8�r��6Ŝ��dz��ъa�s� �4^]A��~���{;�F�{r'�I[�Z��,���6RU .�iˬO'eB�QC�$�_�v�c��Z�Ƣ�?�O2�9.�@�["��U&74�B|�Zo@v�N_�\���S���$m���%i�=�F�[-.g�æ7O�P���T���&p7d������@��A#�/V��b�E�l���д�ԛ"�hoZ_��Ւ�Y��퉗 qLnu�y����?�G��w�C[\�.X)���P��n.��<�6�^��ٜ_�Lu�w=����E��F)S�T�t�4<r9{�t�)���^O��� ڙ�n�����g��d���|�$2�w�Z�Ćzj�K"��9Vt����~���<�I5�X�J����J�0�� XO��t�����^v��M�y�߶v�����0})o}m�ʎ��8�	VH
x�g��m��-�	^'�R�;`��PKʯ �_5�Պ���T�R`[��0��8�/'�W��=��5Ь��<d�ҧ�vi0F"V��֯+�·�B$T�˙�R�W�/%��4�d����]
nh��edc!�Y�w�5��P��Ygr�&�)��4N]F�%�+W�U
tͰ/g��X�"�Շ�B��1.�h4Ƀ��ܢ�`�b�Y帩����4�^c�%�*a��[t[�k	�x��j�|�ҭ�b}����h;Sj��e������p������8��PYw�c`m��w��Apr�X��ȴ���'1_2P��@�~W�9-�9xٙ\^>��e��G�"qĒկ�9��}��]>�_y���l��}0����?����p��+�q>arN-��X��p{]7i��1$\�����]Vo&�����@hE��16�Q�j�nc�_���]IM�b�T��?߼�7mї|Nv�t?�߇��fc$�$֚���2���}z]�=\.D�}>�Rk����p
���L�}qu>�����'Fܻ�>M�i�X��҃o�E鏡w��ҵ�RQ��="� ش��	%���cX�|HVWFg��_xw F����βl>,���������"i�&�zj�sB^��=pc�]���z�w�7�>��u����i�$T9�=�h=�{�^��qj9��P��A�|0�=�J��2Y���W�N4���<�x��y�F�I�/�!B�\>/s��5����3���n�?�=_�[��{�����P��-
_���w�u���(X��|$5�%�MUPH�A��"�^WM��oQ&H:a[�z<�f���޶N��^��x8[14�B�l������LF8�Km;�vي?�����F��j%�O݋�0�?�F��$�A�8�S�����^��)r�3�o,���R�U��N���v��l=��ٞ�<J����j���@�n*�U��V����9�������k%�w�7�,����nrKz�=���zx�<����{vî�{��j�֣zD
��S�iG`vOa ����n�SЬ��e�.r"�I߽.���v�׽)�ɵYF�4�O\���F�E�5M����NJ)��<�,;��:q�m�S�K�l��w\鴩���-#d8e������Q�ԌYM�	o����]��r��"��享�"��H��s�� �����=�\�ՠ�[*C�ʪ��q��v�\7�	���XS/06:?�\��G9���EM�φ���h>������ϾregA���8k�,(CU��
���]m�جjIJ��~�H�ҫ���%f���(C�z�lk����Rs�&}F�p����/�[B�?�"DRk-�XZ���ho��:ᡫrq�蛷#͜U0��5K���}��~�#�^���V)�z��6�'@J����'���i?~[uak�$�(e�>��$d��-�� ��9"Gd�(<n���wn��Bj��
[F)W|��*�c���D��fmWŇ@\�?�v�s��,��uA�(���@!�yy�"�{|gJ�"ʔ���O������A��@�Z, �=z���p����бA$(uh�Vs���ݨ�/l$��N�u���*�w�ſ�72���u�x��^tc&���sz� �>[�(ޞ���1���B8)^��F�>1Lt_��oAĭŝ��u����C�o��7(��:\��C\n�z!�v�t��r �V�C76����>����+�-�>G������I:�^Q�"�*�ih�m"gb2��`|�`<ڸ����n��y8t��Ӏu&K&s��R�v$=Ӱe�S^0D��@#j=�ίw�7���T'�a�������
l��1��l�0E ��K{;.s��2�������S��Ԃ;�w&�F�;��l�3πw�yF�Q׌ Q/��,I�O�����5v�-�t��oalKԦs�x���Zm��~�T� ?� ����b�#N�$M��zX�� ]y���Y܎,�l���0�L��>N�ɣ��A��v3�2�a��Qy�{�#�c��A���^�D�,�׍�,wy6^i]�����������>}�_��7�Z�F"�������O���A�� �lns��ؐ�̀��'��%��tI�J��(�L�PR��`Ɇ�3n$�^&�f8៰ʻf�e=B�//|�Y��U�݅�_�E����
'ݰ�:H���Ʃ��Ќ'���#��4��Ϯ���ߍ�"'Vɼi�ˉ�� ����$�ϖ���!�{ѶN��P��S�B�o9E��p��|?,��#�2^_n�5\��B�"eЕd�	#-���!�n�_�1y��$�7�1÷���f=�ɒ&��8,1����kT+=급k&�oX����Pb�S|V7��=#Ԡz\�n��S�-D
0��3P���^|M�!��՘�4�}���|4��F�&]��&�k,Z �P?��P��4�:SI�.�y��c�L��N�	��^�����4z)'(�\��%2�����F�3�괝���P�	��Λ �2�3λ���id;�%�y?������?w9�����̳���D8�G��RS�y��|�!�i�sf��:vMg�k��Bt�fp�q�	�H��'�������xj�?�6�@������I~�i����LŔ`=p�tuM��޼.�����{5���o�Ԭ*�sAV����P׈F�P�1@J	NF�/�,u��IJ
�����yg�w�S�*7n��gY$������*$3��d>IV��#�)��H<���O�8Y�y�4��څ"����Ia�rEJ�| �����4K�_��>Vq�;���ZK��X���3rK�������MF ��Wmа�Wq/Oz���}&�1���W=��08���G�SI��u�����m��$�c���a�� �+Fb3d|_7*'�8��ZO<�"�kJ�����6o?@C�_3ĂB<����Z��6O�/ڭ��YH#�S�Ԁ��w��S) ��{��Ea�����,T����� n������\Y�גG�
l��[�����|II^-=�72�QeI�v\�I	K����$H���D3�~�#�ªIV����x%+<�G�EZ��3z�}G�Į5x�Su�O.0�d��ajTK{���ߒ�w�0��'��sAF��Zƴ�}�^87�1�JU{p���tS/$7��.@Q4@���X��D<����>N��[�Ѫ�ǅ`S�sf�_Z����a�4x�ֶZ�ƏX���|8�s�q�(��W|k��l�ZM:Qt�E��K<B�#�������Y0 �Z�$��t κ�닒��M�6�%l���tt�0?CJ�scg�p���t]����`75�u#�iL�6���D�Q&�X�.k��QU���4�P�\��۠��Sw��=v rny1�/���Oj���)3�,�J�q��\n��R[h��r�U�F�vN��C��UJV��T��[�Rv���r���7��)f���w���z>��������wDA�b�S��x4u���!�i���(�������e�3��jB��Ʌ}�.�.�_��'��w���׎"ґ"\M)fJ*��7 ,�>T�E��t&+�aX��������-�a߆�ܵ��rB��_J��A�*<[�sYͦ���۝�|�7�9�o�G`a��1�o�b���x �]���-��#I^ɚHu�?�j����L1�.��YT�su�n���v,�k�Xt�1d}  v{��� ���8T9��/��ҁ0��eZh|��h�*͊�1O]�u�7�h��ȉ�|E&� ������ �H��&��^�J�A|G˛9&�>Ə�~&���nhG���$�~t5 �օ7ϸ��9d��#K���o6I3*���3��A�Y<(�K���p�;�Ӻ?��`5�쵺}�w�������< �[|_��z���h4L#4�K�vc��p��7�^��^�&�������ZI�*A��3�1۱�=T�D�<iv���Nɘl���+#��+&�Ha��M�Ue��z9nD_�őÝ�o����T��v�R#�0L۲[��P���=d�s����q�P������=W���Uu�9�yNzZȴbϢM�ʺv��e�Μ��t@Z��0�O'N�U���/<�?�9�bq�#Z�(2�"��Z�c��N����Akw-��p;x�&��gy=�[v���Zo'٨w�κ��&ցط����c��a!���-��7أ�۔e&yn��{Ŋ�z̢f����B!�(����UoJ��2AYD6�]�.��#�"���D���\�5ӱ�o�z�R],*-�}�*ѺTr� ?6S���,��5Jzz�:���#���ӣ���N���q���O��*}&�@ ��r{���#�^oi�Ŀ  �eV$�~*�L����ӌ�Vo�s����Ƣ�rr�.WB��؋��S�f�U��������V���J+מP�)�ov9l��_vݟ2_$Up�o�������v���c�:��*	Z���`n�Oy���g+�4�
n�K`>N�p9b[�����+I���f��S� �~f��x�If�4�޴��
j��Q�O��g �}�0����y�*9�:��$|��_����MSR�7�ܔ���-ۻ7��˕kJ��Nfi2uIL���7}5�=]k���dF�̻���(%I��R���	rp�dZ/Ghޮ��)�l ���e=�B�ㅩ�Y�3u'����C�v50��x����8~�n����8��u4��j�J��d_*�!����8� ��RX��\6c6����LV��n9�X�)���Շ���`?���L����F�����[��/��c�!Z��gr/��/�)����4U�O_I��M�Su{�=�z�&jǩ��E�3��rdxe�OR{�ᐵ��+C�7��nb�eB*d�]8�c;�
Wo��sr�)g�����\I���<�ో��ɐ�Y��S}�2�O1�ʚun�KK|ڸO�&ɢS|���T��:;�+j�Ml�||���(���ɼ%,b�2mp�gB�nzdn�`g�\���}i �5��x�r�@?g��}���3�?�S�Bi �����ά��l,=��=(�>��ћ��0� �^+yh_a%���!��3c�JT��E�Y��LS��Y%!�1*�̐����� o���h�'�Zv��O�ˈS[K�g�I{(}"�5Ƹ{�	�7;��3�=�H�U(���:���NaP���:l���_I�U�N�Ϳlw �����ޭ�aT�5��1$��$���1�����+��27����V�R~�H��b�.�u�����Sc�j������&����|��^�R#��-w@��WO`��h
8���w�.I]���"R�����6��dӯ��,kZT�����j;v�z�* �+�#�J�٘jy��gv�*b��K�T/�W?�D��lv(�0j����D`p��.�K+Ot<��B�X~Ҥ`�����$�Q#A$�_lQ�(��_���}^O���X��y&-��j�}��0���5��V����c�k�#�����? P�\
V������PR��t���ٍ�Isl���B�Cd�������ÔFV ~�Rj���@Y��;�N4�M��O�w����W52�$��5|襙Qr��ڂ$=኿.�B����X��UJ�k�N�/K��kӵ!	z}}��ʽ\� އ�G����'�hEE��rr[*j����Oۭ�b���]rf�\F�z�_>*�0 "�N�����S7Q��,7 �hOڢ��r=p�#�����^���m��yɼ0 �����I��䗾�*�_1Z�(;.�W��і~�u0�IC��}'W��W��(��e�P��%��ͭ5r��L*��_ߣ������́;,�k|U/ ��
����lk�d�j��-?�4�>͞d;���A}���*�՚!{�+G�`S�T�[�{�ޗ���_Et�G~���fb��/����x\,<��BW��b7��1Մ�jgʐ�hfB�kweR2�F��%p�@�#&?�D�ҵ^�U���O�g5�#���\�CD/>��O�?��2s<��#������ݼ7,gd���s��<�?���t�kQ�fK �Q���L�̙�TI3�5c(q�����u~�kA/m_)N���_��Yq|a�U������C���#������
�ԍ'o����t�s@<fü�#�.�I��!c�C��S�x�ʊ3oR�qta��+��"��OeC߰I)�J�-ւjiW=�кZ�\�lL
"���@��ӄ�/Q���b�6��"���hCw�Iq�uH���r�P����J����� T��.�N�ð^KtjX�>Uf��b2Bu��T�P����@u��Y�E�{JZR����^Dr.sl%�z>$�oϙJ�sp����TO�%�b��rt�k�������ʗ�n������*iA.�*c��j�V���x=-]���N�	�@��u��!��t���_9
���n���ɥ\�"G:>kv�������D�ܘ�E��8s��;>�2�w�;IQ��F��(��@��fw��V�Q�R���~(XV� �D��<,�$�����sc�1�4�w=Yߔ_X�ׅƁ"�L���X�`��Rt����J��aj��T��۾�K`U�_qS�e�L3�}����'��N���z�A��[zz��!|�nm�Χ����Z籲�.��~�zQ�.��L�du��PcI��oZs�+=Lnɉ��iQwe�o!i�p�Q���Kk��|���^���Iu���o�xl��c��l�6�1ꐉ-m=�{�z[�+v�3��R��܊��e9�����F��b�p�<c�ε���N�9�����~��n/o8p���