��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�5��3���}K��H!CX��C�T؝�`�Rs��!��e�Z�� |�'��n�P���@8�e��s>�}����c�Z��a$�xAyQ��P��?��7/)�j0ဌ�t�+�%�Q�H	,� X����.�h[R�ek\�B穔68B�n���S�71�O�5�����r�������l�0u�Q���Q��#��8�K���!L'�Z{�Ø�w(���F �\��I�9{~�De�aTܓQX��T���\��4q^�%}�IH}<i34V�}��u�{��=n茡��~s�������M���GIi��к�M���U��� 0�o�b5aDR)�%����H\6�x뻥y���g5����6�F��0�G�"�-�y�i����[��査��W�O ��RB��r�l��ȯ<AT~���&JlQy��xm��� i���y��:���|=rdX�>�p�J�T++�f(��P�����<��ُ�dx�#H�N�Y�8�;;%6�{��)O0+=�8�H @�S�RUA�N+;28�ۊ�C�D��^Á��$b+0�L��W �ǲs<��`���=D���x���2�2gT��죇��N=���yGFi���N�ެW�C�8��S���.�Pj�_W��1��N�VD�p6�. ]�����,�NE�B��J�Ɨ����T�z���p��}r`I�2v7Q�R0;O�ٖ��$�^��/�p�[uV�;V��B�ߗe��^���z��\k��W%{R$J)��J�g0��Ic����U���Y/��+\�t���!Wi�ގ���NAc����֫D�eA.S1���OSoP����/����<^[�E�:X:�4�6��:u�����"�~f�MS�F)tľ��s$�'[�	:�H�����ʸ)�@w�[�0��$��?�T�e]Et#� #�<�����&�-?�3���i��/�X�Hv|������S��ڧ�$�-�ZxP��"/��L�� ���O�cPE��%vO֟�+��H�Dx��)*]��WMoK��. �'�69ߋ�� ��Cs=*Ї�!䧯������-%�G�cE�K=D�\*<��(���C|90�yE��N�L��~�D�����i�>fW�/�BT�l);�9Z�42]�P�Gj̑U���B���t�E�|�_�x�w��W?+e.�;f�t�Wh��L�K@#���Ù���3n�}-k�u���huno�O�">��p�<B�r@�L���y.p�vv�?�L�]a�4�Z�!�����}mÜLl{�F���)�0,�u!
�	ݍ�/toM<�L̝WY�C���SM`~���UVP�2L�^�rޠC����8��x��
u�-PWc���ݫi~�`M	�X��yq��҈p�Hw~�-�� �nD4͎fjx�DN�=2>����ǹ�Q�d�<��T��C<�!�Ԟ/�u��!f�g�S�_�U�=��T��8p�.&�����Ҹ>�+��G���Rt)*�8���Y;Ѳ��f��f��' ����"I�20�I͚�zZ3I��b.9k����αO�϶�`6��L�M���6R��'k�j'���:+�08nI���\��F&i>3��'3	�[a��]܅��3OՋ��)�#���8�¨���
��j���ǓM�4ן�+f�q�Z����p_��ѸFo�X�3.G�W��V��[�,v3t511_g56�;�B�{⌍�6ѐ$4�_>_�&���я<�{�ԭ�Dlmǣ�������E^`-�Ӓe$c�����1 �i�Q��n#k�������Ϻ�Bs_�"#��������$S	 ��V���CɌ#�x�ԭ�ϋ�iw���ǝ�N �,W��!�SSѧ~h�9��A��I�B��9��
α��J��= �v��F/���Ŗ�)j�D�K��ı'q*]_��fh֢^��<^E"��J�����f+7��E>2��Ȅ�M�A�k��F�ܢ{�e��2	�٘��%͡��k��v9�j��tͮt�L��%CX��, F��z����]���Ǖ+�1�7�F	#�
f�RmQգ�@��)�5��a�B5��8tS�t���lư�n�����D�#��"�A�OS.}1��y�JW�lN��؈*�=��]<(���vB�S�gn�����|H��s�/�0��KL��N֯ģ��@P3c;�m��W��ɓ�T� h��2��<��;���t�l�;�ѳb������5^c٨G1����q���$��M����]�z��I�e�fsb:1w�A|��?��;�<�r��BX�hjw�^�㻠[��m��Ek��|gY�`l�WxR����˅�p���k�;��B&���~���0L@tOEp�`n��JwjiS�qo�G-�����|E2=��Y`�I�O�߲g�D�6xXQjں�B�*9樞:�.��ٳ��&g]'�(
�h_!D���������X���������i��Fux?�7����2>`}G�_�fȾ��ȅ���LBf�E	5.�&�Wg���,;߂��%�(� t���h�q����hG.��9�|�����8 �GT!$��~{�HQx{O(r�9��Ow�P��jpì����!x8�[�fO�=�+F�k֬�0�uP2Q/u��������s�D��S��r�m��g\�7.}�܌�L�]s��G��6\F�F�{��8�f�U:�H洕�*��K�S��><9Y�$# Щٖ��'�Vd���|�jP!��{�y�(Z*RjIe�u�j�T�)ն;���}��EZq�T:%�!�R2$���b���HciA���A��~��L |��N|��H�a|�`��W*�.�-J�I���X�:_�/�ĺE5ʢ���a�?���i�Fep�lLT���{�uFt,�)���;�l�E�Z�6[^i^�Y�t:��G�v�v3U��i�� �����Bz���9��) F�^^�9�Ύ80��u8�'��Ag���R�x���eG��e�(<0���n��2%�u>��?�ff�K���jR��h�r�)������P���~~��/�Q+�ֹb��B$c�&*�}b��Y�=�d���X9���q�k��l���O�[x�t�K�|4_�:!�5�@Q��͕�F��V,:����]ՙŝ���P��te�um�v����w�dIn���n}�0���ĺ�Ž@��-}��tV���V;F�9�-S�S���띦�o���$	a0�/e��9
�4�V��8�u�Y�Iڪ���g�|��GA�)26��d�}�Ȟf��%���ÿRgW<�ȹ/�5�d8\t~�t���.~F;���8Js��I����|��ŷM� ����&NZeƛ���el���o`-�i$���nꤧ7a%�Wl�VS�m�D�-����Ⱦ��F"p�S��fs��
�"��>6Ed�́/ܡ�?�	bcXYv��݁�6�S0�-{��_�u)kF7�#3�=��ǼDqq�U[ƆQE�,���,�½c�O{�{�j��I
E ���Krq��� �N��>GZ���ٰ��'h�g���0xy$7s��ԄΕ�����X���tORju����3�XX�pm��u����e���NI>��Psx�.��R��N ����>�,����y_Z�]���z���-�,���&V,J9�;j�w1ҏMܘ���	���Vi���ű^J�Ca�cfe��^��V|/ñ���eԻؿ���@�>�4�$zCѺٶ��[��Ϝ�pvK2KH�w�����^�A�/��x����݋�4Jnߖ��4Μ��jsNy:��H{��o)J�>\�a�.6�J���M�(�d@���-�x˛��:���B���yR��1l _�>y�F��v��]u#�˙�E��4f4�ꌱxh�(-]Bp�e�;�ϵx�|/��=�hG������Y�$T�j��}c���t�@�o�tZ*�lJ;-޸	+9~s�/�����/;�������n �=XW����~l�(�| p �	��z}�D�5�sgO.�Y��\V�h<\�9Dlz:�U��3ీ�k~��{]o�ل]I���j�!�=o�愩�z�w�O���E�a��"�v.&ʄO�&@���n��h���t��@�&"��o��n)f/�j��Ճ�߹)��}}
\������t+M I�*fTB��}���4p�r�;޺S'�5+��U�j�L��փ�>�����~�Yo�L�4��ě�+z��Vy�R�(A{r�(�?UE|�:ԽD�Ȉ�eiV�P.�BL?FS���ߠ�w"�<� !�5>�J=)#�;K��!���J[)1�s����5:��5�/N�Q*ZN&F�(���:�����W<�)b:<k�!a��Yw�J�����
�K���{�x*-�bi�,�q�,pǡ��Z�z��tљm�@´�C�v��:5ݩ͘��/�"{1Di�|���',[�"��\�o� ����wE���^ z[��:}��ǹ�lebp.���3��"�em��a�]m>.��� �#�l��i;�H|��	)Y�B$GtGx��J�	�X)ѕݱ�*��14�'�������!����S3�轆��.���~���󨖤ȔF��0`g~g)�.��J~�jJ����X��8]�yč�������`t�>�7��6�
L�reW7��S(�T�SF��@ޫzQD�x��[�M�Fo�ò(�_��~�3[*Ư'E6n�a@���@�m�ȪZKr�%ɸ�Z��Z�'� �j�$���_n#��ʑ$���G�K�+���wR�u��X����N̶=��@0���+�b��5����of�wюCU�ܝ�����,�7�G��o�8l{ŧ���.K��wnt�oTu��)w��A§�]���`�o]��ILfJ �$���Ó�P��a�����"�?��B�;.#掣������}(�gZOX%�/���\�5�{�Y��;\� �#�pU�,}$��7����+}*�a|5!��W8�O3��#���\
s6���n�E���
�L����m%(�Ta/�;�XYn`��
ֵ���;S���J��7�T@Fq_�Q0�ރ���t��6��g�aB����6[w�9$�]�{��*��|�،ל�R���W�P�Nƾ/z��
�F!w`�-�Cۡ�>M4y����ʘ���2Z�׾M��>���L�Ie,�8���X#�|I�cj}J�n:@9)tptQa��@�ત�5�e����jM����Ï�|S��<Nɽ���˟��zD�Qv;�|+�i�������&,r�8y9��>м]7�&�6�.b�aå��K����6��cG�s��Uyz7�9�@�\���,�+C��dHj)�Gr��?P�����r�k�<�]Ҏ�a_���ߛ�8���t�R�qg��_=���JPq>@'�by�����Y�}���no¬�����T7����}y�Ff�U�1c��s�53���z�m�lGmP�g�;u0 R��jS��l �?N�=w@���T�쇷�I�q�Z1�$����ǖJҏ���Pe�Q,dHS[�DN�ϕ9�8���%`o�|��W�ҧ��qg�t�(r�_P��x�z�EA�9�ϳC:�!Y����M��(6#쬅�Y�{��6�8�B��}�:9���%���w��Xl�!��E����g��4g��ab')��ƣ��R�}��G�xLc��͒�U�S`aF�b�o�+�4㉳^�̚�:�
��D����Y<O*��]��AQ�����V:��Y��[-�Jh~�v���\��,�°qj��T@���ׄ������ٗG��%5�
�C�:a����"zu��rd��gǅ�AwG@#�"d���"X�I4RwS���CH%S E��^�
 f�4;�Y��G1A��?,;�^�j?�Wбz䥼�9ʡ���0tQӄH��z`���Ȁ�P�Z��| ����*�O7���3������"[�at�����W�?��g�	�;[vt	�EL���n�h#Ԙ�,,F�Š1�˒ձ*�[��z��C�+�,�}>��[q4ڛ[GS�5��Z�ig�ÍĴy�� ��V���,�J�F�{��!�*�u�,��UV꛸TT� �G�������bG���Y�R���C����|�;�qYZJ�,�z�w�]S�Rb�
HF�.��Z@�?�)�c�m�!p=�
~��-.�����
�+��B���(�񢒅�kI��Ba�(��ֲ�^��{|"���n	�N�<�`�8R9cs���rB��m9�4�7��@!�[�M/Kn��]��IK��MӻA=�pGPB��v`���8w��x
V�����&#���+���M�V�@�TF��N��%B��1N�dG=�0�#� �E_��B�.Aѩ�8� ��d���WCd��3�n�=P��qs��~}K�aԑ����n��8i�x!8� XY]�eh��Md�T:1f&��Y�|C�*�Lb�[$ϐ�~�2nC��ň�0�ؔ-3,�P��^�NI[}��4h�<��ͺ|�L�碆�;9�:]�HA8�ԆZq��ރ��Y�+��+�Ẅ́��t9@��iu����~��e�=�LtV�S����7�W�+uX;x�q�����Ꙣ8 e��%�6_�dl"�G��=���{/��Q���O�`�8|�!�l���?Vu���T,�}';�n�HI���;���r7B�>+}�&��?��:#�SB0�w��r<7k,�P!�����a�mt��W�^в�4���Z �h�㥶�=��(���s�fi�	�Pv��f��܋��_��t�q�H<�e�3���R���m�!*���p;9����qx1zD����$۔�`�{��=����4
����.|é�Q>�_�M8ו���@y�`7�y��	t�I|�����*�_Kdj���(���k�iY�� q����θ���):�5��Z3��3����L��[����)uM���*���L���VD�!K��V��.>��ѢN��p�h'��� ��T������;'�-����k.�B�#*co `��$�1�v� ��K>du��M��� $Z����1���D �ˑ�8�/�XS�̞uĔJ0��'W��ȴ�q)�C|^�[�	��Dw��|*���,�^�	����9���s�+w���M��"����R��d��g(~m���:Y�5[�ʀ .(`;K:�d�ꘋ�D������+ר�� ��R�OZ@>'!z<��kK�,���GA�qe�a�8���_�N�m�z(9��8���r޷L8�R����qv�_h�5b������Am�\\�X73T�7�J���R��F�]%���H��O�tN�MTr��V���h��z>C��~���_��b?�Fމ����a����~b��~�R.o��&���C��Ӝ�rDg�Iw,a��R� ���7���<��sM��,Z�z�c��%_�fO��^fl��iJR�_)��<��xH5釞�@���*>*��{�H�=[LoF��N2Nq�b��|�L���A
Tk��I� ۠R�4?��aq��:�����G�_k��)C��#��W���S��j�^��l��a��>��]*�z�P��&
E	�[ �XO� f��(;�V�N��;4>6Z��`*����z"��s⼥:�fj'�޽UB�m�q.�(����8Ձ����l�<����j�2sk�2z Q���6f��?>K�ooFB����R�F�mf��봉��4B���ehmlr��bca��9΁����Lg����|Rtn����B��
�D�������A��^Q�]���}����H�x��mt�M���x�FQz��Nlm]ML��o!m��!eL��Ϯ="��r�	��'�n�%��ϳ�5�0
��W\ȱ������?�r#�5�7�U�ݦ��U��i#��~\�Jqy��[�T�N.���-A��;Q@�:�>>��C��o=�̑�7��kIf��>�S����s���N##W����廈
<�J�p~i�96��q��/j�A0(e����r�D�3��i�>Ӹd�.���������@ 9�ֽ�&�{]C��GU��)a2!�<@�o��*����\�E��I��qu&6���1E�K\�
� �^�>��}��]X�u�2�3�����x˰��[�b���a]"��p֝�o�����ǚ��Iiv٭�1�Nd�H�r�S�v"*]4X1�e�lN5P��k�ژx��Ȝ���H�oRB���������N��Φ�ͯ��:剸߃Z�`W�՘&����q �+=)����&�n:n���t@a��9�IM5�&W����䩣�.�����1��+����	���<0��<���_�<��l���SCs���4o�
�D;�W�@-O�u��&G <�$��Q�@���r�Y m��%��.oK5�Z��4A��"&�T�Ԍ���k���ӎ���z�:)ع랭4a��Fd��rYRܘ��Y�%�� ��:Jk��-�KŽVCX�pu��i��ڄ"����k��N�f0v�c+rA��wb����B��Zm�*���=f���Z����"w�Ŗ��~WjHV�1�b�6�[r;Ć����k�S�.긂���	Q0�[�/�M�H&4q�  L��ǐyrOC��W.q��Xty�~���+2e��������
����;��6�P/�ݻ�8x�$�N�v�ko&G�sG(rY�ۣAx�3�&D ��̂%dl8s6,��W���� �����4(�ޢ�����+�E2
m̯��3��2�������*����GD�U��Ή���96��ȫ�����x���m��$�3�w�5�˪�a�h �#����U��۶¶`vQ~�����ӹ0�})y��H��1��X��)��J,Ӟ9��+�2E��z����
 �T������9h�;�j����)p�S��U�h�z�.��h����Rn��I��;�&ϮɜSl�W&c�����k&I���44�3b�T��yX�V��TR��� z
�>��JX�!d��L x.�2n���H>3�gD�yhy��~A�)4= mgk��0�Z�z��~��9�wqgu{�M��~c<��]�:�I���E>Y��|n�j�O��~ֹ%8;�b�����&�Y��'����6��â��5� U�C�)��'���?�+0���R'�H%�g`B8�gh�Uk��v�eH���P}҆$���P(I��$���:!�n�Oh���R7ʏ�O�0��(�
�wTo�x�^�Ơ�R|�}f��	q�<�t;��1<��Bdť�\�^�����>g���W�m���r��S�����5�T(bj�ôB��5�Y8NZ������G�,�xm\E�&�	��$��U��**_�;�2f�P���m��95@)w�9����o@�hi�As���v�ƀlr�O:7����i�����lh�*p�����.?Fx��뀡ƫ����jf�|L�$�:x�	�rK�Xɬ���i���I�� 9�jŬ5^��L2�X�(^_��;��3�QGZ���$u�ϙ\�o�b��M�(n�K�;�B7�k�1�E��0�J��ٲ�=5��a�:١c������e���~�Z�ES���V��?�_�i*���ж���x�N|��m�BK�Z�%�� ��J���(�DW�LL)�%i ӿz_���z��"�nl��DyJ�|C-��Ҁ���в�qy�8����Vv+ޟ5�N��Кxe����SU�).w@t��ٍ`To��POI({�i.���Z��ά��(�֢�>*����']�9�h��R=���e|_�����D��*a�����V�Q3�{��>M;[h}��tq8�&|�|o$�e����OvL�T*�uB��s�	k���g�*G���2���sH9@��x��^:�U�n`g���@�v�2���OWD9��/twΉ��"]�4.WS�:A��"*j��C���&��1��+�ǅ�-5��E�:[�.gu��͙Eu{�n��9�� Z�����W[v30���m��u,����� }�C�!�Q��p�&�鹌-�V�%��-�̣W���������Z���\�`[>1����Y�^�u�/Y^��H�[��	:�\E��>UU�qG��t���w���!|R��U�~�����/ؒ���Z�j�$H ��^�|�$�)��i�(�h!�C7Q�_�u_6.��wvt���ǀ�ZXx����N�����	�J��r��Upxw��$���<����`@�����T�:a0ſ&�W�z#嘳n��I�{���/�my���K�}���o�����7���oe�E�.<oY�ej���Ϙ�6�E��N�P�>��":n _˿Pw�=�-gC����*LT�y��=��.?�I�#7ƄNy�qA��	�?jqc�9�=�棭s��E$ԟ�E��x����HǏ��;�f��ֲ�6��Fp8���GZ@�n�uزK�\{J�%�SB��n��� ��,�ڞ���E;;��v�pu���%����9*D �0�~JN@\X[&hEg�%IS`b���l�m�ݘ��<
@����om��jJ4���K+�Ϛh���ڄfC��	V]�C��)��c�e��R�����)�͈i$* �� uΔw���,L��2a�"aH"��n��ΥV�b�����L�8?���w@ jH��rtX�H ����K���F�aJ��7Q�W���+�nR������CR(K/(��J��N�W��P�?�R� �	���2���������Da��mN of<����m����G�z?�òVhC���:(�`@��1�K���Pw��sz�P�ǪV�ɽ�`��;.B�G4V_K�����Z~��_���	�	.{����ݨE��3��
:�5�y��xZ�o��D���"����GD%�ڟ�w�V���N]FL�ԩ���v�h�	$�_�}��>��O����s�yةfnU����m�G##8����_������/r��iV�1'R���Ҩ���M�ԖjR�V6�L~M4���/�k�t�<��>wyr���:Ȋ�bj�G����,<�F)�
�8&�>vC<�H�v�4���,��y�!X�y[��	K?�ڪb���$z͋�����pl����G@k$W�P��i>�����rp��P��vQѿ�~Z���2��)��	p��]`y�����^"�!ގ���fe��`�� aY��P�����Š(10�����\a�	T�M|du^��4��y+_���ODP-�73��z+�9�
��ٱ%�!�����g�(v���{O?��	R?a�͞:#�,�F��KBG�m�nF���7���j���.��G�~�$0Y���]�2�Y��h�sݨXl���P�a����l�P�5V���g�'�VRZ��:Iax�	Ed�}��a��9������{ �nٟ�P`���q,>�� yz��z�����Cz��w�����g{|H�H|�����u"rPAl���*�ǎ�}�˖�?�9����o\f���W`
� �U��oX��v�8�0��S��v�`��KB{!>A���鈟��ׅ���ޞ1tsM��RwY�3�x��qr�Uza�$F�f��_���ܤ�^�x~�i��[%�_1fj:��"HՏ�l�'{�WH��M�#(��#���\ƊH|v\ 2�UЄ7S0=�J�'#��=����a�Q��
�����ŹT���}�4����qg���Ȩ��]Uy���GT��U�5��S&@cn��{Y^i�yH݆��;$0@����gG!����%�\yBe\���؈y���oλ>��ql[�"]u���)�.?�L�8���W�PT\X�ԼLhO
�s2�\���+12g���#l!ij|{��U;�U��m�˵TD�����zmZ�n��[�}��3VLNB����p�D�@1��3��$
�_:rc7�?���@3�O��,�X9�b���RDnԚ���# `=0o� �=��'t��ap,���.�ma�I-��f0+h�hP�mQf�'t��&����_Nc�<��D���xC������]C߭f����%�i��?8�����yR�S�Xbè~[/o=D)"�H&����7fS7���èUĴ�ټ�S�bi��C�di|����zii����:,]�R��M�z���Ƚ���2 ��70O�X��a|f[0^�2u��,�G,,�]v���ߙY�1*c	X����v� �Qxs^���>^s lkR��@�5�
A2K�m�E1]�^J4�_
���h��&�l�}ZyO2�:�M��g�pWo�5N4�ί݌R�W�����M\��qwX�{�Ө�Hd�dR'��+0�S�����2���.s���2z��K�;�${  �����e�#R��W��$��xj𪬵]<1N<��Tl�1O�K1���U��ID��O�(��_�^�̦;��"k|�:ٹ1���䤴S�}T1�(؈�\_;L;��5�u��.i��5!*��L%�����G	�Q<Uq^�uLG�X~���D����U��C[��|[^�����4E4�U��u���\��q?��,�M���<�a��$�ٮ�P	h��dq�=j�ﶇ(b�g�n��b�B��4�{���1R�v�q��=z*�osu33נ�������1}.S�Y��2�R�	�OԝhA�K{��[!�j)�l:�s�q��gE�A�r��y��Z�Pu^���F�$���b���}4T����fe�Q <�I�ʮ[�I�ي&e��qk��'�m��������QL�VR�A��Ӗ���dzO������P����6K�.��FI7��y$��>� &�D�a�yR,���U5�e�Muv�AX�q�#���|[��]kp)���Fg��^�6��X��B��T�F��>��ې�s�׍Y�\ko�����y�%k(��a���w�)����h��)��Zd�M�����Hi8V��Y�\�~.슺����^�n��ڿwu�]���L���A6W�X�Я� Q�,����x�I����j>P�<����Z,z[�
c}|K��S6�8�R��x�G�䃳K+�[]<�5�K��
�P��qXqY�igj��n����Tf,��������>x�{�RzVT��6�;j&�0�pjj9X�Eq�u���**�w7U��4*�O��Ɏ�Y1��1����
]}��n_�P.��QϺ98eU�p�/:��������ؖ�wW��C�%���~��a}�i
-�����@t�b��OE��u'���N����%x����䍡p�!�(hҞ.u\�� �5�Cs�~�Ø&��LH������3o�#i�mo��u��$��pR&�í��B��ۅ8��M�7Vb �U � �7r'�W'F�e�o�D5����>K�I�Vq��5W���V.ك�_G�8�o���L���;��,�����4���sl��ҫƋ��_�t�1����:���I�8�(�������Y�C^)�&�v��s�L��<�e0%�U;ޝR(vWONp��T`#,��������R!��1tߛB�zA��w��˼�7�����`�/��ڹ�i5�hF�@:�����u�BP#�ZMI[���]�M3jQU9t�=ߧژl���v�Gu
�S�D��ξ�ڻv20R�����Ҭ"��f>�ThqH������İ��z��s���ɘu+��!���/Bi�ݛU��rV)W.���]׌^/���[��T!�_>���WЯ���I���y��SRhAk��sd��&���KQ^�`�!x��Z`�.��rO�؏���Z�,���PB֞\Řެ��%��T$#��$9��!<F��)����)"� �*	��� � `1�M%�f��ùe�r�S�ݽc@YD8�CmJ�)l��R�>��1�B��r����P��l�����ӹ�&�?1F�?�O�dD���
�`�jG6��4�}'�KI�5�Ak�sf4�W����P���\CM�Q��ʈ5wC~]�I�Z���v�߀v�0c�@�w�gb�̏�_��:�3<u��zg�*W�^d��:���b�6>E|����q�#蕧q��\������p��>��zt��8�6�T�M� 9��ֈ�u,��Sr6ù�;֮��s�G1j&�Փ4״JN� tH�8d�	fW�R���uE(n�=�C��p1j��"A��h��<��z]�%'hU2�}��\���][L�-4IU�S���9�|�(�!W2��1�``�Y�N�%����+�T���.&��`��S߉�0~o�Q������'��tb�pm$|�$�!y	��{��Q|�<�	����H5v�N�ptKF��/C� 
b8��ڜ���|+<!Z�x͛,�He�g��T�3�u/*hvkn��FϹ��#m�:���~^�gt��pw���|ryw��{	�x��8"���~��ʊ	���9���5;{:b��>����J&� �H�2�X�2I�/��~s�@[`.P�8���0��2�)v�Eb�������wFk��ua/{�ή�Z�����&������9s�q7؟�i���/ğ�C�u8>�3�P��r�4��h2^� V|R;-���B�"�}Z��=���
��2݀|�k^y���%�5yh��vs���hAMWQNAe��o�1���L�U��<F�4��L�*��¤q�IYt2��5XSW�בu��'ة�\2�O3C��_&g����e��Q�J8`�4�sX[۴b��S����E�k��v�+�m��0���1��MGڳA�%/��~
-���D�cr��Ug�@�Dg�_3�C�_w���uK���P�*52�J���p��H����DV>N�A�M�L��vKU"z�Z{{��jb�����|T���/& ����{����=�;���	�G(B,���� 7����EOT l��� ���u,�i��Y齳%��ήtՃ�eO��������1J�Q�]�Ժ8�F��v_��K1>hE��1���m����K
�������m�%//[�Y5j�}5��Ҽn��J{)�7��3'���H-4����)��??3)��3�C�D-�'���oN}$��wm��.��;6�RA�t�w\CG����a���yc�J)�D�������G�����;
����^
���H#ϣ�����H���l��+㝨��S����5�n���xt�h�35��X��+Ȓ�zxs:g??P�Th|j+?����T��$��h2b�nB���ظIM�br��*Q�(�}��0����0d����LKВ��^BP�?L6Cӥ� �������9���p�'���wa��-�|V��m]��2)�j�$ÅH7c)fS���e$�6��t�V�L�o���+[٨NBW󻮚8��PLc��������Ā�])�w¤�t��+Z'���b�*������u�@|��Z�J��fg�M픧>Şk`��o��`�ڱ9�T�=	~�o�3.;�a�:ܻ䮽�ߜ����k��?�J�YQ,ֺ/Wֶ���&���$R�͟��;\�$v?ċ�s�:ǳ������`��Nߝ����'�[cN�d����^�Z"KS��D��_r��{�7�K+���bΧ������ꪃ��M��R�U�U��ti��%���EoAX�ɏ�T�[-��q.PZ�/�uQRɋ�
�:[��ǏI�*��G·�)g�z4���sz1Sk�{UX�߷u�T+娼.��|o<��� � D}�S�z�_8��6E�I����hH:��v�Ár���L
��y�De��;���ԣ�*6�tqo@�a^��TN��Ρ�(c�=��O��B��X�1b�%�N���'R�i뢜���;�7c����.ۮ���ze0�p=^0NK�;m�Rݻ��&� ��r��a��`���~�?��y��Op*�5 �d��Q��\�L�}�;��"�ߋ;K���vL�rj�1C�+�n�P)L@9`��
����L�����O�k��9!�=�����������~��Fy�d��4�sdwO%�/r�~��@�^&^Ѳ٨�S�pz}�"	r�uPjg�v�'k0Hѓ`E˫E�����]�T���Z����6��ٸZ'�t*�,gx�P���W���'�"�~-m���p��8=	�vɨV�gV�S`�ķ��+-��@�Wi�yG�rY�%�T�/*1J����&!���!�N�^j|��B�Ҍ�7��B����5��4o�	�Ju���C�1}��-�<�����)��a���n���;B��g���tZ�{�]���J�7���b�0?�V1ޙ�23��`�dLm��S�1�+w�I��Łv�Υ�����#Dz.'�8�A,��8Ғ7'D�z!�#�F��N���$pW�4m�}P�T�b646�=r%��Z�t��DyP����x~{kR��m;�9�f����&�܅j��=�v����������wu��	�����v@@��@��m�6�`G�K�^����⅓��-�>���'9����LV������Kz�9���*Ma�D��!���n�28��M�<��m�q������Dօ��_9$,��J�T�3a ��Rk���
�S�w��(PC\�8L�_G�-"O��;��to��X�>Y`�\(c�J+�&���V��>�43%�!]j�q�	z+Z@������b!~</�8'�kFe3��K��$���j4O��s�u;Ԉ����L�f����v&�U,�Wתoo���
�`�wxY��ب4���~�8��}j���8ʔ��e���"�^�R�KʡE��\�����?�S�������PeƠ������;�q|��;�rL��c����.}�ey
�s~0K���bK��pi����R��sh��)��a��3r�*B��:S�j�ԄC��Q7k�l�d$���Ǉ~^�������.^e�[��1���?�~^���$מ�����Xgt�Ȓ!��w%EŬ��l�Ě��>5'��W3
d��W��魋���K�:]6	��*8��ǿ�gb�z��,\���-�ҹ�=�Yo1�X �5̍o�qB�S�gJ��-c�W&N�גH��˹�XD!�[E;�4z�
Q-{	<����d�p	��z;ݐ}��Ц�ҡ�}F��*�G����"|�9-!���Q�yCy�/�>q"�A�⿺M�����y��z�N���d/�9�"�K"lvZ�zf5W��_v[{YYq��s�[Өʶ�G�7�ޢ�ۑ{���xti���4�CIca�5��[pI&vx���6>j�Q���0��@2z�E5_�0.��7jF��v~�an��"�W�̞��8����_���}j6z댃��h�S��՜���Yz4&կ���~,��E!�8��ޭ��9O�ϼQ���=��_�TL,� �Ct�.����|�H%�N;��x��C����a�M�1DW�i��[/t��jڏ-�� �c�:����� ��;�i���fa}r��M	�$��r�l&:���A��t�qs�[��z�Z	�ʶ���kݿC�[-��b�֦�<����6x:������<�1OyNb#c��#���E�k��{��������eJLu�%��v��pT�M>��!a��{�z N���T��?{:*we�9��f(��8�o�zz3)UNp-��<7�G��(�C���z��V��
j��"���WX���'�&=R���4g�Vi{4�;gv�Olāa��J���WZ���������{�1Е2����V���4@�Q�A�����Q�
�&9i�󫐃���>���q�`�8)7g��n���u�p=6Z�Wq���NV��%�a:}��6����9��s�T3M<^Z���IFEmĢ�~c0x���!=�#���
��|I{����%�;�>?=7���V��]����~�+o��v���DA��w|�ݢ��D��j=����N�u�DC��>��_�S[~%��PZ�ygmo�J�>����9g��X�Fb���0��3�h��J�ʠQ���ֺ%P��>kDM�qX~���S)���Nq���~� v��G��6�-�1Q0(���* C�֏�g��ykQ����
Pu6Pz��.= )��}��sΊM^t���*O�exv�f�5oC�=�z�r*���ښ�Zn��3k�p�>C<�����y����eM�/  ك�����r �6j8?=n*�v�3���舺���H�������)'��u�4�V��6*���gOH�0�~ �]�\�`�Q����nn!�t?�>�lQ��-�h��i��ǧ�(`L� ����6��~�3�Wz?��߷Ac��|V���K��f|8�=m�.�°�H=O�b�]����Q)������Qp7Y��l�l��PV���N��"�&�x�|��\�բl ����z��K�,"w9�E�An����6�)��.:u��TD�`���jlw�s�`�5�G���K��X����効u����2źH� F$�Z�W�?