��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�O��?A~'�^�a��嘝-Q�'��"�"._��ψ:��Ψ�n��.�)���73\��	9�}i��V�3�~��}���4�����፴^�F��� �Ԏ�Z/m��7��_'� �=���A5D��[e�����\F�q.�Kx��us:�;�:ǻ:�K6����������u���)5>��S9��̋�6I�˵^��;:���4�l���Vэ����t��@���O���`o�����N	�4k�q��
��#Սʌ��b�8��[�T���~.kҧ3�r�3	\a$q\i�&0���mr�mOc����ł�~�QbS��v��y��.��t=>,�sY�VS3��������l)����-�v6׹Umŗ,�*���Q]��!�[��Dv0���N�2�eo�Q�ت�Iܸm!���}���A�)��#y.��~��������Y�[N��2���3j��7iz���)�ؾi��o�T�˴I? �^gE�� |�r`�	��ͬP_�k��?Y�<ФtQ�ފ��?��q�p¹���+��w���D�Z�M��b_i9�,/�bB���L�@F���c���x~K�����~<�.��L�1�&lp1ʏ��v� ����9 ��󨚮��֮:�P6�V�A��W~�q@(�.��	��A[����G��0�?��%�f�TW��r#��/�>�D��~��@:�C@'J���0,�u�J�?N�Z�֚�(�j�3�}��p�H(�vf��ʲWHQ����3����j��w�0�T笿j d�_��T*�yh�:!�&��OoE�'�ۡޱE�k\�$|B)X;O�Ğ�K�^s5Eo���� �3�/�R�����sS"�7�$�Ђ~ϑ_Ԟ~j�٣э�S�k�G�O���� ���KF�.�r��]&<'��C������%�e��>�I#��J#�\Yc9��i�$Wb�*� P�Ku�&�COP[��������Q���[�QN��;�Tn�t�=�ŭ���@�C��y��s����- �yH��8R=��gv��?�����hYe�A�c����6#~��\x6����X�oL�=*t#�_X_��Ce��a�v��1��oi���=䣌w��X�J���×]�>���2O3�T\QK�k�q�}$#��laE�	�#EZҀ�U+����DQ�a�e�UU&�d���1���;x��bwW���[О�����S��%��jY�a9���nJ	�~�v���h8W�N�M7��%tPq�ə�f���B��S�I��ؽ�
(=jR�d5�Ѐ��ak,Km��s�2���λZ(=aAZ�9�s�A�}�����zD��Y[F��ORO����%��O���ߨw�=�N>ib��!'8<�M�ۅ�("C�m�>ؚ>�d�N�K���ӸN�!"��i��-�Mk���U�_��1na�1�,���0�}���u�=J^[�)� .��!��Q���?�j!I�4�������pF},Ϥ�T�;e��	G?�l��k������Z2�N��8�$.�À#�'��&؀�Wpt��D8��.&�fV*H	���!c�`�i~G<�C�ke(����휜}?�3剒/�05��c��N�=MdJ����`tn���9��M"1��X�>�U��J�nщ�����.J
��fx��gx���A�-�`mʖǻ�82#�%�Kg������D����4�i�Yi��/C�{mP&!(���`��]�oJ��^�>G
�� m.��?�d�[����S�������O��[D-�A@�<�;KY� �y���b�i����i3��{7�[Q�D�S��W����Ʉh�0�Gi�/���`�߄��o��]p+���D����NM��H�jk(�|�ɲ��%�ԥq*��C�iG�)X1��"�UpFDL>��R�/�N�I��B}��W[�2}PZU�G�I�"�� �W!�yL@ͷ�j}N�^Y17*��1c����C��ޡ��怒�e{RE�uh����IspO��� �zwQ����Ef1{U�`���}�@h�+�'
�� ���v-qY�c��_�� ����Z9
��1/v&�󉑠H+`1�}9eʞ�lc��ޖFU$��3 �����j6]}n��nK/O�[Ξױ|�Z=>�����K���^x�7&=�ڏи��ۂ>�oj�}��e�g�>�0��|>ef��m-����=��G��l�������Uas0��S*>/(����j��n\.�ӡ���@`�I�+���r��;2��O��!4��v��=�<+Ӟ�����}:�*���8�Z(3T|>j��9Ja�ӣK�o`6�h�de�ꢘC��Ɗ��j2���\��;m2���J�䷒�x>Cl\"��x�q�AY��jJ8>�����������9Mp!F��0��1���M�DS�D-ͤ��>{���0�����ors�!,.�ӲZ2�	r���.�2޽˰��L͔�;Nx�j"�¼o���@����F��nD���h��;��QΎ7�Q{������h�O� J@�B�د���C��6}�4���vy��L���u�GI��A�~_N(��kJ��S�K��5'�w �;��˾��#TQƒ!��5l�&O�a��4��di6sW����ĔN�-����s)�m����G��a�O���Ω�׬�J!��H	>5��ׄa�����r����s��Q�U�]��h�Х,��R{2��hS&]��"��� �p�3l�'˸D3�o��lfm�[Bmv�39�k����N�.�ҷ�OnG�v�H��R�6����L��ǟ����)^�l��>홢I�?�h>1;\�n�6������)/9�C,3�1K��1�*�n�!鵑����L���]@:u{�p���X:��v��?R>���~X�gݷ�`���0�A�
�&��/;�b�� Qf}���S�$�1��ꑣ��q�?Q'?�ZhJ����<�W�b��;����
�*�y`�?qe1�V����F����u[>q���lN٭3�䃃�֠����0�eFn/c��Jُ�f��������G�Rۭv��1�LJ��x��(���(�/4�xk!VK��æ[�&53\.w3��Eۦ2]b���&"7��ړn3��Cm��ǻ�l��a~������L��מ�0-�� L��s1�ܔq��A�3������/&�S8/�,�w0!�5��hQ��� ���X�#>evvI�A�����`]h�r2~��6_��c2�=N5��y��:�R҃u�+&FV�:s;U�S��Xu�]7��YU�(���
l���mi�|z�
����	�!�*�Y���eP�`Һ-�;�o�]��266��g��>2N�Bb����diY؊B�"n�&���a�l�N�ȿjn�"�Dn{�+R�q�5��eIA&z�t;�`�s_�%�����:g�8�:3b�d�0��w�AY�����ԧxx=둪Ӷ(,|�eD���>Wzk�?`zn�A.u���� �_�tF�Av�2��-d��Q�v�R�|�����5��>;��>�@@��U���H��E��3:}7aR6��u4����ʑ��ؽa�~T	()z.Ti���D��&LQB;{ x���F\��J���k����Dv������ʐ8)����R3��8;���	poA���g�������q��=��s�X����m_GW&2��@�H� {h_?z�����Fh�;��q6fų����猊M�Bhbџ���yPeƢ~�ϲ��V���z�9�f�10!�q�	�ab�v�S����K&��y�ۮ��X1��fo��.�����B���R�h��!X�����;�X�Z&�̾>/Q��2tlK���5�+�L�%�t�f���������B��Dq�����<e4����הS�C���v�]GK5y��+YE�E2�ϲ����`�.~B2Jʞ�?s6e�j���3������n���sۈ�N�F�Q*n�%H���!k�Z;��l&Z�)_+D.tn�+=�j9�uT�:*8�؋a��.�R���H�!����_�XA ��Ma��yhܱۘ�C�@��73�V�fN�r
�;���|�c=t�s/yxu�i��S�<2Ħ&��4]?S�D��Cz�� RkW�%S�����.T°04@z�%�'t2m��1&"NR���3�f�8X|�٬�=�m͠�*lXd�<��d<d�f�Lq�� so&�L��)�6N}���`#�I��g�a�ˠ���7��t�}o�&~r�Nny;��H{��������-���j%l��*}��ǎ����H7��Z�u���"^G��6Σ�װ/�޷�#B��d~!�)է#E�osf$ܒs���3�w��ۢN����ɭz�/b-Ow��B <��y����e����q���R\�����U�	I+p�t3Xi3��[U�p���6x�(�nu�O�@3[,d>|ivg;����$��.y�
�����ҠW�@��[U��)��wϮ=�(�����kO]�	8�bC�{���J�6�ٽ��)�(f��`���p��.� ~�n�
�T�6sEe%脕%x ME%)��J�^'a��B�4
��B�u�U�Ќ���&y(呮,8quz��y9d�xpExw�2!�mB.���Љ�gO