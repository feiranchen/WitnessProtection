��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�5ߣS
ؓ%�v�~p�o�B͋n���n>_g�\��ǘ�'�m�!��ys���[�� @��B�h��c�����m�TJ/�OL�'��c��	�#�N�.zX�K��%C�K�Y�_u�R�K�B=z��i������^�;�
���)���c�I�f�FW���*zŊ������h�8� ��0��Pq<�o����},oۨ��-�� 0�=�DO>3���T�Y��ZPQXv�ibo�k.�܇�xH�E��,��Μ�+�1���l$��\��p�P��>�L�{��: x��L�,���WH����^�i(/�!b�rĹfs�q�AĽ��ޅv���s�!��d"nS���C}E�u�^�|�����aFin��7[������q�A�r�H����N�!����x"]+��L8�#wG!0s�SJyRս4G����:*7?��_���� ���Q����,�:�Qj?��:܀߬�>�h^�oK�$�Ei�j>�M,�f_�*�Wvͷi�4
Iqi7j*��e��T��M�3�8!��ɔ�1�lQ�e*�5q@c���}���@��8�j����*�g���h�E�q������ ��;�}|��2����*����/Wp񠊩�d8�-	����l�.L�G�T�`��۹3t �":���s����i!������k��������3�.�&��+�~^y�[D��|j͠	�+�z����A�c��߸���������~VT����h�B Թ�Կ��B�"�Q�ov>5���Wbc�Q�KH��AT�A^�b��r0�?&�t B`ө���o!P~�`���)/n
�_/�nb<?Yjć㡯�Ĳ���_������:���Y�2$J-�^���-�`9��5wN��*�6qsq�>�$���P�6
�0q,�Z�G�N!a�au5e�](di��ba����<�̥xM�Z�������w�U/$J�y��UG�n<</RVCUw.�>�6�Գ����@�&�膟��{\��-���cd]=��EH�Ua��̂m�$�`��ƧI����~be�}	2�j��aG fs��I�!g&�.�q��6ǹT}ݳ����G��Y��\$�鈞.|M`���IY�ʩ�kA�/��"����,��g�ϔh+oL��<�i���8�i��J竽��`os1�w��\%�l	����Moc.���H��������O�5~ 	1��!.޲Fg:�?�E�CҢ��>I�0��zZ��t�'qiBĤ�����@��W���ӷ���8�?���
�x�<��ϵ��7�Iı���[{g�M��H�P\6�%�`!_���2h��y�r�Z2NJ�b������U�dk�":R��A7ՆB���X����c9�mN=�C�>�XXni��d��(����#�x�|p��Idp�����C�a��y@� F�����&l	H�fx(q���/�9ŕ+m@�����gѹ��V�WKԱG�R�oV����%�m�Ñ.��5��n�奰>o�h�ߊu)�� �����d���V��<�ۛZ
#�?1clo4�`3�ߑ̧l֥�¬�����S|`�{s͹\q�����CLj�:�yl$L�sZ5/��f��@%���OD�h�9� {�Ɔv�P�M�͉F�i�4���������^y�}N�����G
3Ra���s8+b���E_̜��Cք���S��Y^�I8#� I&tX�$k�������ۤ���b[�)1ˈ�xB��I��-��x�[�b��V��,<��E�dsb0i���{o[0D��")�4�z3�b�)�N���q����8B�kw���Y�H�F'�A�5b ������n��hpK��*�[pp�L��I�|��E
�]��#�Ɠ%��	?��f|��V���� -����-uU2w������=���B+�z\�,�b#	_�7�s�dS�$d\*� ���z��MӟK�{^����'��j�[���- �0'�c�*�%������@˨i�ي[/es#M{�l� "U6�vc�G��[fZ\01��!�\���D7<����ڗ��$�Bܪ�%�NF	-F�dm{��we����VsD)�������ּ��uc��#^�h��PV�@ߍxM��B~;)d/4ͅ�e�~7c4�� ̨��Yjj⊸��`x�H��)O�ْ�d�>{X����	� �n8��~��~��k�÷���#��4+�X�j���i���A|M唅x;�F��l�	#���?N���:�qt��I�{CM�m[��0z1�,�@���̀�ƃMg蓑}�e�)oj��
�y.KF��V�}p,��G�CbR���s0mcˍ�5�Xw��N��i_��xΊ�S4,T@zB�#a�!���m~��f�������w�Z�:E~�u77-i�,jE�o*PW#!����-�)���	ms)�}棋)@�m�7��%b�ak*(���,G�A0kV�OP�
����̟�f|E��u��- ��2b��fF�ֿ#���}Na(�w�'��j;=ŚxZډ>N�q�#�hK�%|����=�/cK���:dj�!���M*9��y��H:Z����'ҍ}2�M�2,j*���-i"�T�+ |��^Jc6�ld$H�`d�<����,����^�ѡ=���5�d}Hk\�m���A)P#��,Z�Ne@q�_�Z0�
���z�qf�����){bU��J��/�ZY�҅[�{^B3+4��,�:��! V�Ƥ:>�Ƞ�x��թ�_��@��x0)Y�9-�Ip�r7?Ǹ'|R�B����;�#�':�r�l�tQ�7&N;T3�q)��J�9j|z�\g�1�y">FY"Z?�2�4�a��f��5��+�o���ݪuyz������"�k���rk	��dQ���#u�F����&��Z�����%Na\���?�&}A��3?z9��yy6MO�H0Z�����NǾR�=e�[f��O��O6�tg�Z�Z6n�ǓM�[����d��[A�#.q�1�N��sCW�9,5?���*tx�ٞl(�u��dǸv���n�`�݃;{�˭"u�w(iʊ"%Ҵ�d�<�h�x�p0��y4�(.�w�թ��;D7�ܠ8yѦ`H%���d��E�TQ�GM/����z1�eQ�cU�I�9.]�v#��p����S!0�)SA�v&�-XZ�ie�`��|2��]O���7(H�-$�n�;'�"���&Sx�=��q��]1��� v qB$��s�(_L����S�����F��/���7H�k��X9:J,���c��郇���%�4�~'L��Qɍ4Ssn�z6y(��o�����h	��y�G�@�f�ë����rT���(�:��r�&vۓ�� w���𚛳����lt�-�����-q���_�3��I��K�F9��!�D?���F"���eg7�{��l�̩���8�V�I<啨u�-��'�^ iu綵r�l	˔��R-�n����s��� ���{�"a��m3������n��p�K�ء��@S�.�I�Ą\4`��l���V�1��-+R�f�V�|VI1�ʍ`��zX{G�m��o�>��J���w�Cd6�����h��ߛa���z�6�o��'Od��<ګQ7����9�00�V���}8t/#D��\a�uq&?"�D2L�,/�x�B�K�V����H����R����e;��b��h1̛v�sxB��89�	#�A(�[��31�Epj�~P�i%�Da�r�O�<&J�U���c��[%~B9� o�1��$����熂�G}�٪QkQ6�_������*f�M\�����߲0�>��z_�ZX��
~$�����K�D\�C�DHK��R�hat6�čc����h:�7��o���J�����$Txd4?:[�Z�4nG�Ht�����H��_�	�������5�|��4c�"��&}}M'�Hߎ��d9ut���w>����Pf�g��ln���B�@�����c�B�3/�~�輗��g���P�U]��;��K��#��2-�C�qT�����l=�0�?%�}JU�	:vpU�]�O�m���Y\T>!-��͕�ߍ��k;�����6Za�*��U����!VYzI��K-Q�����Bˏ����Hj&�,�Х��K�ib$�ɱh� Л��1���$A�q����e�jGW`�'`�ZE�ϲX�,�Б�~s�l_�~L�y԰}��8��r��b��-�Z/��'C黻݅7��{=��=�c˂�z��,�%�g���O~7I��Ô���6=N'�}�@����~)Pa<9�
/��;2���,�VgX6��T,
h��Tn���:�O�'l���9/��Y~����p��u=r��ڈ�ɷ^�D�UG��^&��ab��N�3��z��r�M\Ӑu=�ɒ�X������t°��x}%��^a���f|��^�g;%�G��g��Q���}7A�7{�Q��҃�]�,'��SH�� ��=��lȂW�6)��J{��l+l���9���������	���o�׉-�� ��ؠ.���`���A:�����<�� �>{�)�C���e�W�ٕ|��S�������3Pj��1��%1D&�O;�����X��O��#f���]�W��I�dJu��M���l(u<�1߱TVk�>�1�B��ό	�� 1 N��ˈ�8j�������:�~�� k��z����	���܊ZJk�TTQIB�4�_���ȅ�7J6?.j���3!����r���a��@E��B)�(�������~)<I gWG�2"�NӱH��U/���`(��x7k
��G�w�H(9)�c\DݺKr��^S��b��L���TH� 3���խw	W��聆�Ni���f��aO�(��7W~i�M7B�s,k)�Li�s�z��5�y9���m� A;��AFs?���w�7%ݠM*�������y�[gկ`�fo�]���S��Y�|��:��됟eu�����Q�,}n�;�"-D.�M_y�}�[�<��D�TXHaE�_`�@�l��- '�i.V[�i�1ȴ�v�hM�pku�!�8��iEu�K�W�Aڐ���[�Y�S@(t��@]ۦ��%��SԱc���O��eiͻb&�>�m���R�gi�k�<���u�,�x�h�[fVI���L!۝�{
c*y���wy_"8�����~�l짜=>��� 6��d��Ѹ�a,������&>-��ˏoݫ^PT9id�]�$R)%���Y*[�@]�Rl��:@��C������IstY�zV�Fď�mq�
2ݮ%t1���)�\�-E,��@&�3X����?*[��Q����A�'e;S3�^�Qw��Pm���]J���	rV����M��5�l�#jtnK�V�sJ[��d^K���Y�^?'՚����׭LS�wB`7���i��GjU]�[,	>G�W��>����9s�\�{�.�_3Wy�j����̑TZ=8�^�h�:��������9L�+I��m���"߼��f�]�*�	@�i
71#;d��0��fl@"�/	���3�oS��_��9)��؈�s��S�~
��u�qUo.�b�p5U/Ͻ �����=fEw�Ȱp��� ���5��Q;bf�9R&C���s7�����O�FX�ykob�3�W��r9�J�0�ŝ�����I=-���Z��X6���L�A��8�إ��λ�8D쑦����q7��)q�Im�
�q�D����!~�>�C)���w*�G]<�̈́��<K�^t-�E�C;���
���U�jz���]2��JXW���1�J�;���w� N��15ńc��i���:��VD�{����l} �ƚZ��1Dn���x��-+m��ǔ?��.8��)R�O�EK?�Qn����lds0���6l��w�ՙj.�|K����'S�V���Ȅ�PgU\�i�j����";)S�-H�r�`]b�{��,�8eǢt�h��)v˥�=a�Q�xஶ��ߠ�!�8�Ix��f�m���7���� t���Lǃ�p�վ���F�r-��XVt}��b#��I�>D5��(����Җ���l aFn�L��ac�!�3zM�l�)C2���g�Y�96½�|�a
*�a�k��?%��s�wy@�=��;��F�����H�^�y�8������C�:�X�j���C*�T	��o���0#��X��@i�!����4@n���$Ut���~����+{�
��["������.|��[M�����^υ�u9Ą�ڒ;=���=�<��F.�@N����P��yZ�=�}|jB����h����e~ ��-��y]��{�M�T89�q�Y����<�LI���
9b�@������y�Tf���xF����6i)f�MNE�&W�6o
P��E/X_��r�i᳁ǩ��N�p�<���k�R^�63��8+�AS�D��&,/1"�C����KE���ƞ] �Fhe	8jZ����jҦ�Ɔ�B��/r�9��|��s.8�s�鮎'/I5�2̽2ڰ�����I��<����K�����[����x��\u,yZ��z�cv>�[7�F���BT�5�@���J���M���]��>���%l L�wP�.^�%��q�EH^,����_�h�P��G?Nj��Xc�̖V�&��+�����h�[�o��Q�F�	(��a�Z�
�$����/��z��R�(I^%�Tdn � !H�d�y%r˹�7���4�5Ra^s-���ʩ��-���x�	�W�����n����vaI�Ќ�}.r);�~�V�����r�0#��%�F� ��/N����J�v��k�DG��X�l��>��\<��3u�X��$�R��`���۱�(�A�7��Q�4����Z��.;�Z�7�^#���;��[��<mm��A��l+Hcm<GB��KEUR�>^,ә�`x��MХ� +����0"��{3��Q�W42�h��-�����������}מ�*^$�>W�-���}���FM[�����Ҭ����e��,�1����r>��t�i�t����Uё+��|ɍ�u��s�G���+���I���wvd�pDѥ�V<X�p7�
3�A���Y�Pt����1ٔ*�G�VO*1'��Rsw+	�E��-���%�3a��Î�ӰEW� 1K�c¨# �&� m��X ����~ C�ׅ½c�Z_GoD�����^���!�s�wO���� �O�C?��X͖oqF[ �o`��?�'�ʩ�ђ��s���Ō�LWD��#"�+(ۂ:�ZM�:��T��/�{|U	q�PH�?�Q�E%y����)�#���Dh9�Z����IVF���䕺:\6.�	�o	`��EUݨ�$��N���gtit�/ʩS��~��� ���\
P~S�۴Q�e�"�5�!5H�3U��,k	������p2��g��� ��PR�e!3x�?��d�Ñ�����q��v9��:��)�V�'�d��<d�:G�'<�Fm�G�<����J���_�{iF�e4sxu)e�˶�U�����:l��5);���6��a�e��������!4��H�	w?�+��=H����#�>���K�G�B����I�%�lg}��Bԛ���nipoה�(�A�n��A���F�wl���v����h�?M�7�S�'f:�X�c�����2��jQ�����It��mi ���?Ȧs{����OԹ��k鉳�ĥ�n�~�L�s�QҰ�fQ�M�_�LtD�	es%�1��*��'S���3X�����~�s�5���4���YBs��V�Ȝ	cZr�d$>��=r���GP����_��&oI�^?������7O�u|Ym������� �.�|��/I���8����58 |�� )ѱ�h B��;�+ ���^����F|~��1�v�UF���A^��Cm�'��˲�D~�@�c��	�6��z���(��B4�)�DxM}&���t(�)C��C��ֶ��Im��!}�cLˑ�b�K��HK���Jy�mW�����Q-�ș��Hh���]�& ��=��>�k�����n=2���G<h"2�A4C,�Ϊq�j�.l!�Ho�)�H��͑�p;�3>�����5�Da��A,_�U�B��s@��s�>g6���Β��tm�Bq-�tC*�:���<���cO>]7@Je,~A	"D�g��P�M�}��G�89��{��`�V,��5!�
!�ξ��:Z�(���Vުƞ��h�O1��C�C$��W�#���+r
��_*��Y��-yA[--�'N�_�!�"�6��e��	����u����w� tfw���|�K5?"��J����H��`x�i�&ox��u�]ڤ͖~s�������^ⷙ�Kk=�.C���I{�l�_����n*&	}�8��t�ϊԉ2�1�A�<��#AGV¨�j�="�����:ݖ� p����ve=��(o:^Ed�p�����CЏ�F�w��7���Ԭ`r��	)��������Y:D����x"3�	�$�S��| e�sUt��;�(��sR��*��Xr��u�Cv���H��&. �+[�l�>��5FLqc�3q��T4��"i�|la�	�Q,;�ۧQb&�����;-�o����UkϞ��R�l!\~��w�t�|ڄ5�ƽ�+����<�?�_ޠ-lKD ���������%0[�ΝB��վ?]� WhSnL���Ī[Bی?/ь`����R��Y0[Y��X�T�a�CM@���'��։� �r̼���GoO��������H�a���gg�N/ٓ�fA��1Rϊ���D����SU̗23!�!x�mp�3�|M�f_�]eR����@�v ������p��������?T�]S�!�ث)������K�T��|޺�7]Oy�b�F�\_vp"Q-}bFPu�\{H&�)�#8����s7Ɏ��[6��J�lkϜs{+);|׸d�
���t�oS��NV<^A��֏������+U�|�FA�fKע~`��P��@n/�(V�yG��R�7-l�OV�.�7/)6���\=�^dc{5E༬�,��vC e�s�f |��
1�d���\�D� ����é@����yX������&���������0����0���貋��jHoqʡ&�T�"XG���D�,`G>#
�>bHТ�LgRj�Ϩ��J�d��j�$�|�,��栋f����N��ס�ibD�eQ��nj������9ഫ�ƣ7?�pV;���_K��v��L����@qX�3�g�~� @/-��v�U9��ǫPe�y�FO�Wy�[��>5�%�>��D��ƊZS��n(�����ᠼ�=j���}�c�-��K��g�*���I���Ml���N������(]q�<i�p["��l���w:���-E\�:4�"����.�b`dDr-F����L��1�	�Ɍ�>��9<,�TSKv�M��r"A�w�
���|&^����ִ�u�ٯ� �Z��h�:�] ��b���vBW��-��nG�9(Y���ߏ����;�$R���E�l�rY���8��������x�m��J\�W��(���؇sە�(�w}�ld�����g�4���{�Qa�0jDh�6��\b���Ir���%�X6�A��^S�l{�v� ��l�Ƹ�,V[ ]F7�yA_�-��ٶ��M��g�4�x����󆲗�5y>?5fYC���w���� �m�-�����B�f/+#&%]@���v&l���q����*8����	�g|Ю[ߝ_�}7eA-#"͞�+��c��ݑݫQн��[&R=!��l�,�ngi+�;�K�������=g�\qt�Y���o�֊�� ��9��u*�,}���f �֞�3]���P�@s�d笢�M6zd�.7��Z�Gu)'z:Fw���~���ﶥm]g̲r���������z�B�B���([�os� �bk��x*
���Z��6�C�OM�~Tv���^���h�\��ﳠO�� �~�m��h�%ȝ_�.�m��&��r��iv#���eL8��4Tw���T0�e�(F/�����=�)�QHGl۸�c�����:�"�)�B_Bc���v��!�)>�ξ$n�B[�H��^6%�p��Ő��%���Xj�V��0���N��ʔ�Evl���>��Df�J���TH���QHbe�'^�7"���o��;���ח/L�`�gz=�7Q��Ԅ{2v
��ਓ�-p'|����)�����4�"�����Y���e�%�
o��h$�6���������Q�,'g���B�6h'?�R��}���~��%6��/�F������10�f�6�p�D׌��'����