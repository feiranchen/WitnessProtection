��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p�l�z�����k������2w�%��G����cׂE�D��dF�����/p��g^���҃\��%�KҰ�}o�AҍXGܕ�_Ɨ32��ٟ�l�d��'���甹q�����pⰈ<�Ӟ\����c�N'�f4J�R�����*y�����9I~<'��Jzh�p���0�!����c���})󁊾�bDCN�,��L4��gQ����\&?tϏ�,����~��lXE<�������܉3+<ܥ)�v��>q�|(P:ס9p�v����rsӒOl9�,�+����(_7�@�
��| ,��שZ9�䑂	�U���x��rL�^�`>��&�GRD�Gt���F�l��j�7/o�*�|�vm\��&��/��!��f>w��|BW��h��B��l������;qE)�0�{�Eˢ}�����$F��4�$B��8ާ���Z�c=�B�jZ�;���Ѳ�z��㓉_
�3D�b��yw���Ed��[�,l�����aedc��� wI�}Nh�"���������8A�!0���@�� /r���މ����1�x��`��Ub�%�X�<�	��I-j�D�B��eBNdk�C��~U�=�]���T\��"��R1$�&Ι�4L�8.�������y��?[�[�X�%���ɦ
F�4Q���o���
慨�����0��4x�m�^m'��@F���w��
�fr�n�A�(�΅�)��#�g��wf�"l�Mu+
����������׺"�R<�2^J�x�]����V���ie[���?�UJ5�E��ra�V�,���[2�;�� �z�2�[��ZLl$���̺#JF33�1a,�������?d�&3��OAr_c&а�:]�G���}-�:��<���p��'���Y%�����R��`%h��ۀ�п���N��Y����վ(.b*A���1I�P(I�GC������0�e"����w�਴H�,_�w�`??O�şf{���_�C�jF/J�!�E[�1���+��T��]tQ���.���I��
�VL�.P�ud�h�]%Ikp��q��,:A;��k̓U���/��H��ȋ"�n6�1�t�+�*�w��W���E-̹����c��ɐ��'�]k�v^i��A��+L�USB���{p������P���(%3�QXR����sWp� �r�0#�Đ�m��_���\g��Y*�
�XoC4�k�''W���Lş}���$ϵ�(����N^��z���|��v @.���_ն�}_�KR�t��~W��ː�e;b��1^)�"�W�VÄ`&��;�Wo` ��;�P�m�~P�U�c�&�#�V�Q�}~&���(�6�&�ד� �l�t����N����+0�D�s���)��2W�5,��;�X�J��>���{����yb�֞�09
���ݙ��K�����sc���_��f��J��z��>x`��WϪ�,&[8�\w��茈&�'�!��?�xQ���X#��[Z�y��A� ��2>�C���w�ܕ���m��p�o|���ۭ�d�p��Պ=K|��2ԍ��z1\���U5hp��.�G������(��!�4��hWb��zu�Qic?6�+jdOkiTQ�ɴ� IˣBp�u�*���t��s��ƗGj��.<�A���>����U�f��ח_�ܺ:0�k$�����_oN��ݓ�J����7� ��d�h��}��[���p�� çkD{���`W�R[@�>�=7[�3����GS����eW��(�C��Y$�fS��б"=�*��z��˿��]�Gw������i��!Х�����(��'.��A��A	eaU�5�՟]#wi��O����t1�,jɂ��G4��]�U�
ߠ`yꊀO�+�5>��A)C�@��5�?J<^���%-j���Pt�'	���!���G���𣸠<�{��y �[$�xo�-��œ�%�%#,c��qf:N��<���߶f5�R�tL`H�]�	�.G��3�'�|/�}�HU֩�[HW/|�� R'�5K���oΪ)6.�Z <I϶W'�x�����,[����[َj�J�d~ɣ(/jg��Rf�_�_Qq~�Qz�i�1b�)_��EDn��s�Ho�a��N��-u��0���}��X8�\A�)NcE���*|��I��8\�L�]�h�T2��3	
�ÙVn�-KbK��v	Q���<Ba�� qObKgS���j���Ѕ�̲鐅�x��a��]��o����XdN�k��ɹ�7����l�h���G߆��f>H00ؐm�	Է�&ޢB
�4F��]߉.�AhlM�mƩ�ʡ<�{��m�������xae��&�	�KJ�ڂ�ʄ;�@�A=:��su2�_�e�[Ÿq�_����,S	���H!���R������Z&J��l�c�����M�6�4muV���r+�~�5�+�i��k���K|���Ja.qͤ6 Ҧ���j[~��}�X󾆩/���Sׅ�4˟C�E�P���?�b>�����}R��Qr25ִ��3h��<�y��?�*C�ބ�P���T-o�!=|�nZm~$gKÃ������;��Zw[��m���e5	�ڏ���t_�c��Ѷw��B���۬f�Gy�7����5<5AfD�`�T�-PfO��$�S���ŀH�!������+a�%6�1��<%&7#E��s����%G��PP-{�dz����d;5�xO�#M��=�>�O@�L��-5�l�]0$F�X� �wX~U�[��#�%^��io��{��ԇ@5���C��\r�I$�VeS�HR �3���4�^J{E5�v�=3�Z��	�8�,�Xx�K)q��m_���T][kRe��r��oI�a��D��>?�(�I�5����TmWx�l�䗏��]��
�8��{����s���+������d� w.��@}u%E��ـ�
,�8th�*{}_<��*v������:��������zX�?�'�>�W�:�Mj������-�2dg8׺�"��p��b�_�G`Z�4mv��؂�5.�<Z;	]K�H��R�K�g�U��
B�A�[��, J��#��w�����#i�R8��J�P��ʎ���4��
hV\xZ��76�Ϲ���hؒ���5�#�Fxt��d�o��;7ˈ�b7��!�' �Pð����ȶ���	'X\�zW[��].u�ҽ�g�{�fF_6��>��?"~T���j5�t�%/7�	��^X��;z��d���A��L���U��2E�@�������S�y����s	f?Hl~E�{Ad�<�&<M����lDߩ�����Ԗ�:-�,�H\�8z	�.��O���ʎ驥5�5�u.�ޱ1H:�
�8��Q�m[~Js�s$PP�^�ʮ�p3*�hHY�),(�7k�⼎��b�,M�fo��z��~5/V�$�;�y:A1�w�6��o)�A��*�4=w�,�٬�� v��m~����3��Ƕy[�������r:a�*���#c�0+sM�M�ڋ�����aqy3Gz��?���&�� ?T�	д�nH�".k�QGzD|�f��FME�#�̥"���0���K�(�M�\�y��ʏ��׵Fk�����Ls8�-�8�w��&+Z���a�Z���my3��J��׽g���|��S�'ɟ[Ҭ�䨌ˑ�Q�}�B|y�������B>�q��w��z����ﱩm���:9��������˞݀���ݞa(����#�G:���R�F�r���%,�!Z�K�id�2#2AŖ&�[��f̡wC߹ќ#R�A�zP9&�8Z��G�����֖�!��bx΁^WX�x��e P��m��I�#�.JȰ�=�_�w��*�\�`�V��K�_q�.G=���XE�͋/n�g^�^�?j���L�i����D��а�6"�o>S�b]h��۠$�M��E��ԑ*�gKs`X���~Ձ�8�3��݌@���)���3��)u�> p@t��R�������#q�m̻>�Er����ƥ��1t����Td�e/���E�T;m��^E����t���!��6�"Ϋ��}�Iqu���#�:��E9�Zd�I怀"� ���hJI,!�T��k�B����AL����uK�\�p���rZ9���z�o.�ib*��M.���:�L="�����w+
��8:�R٨a9��BU)!�=��NK�j�%��V�#�$w,����u"����Ce�~~�.���^�B���V\P�W6�EQ��w�r[z8I�"�yz�"9�ʺ�q��X�� 27-�"u�U���1��ts��Q�`&�Ԫ�����r'_A,�k����q����摻������Z���i�3�H�q��c?;QB:׆�F����\�aX��h�vPX��1=ʲ���G?���+g0��C�������٭"�b#�|����V&]�B_���:�T��S��	�
�r��m㷸(�\�;���(q �[�q�
8��$D���<H�*��o
�m�iP�.Ֆ�E����\��� �
��)�QL�o[b4cz���'m������j����^a���e���l�� d� �E(JN�����Bg���oC��@�Oh������̫�|����q�S�����{��>|k{@����� ��#������1��6��C���(��F��&)�©�ø!��7�u,�Dt<�����OC#�iT�����Υ�Џ&��	HY�3�����Ϭ����C����x�&�$����Po��D���T
�pjE�;�I�3�u�,�-ȁ��m�"x�����g?d�F,��K����:�=<����s�˷�'$]i^Q,ϫ2�7Ѝ@2d�"4V�����1'�tS�����۴+����v���X�A"��L����[�&��'=�	��4�vJ��| Ԣ�����܍�LA���;�`]2bF�쳧�<��8���\t9G����k6�u`V���W4����
���?-��"VT��N)]\����UӃ���G�l��O@x��&���e�.J���E)���K�d�P���$�m[(;Z�/�0-� 	�>|U)!������L�Lu��5�-���Y���yYѝ*��l�ɰ%�`{t����GŪ6��8�Ic��e�pLө����A���N�`G�I	�-�䆤�|��P4�uL\�n̓���Y�P�[Fd���-o8`��i8���)��W�@�A�`t�)'x���z#ƊM��_��P/Wh���ڥQ��{ sb�n��i�Xd�\s�C#�Lc��#�-��<n�zq�<��IJBY=L�����a{prZ�t^�0���	&^4����CL��� wJ����]Ԇs�V��I罘�Ú����4��	�p�e�/�A�#�S�D�<�5cdN�Ĵ����L�$X8�xC�/Y/3A����=H Y��3������p��b���ᅕ)��B5��o�4]Ĉ�\�I��z��\V�i�O�rF�\�J	N(A�d�d�)�V1����yK0���'j�^R���Ȭ�Υ��8�\��뭢�d�6Ā�ԹI��3��;SQ������ҙ�k��R���_���lB���#��P+b�� ���V�E⍦ �cT�O�W�S�D�9$t,�\��	�s��H.����.D��_�ڶW�����<�ŗwM�m1�������>��2l�/��t1�����Uf��8T�ޜz����wa�H����R� 9�!��%��>ڃJ���íN��>	��"�I��8آ����w>��C��^S�� x�dH=�`�%{����� �," @�-�RB��\:=�>W�0$}淭Ԏ��}�io�w
;��y����=^ =�ދ�,��k�{����&F�SA$�C��=Ls�n��=^T9�(���7���a��<Uv]�9%�<�g4�:
���� l�$�Kj�ɓ]�S�R�/�DU�{��u���î���H�)R+����
9��,�!��;n'nz(��~�r)�Mf+� ����
bF��y��Z��a� F��l7�b/~Sm-ӎ��F�<�ؠ�7��� ����ڽP����^� G�n�LϷ���G��u=�oh�y���`���_����͒i4�4��Qi�vc��E��i�[�\B|��W^��ezJ;%���>и �L'�¡όkC�o&�����"*b���z�`	�`wR��V��K���Uo���})���I���{��(R@���ԩjh�\QpLfG��6��g��54��������P�./����A*�3����bpM<�'�Pf �X�P�jZ����hjh�
]�/�˭ha��(X��bjD���'�5���,H�v5�/P��$1�{���O�S�a}�(!V�*��;.��KE�� �������  �����KTJkge9J])��d�3�;:}8h�(�ZK��[`ַ!�XGk�Y
�z*�+��N�Z�n� �k|��f6ї�M��R��A� tTi������Л��M�pƚ<~��w&p��\�ns��	���t���>��iS+L�濢Qm#�0�0�B��F�#�|���%̇����'ף�Ɇ�Őu�� ՄY�pj����<-]���W�vZ�A��J�q�;7�b�ø�<��Ѝ�K�oE�
��z8ZE{!�>+杄�Ebbָ��	}�r�r��v�=�Z�D�Z�ͨ�#�
-��!!Y�%%z����ǰ���Ŋb�#�4�=V��x�p6!y�y^wD���N,0F��r�D�Ϲ����4%&��Ȼ���)��&�r�.�XO"�Gi[�; �6�����h�L�9��9!X��]�������8"QU��G'���F	,��IU�3��p+tְ�#1�ף)�1�^���|�%+?�X𩟷�l����U�����*Y��l��i���>����,s%/97޼� �8���q����5��V0��� c�v"�_A@�:妈����YE\(����.TWD]{�����e��G�k�7y�q��?���O���ذ���v� ��j�!��ǻW�ԈI�e�����yQ=�Z�Fjv-8�U҂EH�os����iö(�ec��Y�o#�n����+��2�7����6��dgb����	��4ߵ#ȖHR���'���u����_�::�A$��:-�%�1m�'��c3M$��1�W�G;�QgQ�:���ݥ���5�E�Mγ>n�mHF�P�A�U��0�x�HDE�K�`�@�rǼ��uɍL��<���4��V�?R@��(���a��aː�;���j�?i4\MZz;�ͣZ�l�}��.���c}�?����'5��Iϧ~TIɊ%E��������v��д[�)��#x�VQA��������������7rL��Xۘ~��-���'�������,:���e?[s�<⪻3wq��4`�A����Uu�T�#VNi!tVb � �6���wZoZ��p�Yk�# �JdzA�����E�������<�a^|�����R���Fx���*���6s��n��=�g�?��.�>��y%}|CH�b��/\{����$��o�,�FٌA��n��7j������A����௲$������3���/-��(�:�ir�="o���ŀ�M�1X�����@Lq��?�q��:U(>?c���Snz���W�K���LvЫk����g?M�%��Cf����,�&k�1b��١>S����,�z��q͛����2��y{�ۀ����*�T83z�Ϯcßw��S#��G#ޚFi]JIH�9���-�Q�1��D�Mr�q�~%(!�(ָ��;I�LM��7TͲ�x�,{��U�ް#BsQ0_��׸b�g�i��	Ș�/�*��=>��fq�t^~�'O30ۂ�l����?�?W;ŀ���B빿�;P85s������$��>p���t���`��83�W���d酪���z�b��&b��7'��ֽ�q��ckm8|�� ��QzcHw�`$k�9���)���m=ɞ�"S��kH���l����2p�����@\�m����1�i���B��T{�j�؎Ր�kSG��u���\�0�	c��u��	�5�-6�z=��x��PGcf�)�[=w���8��Ԝ�?�uf��(�r6>_���~�%��Z� @�P�VV�:�D���������_�H@�1���F�zUa-ΐ;+Cn���m��6�]&}�0�,/��tQ~p�O���<��Z*7��y����_��0ze�����М�@gOj`�*ێ[([׉��	�E�N�9��?�-ق>Rǁ�M��݂�l�]�W4 C����(�-�V�Ge��\sIع�'K���:?I��CW��u��F���ȇ��������gGx�!�ݦߜ�O��L��$�'�h��ۮفU�W��#L�b$`RɌ���,�8Y{��h�q#�-�yW	�1�}R��&��&�NK��z��\��Ƹ�D��L=��w� ��$�z=��0f�]`α����㚁=�ԣ,��?��u��20�zE#r8߯s�sZ��8j�-��汲2Pv�����E��E�e�dKK��N܆�!'������:�x:����z�!�m��1.[wfB\p4�N5_��BtN9$3�Z`}��`ϰKh�t�	�f,�;;My׍�i�7��2�I��#E;V
���/��g��3ܸ����zt��s��k�,@�e*<�>�Q��L��f�RYEn��q��̷9z�=�2U�>����R{:m�T��KY��@�37`�;4f�SߠϚ�&n}iI�ㄣj��i����A�Y�|P`��B�78?�Ds,�;�8�;l��.�<@�>]���Ǹ40���gN>���Ĩ��e�.��(�m��Ok�Y�����7�h_d>>�I�~�u.���^��$T����-i��ф�#����̾,@7��o�3��āSs�5�	҄�O��Bk2W.�$K?ƪjm��e���^�'�Y�z�#�s0�P �~r��v'*f���J\
E���sg��$1��]����}G`r�-d�@��"���eO�����;z���pUd�:�v�_�<U)�[!�'w�y5U�RtY�2n��1:�L{�t���<� �~w{��8�n���cӬb] ��'�Z�>%7���j��p�V��n���^t��S����Z0��d�<Or��o�-�.D����}��ē0��2�}�ᯕ�2�@�g���39�I+�\�����0h���*�R+u2�`ҥ!���荄w+��\ľ���.t�ɊlUlՌN��^�"�ŵ��I΢~e����1[��EQpE� EY'1HসQҹ&_�y�:Y���錃'�3t��Č]�X��#Y<�Fg�5���t����<��t�q9M���!};]��Ň@��ޮ��*Ţ�Qs�}�*m���;��)�'k��|�^�������^��D�7N�%靊&�H���^\b��&?�t��A.��M���߆�g2�>��Abs��}86�6��IQ�XUD
L���΅�0ÍH��ψ�V �zv�Zas�]k�	��"�xy��6�l��N��/Q�:8_�9��I�}AD�"�m�� 0��`Z0M6>k�	͖�
�m;����omn@��Ni�(u����I`����}H�Xh֯]!��)suNΊAZZ�.����?wG��~�d����X�>��&Pg�TЌ^�u|��#"|�ב��<�/�|�:Nr ��v��-��	��w�̆����!��%N�R|��u/9��6V�7�d,��+� ^�I�{och@�j��I���U�NO�E\�[�,�Y�k�g?(	��O?r��!�"�{�e�]�N����Z$Z�#F�+�9&C����@(�ó��I~a��8/�ϟm��~��܉V�ȎiY��9.�\/8#H���(�	)�r�"����*Ӓ&ǿUbҊ�����dI��k?{{:�b��<�Q	>'����Z����.q��sx�I����ܾb�ݢ�Q�;Ҡ�g�`�(�,�����Ŧoi�*�7���%L��9��7c��ϼ�"�('�wزaT���6�t�cw5O���!ߴ<���3 ���vo���_��i�s��΁�gT�	D�tM�˃�YC��������1��|+|zG4��+׆>>�Oh�{�wMA�h�%�?bQ�\�����EY��B�&��}�^�YtR|�n�z'@4s��I;e^�p�N�3h�k��)��2CH�w��l�z���J��y���%��h��E��0���x8�Ai�f}f'9��G��AH�yy�dܢ�P�.���n��gl��_ԉd:Z�EiݞČL������E�����VV�D�����'.אH��љ��0l٧��Np�-�ڡ�p�~sٕ��QYpR�2��kOv��zՁ�mn�cq �ٮ��g�@w����:��FdN�sw�#�|�>���D�F|Ľ	���rN����Y�cbɎvR�����Ub���gb�W���U�M�<Z�B3�Fd��
#`�<��C+�b��tG'�Z�=�6;�3k�g?��R ���`�4�
u�&��}����jɷS�U?!�🀸�Q��%4?�*�a��Hƴ��̐�j�{�+���y���7�{��:�p�#v��r?{�1���ٕH)�mJ�C�b@�����Tjl�p��n�"қ<׋�%��g�(.̖X��K���S�Jw�mGW��Ri�Bmi�6�S�F k)v�l���-<J����z޾�M�W����7&^@�Z�� �"��0U�\_N�]�z��@��X�p�sv�wȐ�y��w�u��I z�]����Ν0>2\���:b����©
1T�W딢�F����t,į�+���8�r�x!o���@�t�Өѵ�i%�C�W=�=fW��+M�3qge�d��@�8��N�o�S׆6t����)��'�**>����0����]���e��Oj�'�
tK�\-�ܸp\�~\ӷ��W6��u��,�ȵ����}�D�6��N3�{(:�~\q��waLtbV:��=�8Gъ���A�U'�jc�� ��������pvF���%C�Œ�F�-�[@yNu0�.����1�n7v�JK^�Kv�"��$��s���F�݉�bs��4*�u{3Q<�W�b����=YM��Q'�^�<|�ʑ�����3ݑ�ϴ�\S����l�߾��F�SG�F(����=�MY=&���s���+��t�8Q��Х*N Bnt��
F$�R�Mo�����?C�͜eFgȒ����d�����H�B��g�T�K��*��A��(XdQD��c���u��1&l� �)7[_�)�����Ml��i���D�0���v�Tr���t3��l�3�R�� �T�o��J�?�hs�֞y1����7�-�P�1��G(�ZQ�����*5�����>��Υ~�*&U�=�DU�-���*�&6��oڀ���vX�H�G(n�Y����Y<��i�.*9�e~@�]N�}��VG��/嵚�`:1�S����^��P�L� �vaD��t)߁D��_�A=�^���Ly�ZrH		�a��Rv$����'��;N��Ar��i6g"u"(penO��
�&A�,(����A�!�k�i�3C\{��
M����U,�rc"��h��q���(�3����n�IH��Z&.1ʣh/������ޓ>n��!�G����P��<՛�����9+H;�G�X���V�o6��$�s�:� {� w9��`\1z;� ,�M�o�Y�r�F��Sg�O�\A��Ϸ�V�W��w$��"W�tp�|{�8�r~Q_�&%�u��	��]=����������UW�=�:~��t�F�8R$�1� uN�Ht.^1����������rY�sN�K!�`<6I.t���W�<~�!��՜�;����5qֳ$�<�
���D��v�����EΑi�!�f�n1�|Ù=�uJ��{.c�U��a���y���x�ۂ�=�s��wm�u���י��j�.w��y8�Sp��:֝g�<�0,2y�.��g�P�m�✌�a���=M�8]A�� ��_uˊxסg�u�k!}&��
oA)�E͜��9&'-c6�-ey%?��z��H=�R�y{�3���,l��������݂��,�M~̭����_[f�M�>%3�����4���?#��g��^"z��͊��'�S�2?����'a�TJ� �Q,�i���m���.!F���y��O��LXN�B�������;�${�*	�_A�x��T*χ'�����տb||��3�1^��%�	ԭ�ڠ�ω4<*hg^%gWu�I$`��\�%�[&8�!����Fۧ��`���m�s�y$�Q�}��an�������R�Qvq;��m��w3�0�=}c�s�
	�Ȏ�(;"�k8.��o�	�vKcQ��F�0��y�K�u��/)b�^{z
�rZt
fn��HӸ �L|��K�,��e)����^����tNt�, �zޓO�*�����	�PJ����MހZ_��4l����sE>lU�<���ށk��I�S�@
}έt9��衡;?z�Ј1ޢ��M��klk�?�=���ЍP�ǯ���l�=|�2M��W	9 �x��qV��`��{�r|W�w)da��Wa��k����B� ����V��2I���x4J���u��o'4ẗ;�^�>���<�"�6�K�/��,�|%�O�?�q�)_7U�n`���|嬨6k~�g
'���N�c������6��\�\H_֑��QG�Gg���:L�-�s�YN��fؽ?���-���R�Q��iU��e!Ѧ� u�jD�!.� C����6���`G4�XΜ�ڼ�g��X5ؗ�s���Y�ʨ������ނ��Jt�f\�>L�B��E;��J�:���.�3�~�?���bD�w
�`ߦ���l�2k�r�`ga;�Lh���ndq����[%��ȅ�ݲ�1������8��uZ!}K�:��T�w`���nb�RϜ�j���]D�4�UG)�@�F�&9�/���E!�F9�� ��Hd��F �H�g�&��.{���s��ňb5�LD,��L��-�#3���#s����+��͞��L`���ed�է�I���x�Á�i��Z��P���r 2Z�pׄu'���I�m]_��~	��:�v���N�m����^��đ����5{^�n����0���J��dX�o.�u�L_���1:s?^ /W���c���H&KV�Z�B�N�+_��F���Bxq��tGi�v~F�"I�LKf�u�l��^Y��m���m�=��Ft��q.:�?y��ԛ?���B^jj��E-�u�)��<����ɍA�c 4�q����n^�{T$w�����d�d�����x�п-=6��r�k��RM�󒹴�GeZY)�3�"�/�lf򴥲�E�]����A�;Ș��0�֬e�Xt�Up8qe���wP,Jo��D)�A|$�lk3_��!���tƂ��i�&/_���7������Á�\H�Utf>�T��t�w���9k���.?k��Y(z �K�y'�#��b�G����d4&�L���
(V���C��9��n�'�+h��nS�{�C7��1^�airz�
���>�pH��ߥ�w���49=(��; �s�G�B0?�$����r���?+)�z�,�f����r�].�$� W&���)�n��Jn�h ��Տ��-�Gb��	�ԝnc�>DŖ�Cݵ�"�Y��E!�>�wP(9� ���[$�|���e�Ȭu�^�\�P�u���Z���/Ú���ϝ�wf1c��޴�-���Wq�?@o+T{��̓�G��װ3��4�O�7�P*7gm�EbZ	��*'������`ʴ�~��p�l��d�aZ��Y~�m�-�����//�p #� �Rʌ�V�0D;�|)��/J�V�R0�������#��l�~d*uq&��o��x�z>��� �v���Q��L�M����E�RlkQ,���B]ܙ�yF|�)VMzix(�O�qn���o�kv�K��2��w�����E��I*H���H����8�IK��&(�H�KBY,�/_*�j���3DI�A Bp�2��z �|�Q�p�-��r��ƺ/٫�)�B�ulC��xu
z\
K�A�h���5�:�Ҏ�&s�ag��͋UC�ȯ��b�&ȃ�w�}���	�I�/��a��5
M[m_�am���Q���t2Yǳ����A�[T���J���:Q�|�8Gs �sLõj���C������y_�D�ۺz�V�K���ji��9�B�.����r�剹��M�Q* f�����q�Zm��AN��O�91�[���N�;uDQ�	�#|��3�GZ�� �oX��4B���iCbZ'(޻H��w\m�R�4"^U�ZRC&�P�|�'�Р��[��|Ȍ3����oEJ��¶�us�|�sy�w�Q��
>���nArz��d�&�Ɯf1h=��*��=�=/�ONj~QR��J�	�(�TT�'}Q�a��W�<Y�D�O��G�iOw���T��n8Z����D��ۨ�+'�,�5���
<����9?�^r0�y������T�▂�X�V5(���Ƿ�z��l1�Z�fGPҰ����:a��9���q?��?���i'�\�p&*�*^H��!�Ǒ���<�W�uU�M�Rz���g����HZ۔���7�Υ7W(괻���� ]����NIh���l5.���߸��
��7=,p3��쬺��4ä�3�4��o�%d�D��Q`���Ǆ]��>�5����l4�3���Zd-��il����mW8J���5MU���B��s�8o=�ՃC8h�ʸ�F$�%w~�\9x/���x�cɓ�!��t�<�j��X�@1�d����3���m��;1��	��Ht\<�B���me���fms�39��P��*�Ob\5�6uf`pb�d�\�v=�1kY�{������6R�110�?�v�\'�,�D��V��x�*BK�P����F.(���ã��+�ʎ₤��j��3@g��Pۉ� �?O�#�$�
�oڋt� �͜ˮ�؏�s�vҴ�n_š�����{Է�<�2%#2��*&?-
Eݍ�xԨ4S&i���pIw����[����ky4�ZAHJ������ۼ���4�/ۧ��Z�w]���|h,�mK���br!Z/53u
ʌ��{��mct�����;f*O�֦AW��L@�)Z�
Q��� >?�t���'-2O9��ϮF��x#�dfG�_a]��p�;�l"�r���U	+u���|��QȲ�27ht@E��%oT	��\�	H���	�!#Y�/��e� ���շ����mTأ��D�(;|캖$�����}m���T�^���'�L�I�KP�R<�U]7�8��"�3|������5�"(H�ԓҫbyZ�'�O�.$��[���9N�"�,^y�H�lh3���F4��hœ��\��zdB|O-��.5(<�LB�(�c�����	���L=ţS`LY8��y����u�6[E��D��'J��t�gW��͈��[���7��΍�?$r��Ej�D%��˸�FQ/�R�,�G�1/n���sH�� ���ӏƥN���e��!*�dly.g�EH�� ?���%q�sK��C�x׃��pQ�M��f2�:���Q�\~+��<���s ����ʎM���.k,Y�D呼�Q�C{�ϟ�<j��Ih���)
D&�شQ|���z���ID� ��s��Bn}��1o��`����5y[�|4������*�Jd'
s��b5l���C֡�Ċ/
#"�����`P�>+G��z�z��=&<qYV�@'c��06TR͌�|���\���2F+^�����9�c뀵-' ��U�؎(|&�ț��z���=U)M�"�ga�b~�������z>g q9���Xo ��bv$�15������m�8�v��X=PR8��̤w����G#�^����,�hM	�О*�����,]&*3
T�f}�:��ĬzO����4%�&@�Rq"?)��X�R�ˣq]b3����MB�琾�YMs�6�	̓���aPכ���V1��0��ު��?zk�S����N/>���[̤���� �6����Ԛ�5+��\a��G�ؓ�:E��f� �ҷշ�Eĭ�%0r��8ˤ�F���WD֖�[Kx�. � ;8Ӌ1j��2)�&�J@v�p2 ��G?:Ӓ�j�
�G��yX�6c��패{yM��T����2�����p�+�����{'bh&��1��%7�;��ez���$�46�=�<ƨ��l�jWek}z�!�ce���&7MK�ʽ��B� [	��{8����i�#��Z?����0���,�Q/�é&m\V|D��̻=�	����l� we�a��p�U��d�T�G�/7��J1����[��!��E�[��Oc$+��!J�MO��&�3m��][X(�^�]7S�dB����������+��ø5H�*�F�������H���jU���ƈZ;�J�dͶ���z�&�4�����ӧ�;u=�z�N���~.�ǌ�?	����νt��aRRf���t���5æ��&¿]?�=n�u_dY\�����1��"���ǁ5������O�`x�A~��s������)�7�4}_�
x:��=��T��Uu[ڇ&V
����+�Y������n[�C<�k��5�a�J|�1�n{*��\t͗��t�F�]恕+a��J�B�+�u-�$��c�]��raK$�	��j�u�3���g�����՝%��9�;O3���	̮�B��T-o2��i_Η�X�b�I�/؏@����';��"G	�~�j��D�ׯ�j�6�l��]�u�
��쩧RL9¨��3��I���/��z�J?!߁�LQ�؆譝�6��;��V;���X���%�����f<�!�6?��E��['��Jt�}.����ݗ��O����"Av*t3�U���@s�B�=GnH��8)�:c��E$�%�.|��_ij8�ED9��Ú0���ߕ����r�F�E�%��8�n	�����q��"�l>H}�J⺵�[4���@��m�v+�[��i{�_��b�kDR�<������c�:���\�jB͍S�:r3��Z ��پg��-���T��Ԭ�D��d�U����z����Վ�ʚ����!*)�9B,L��oq (��� J�ڲ˝5������rg�MZ+����q�u��7�\_�B9��fN� �e�_r��n"��Su,��A��ɍ��U��:Sh"ǡ������C,�U3��D�#���:NՓ�)��`D��4��)��O>��I���,���T.H� �5���Λ�Qn�~�:ۦ��A�|�se�t("���J��-�Π��PDV�a�ѐU#>��?i�?.�P���P֘m�X���G	�#�Lh����o6	��S[�oc0Q4�e�N"d����g�.[�J����9�V����?:�HgxX��qhj�`���L�	ʍ���N$ӐlQ�Q�o�=K��|�sp�ӽ�	��a�r큂X��x���P�v{�A��<QF�=۳K2���Ry
)���D�7jWY��W��uɅ������
���5c:oe'�����꿤PZ5�e�[��۔�J,�v0^oQ���㴠����"����$mp[�-u���]����5��%gu�C�~�Q(�%�P{�{�@�p�c%�}��9�Y��z1�3;�o�Y�?���P�m�J��VmH�N?j�ة�,㨼c������}�I��"��dl,�I�O���omE��tWi�CmL'N� ���N�'���b������(�`}�'3�~�Jčux��� �R)l��9�v�c����+�I�9x?�ǚz��üߋ5Ow'ٗT�,6�|:�41�[�u>�wh��4=?@���m
*���Q��2����o׀�������;0gk��V�z mVE�E��׵z�����ܡ-����t���̂a��~�vT%u�CYp��y���U�ά&��#�>"� �#��'b������\R����fE×���V�A�kAJ�;.��L����Pj���(iOe6��Z�5�K��4�t�z��h!�[�:-T�
o��y*���
U,�Gõ��-z �c8�'7��MFj	�r���Km���*��G9��Ȋ�� �_���{V�]�ā�9�}�����=�Y;��^�����8���,-��=�IP���R�1��� ��z=#A�,#I(�'%O��.59�d1\�3�H��Flɰn3����V�����U�_L�%��"5*�9���+�3a�S������Έl\�,V5���@�:�i.��P$�E����YW(�����Ck��i��?6�c�Q��� Q�\g �������Q�z�M˺�H�M&�f���U��a�k���B��9]��_�T2�4���R_��o�w* K�3�|�iQm�WfE��W���O�i�Y�rzn��!/'�	4������s���RT�����z8��k��x���ZD~����C�֗ �5l�g�i��EHdJ����p�Z�4Zsz��t�JU�z��+���&�b�~�;x\�����	{���L��5ۂ��pl��H��F�h�by?�i������-uTνY��b��9��;��s�D���
�֛��ȁ��B�d�ȁ,����ɑ9��m����*~�N���lrd'嬌8���֤�8��sA�;�D�H��oA��@����c��w���D�K���YC���o�~I[�ڍ<Uެ�Vnլ�^3� ��R�ݡ�(	E��E��RR�ϙ�S�;��p3��~����
����zm7�C���j?`U2�u;c��&��[6�Yc�02gc��as��+�Eh<3h��b��`C��-�w����e��P�0�}v�j��$�I��Y�X��p~e/�إ8ǅleuc������U���]4f��,V�胿�W�G����b��l�kM�ԥ�_�wz8.��$��ޣ�\(y�j-Dc�p�ϡ{Ӊ�<��I�]�ܾ�A����}*����FuL�"/�D��|#���ǣ�DY��c�N�y�uU��:�r^R�fhL�3ۙUn|��[�e�p��Z���L�Wʖ����4��R���$�Du@�R�8Z��]4�2)�aw�3V�!��
u��-I�况g]>���ә�m�p��o�3�ӌ1�΅_Hq^E��f#�i ��^���q��rvk�ǆ:/��[�����=淲?.�Cr�*ߏz�C^*���P��u ӥ3�2����8�WKX�w��ҕ8��uҍ@�m���j|ۮ���$� ��Ż�H�moԂX�ҍQ�G�8�w(�E~��o3�}v���`�fy����7n��=M���*�xH���d�M��O��-��0���|vǘ���:���0sE��O�t�M����5�g��\\:��M<|�?�QI# Z|�o����߱ �8	�J�����A�>��3�CfNV�t,z�:�$ )P�3[��J,��^��{���G4;��7m2�JK��U*m
X\� �
���v�=���D�h��_����|V-*�[h�نE��v�3��8ӹn{��0)?�^a���;{�Z���,T@��G��_6zj����|�-�u/�v��}H��Lbdsb��L�X9y��~��_q/-P/�m�&�d�mk+Z�H]�5���OL�Yi�����X�כ�t�Uc�)�%�*0?B��&k����mE��֝�n��J6���o������Osc)+zo^Z���?vC�!c��V��O�����j��+��|�fc��?d��L���&Wp8��P٨E���/@}S��z�K�����<G�&��A�,�jL�^�,��&:d��$Õ�z��p���\�#�T,Jw�kxT�e�w��&��_��-*�p0}HzU8\Mx�ױ��ZĹ��x�!�H<P���9е3�#~���X�̄z�< L��疈����A	b��#���c�����t,\��(�����}p�f\�B��_/H%
�3CS��B沥X�/���i�S2�����l�b6�Ig������Е�'�9)}mh�(�`��FY�T�.�f��� ���CM-�\��%�Q ��3)�N�g�;��t����}	��h�x�:_7Pe�ޟ׬��2T��6�m�z��]o�ي��K���#V��!��~q�A�[����ᝫС=M�Q��݊�Y�{�O��n��S�����g	�1/:S����Q�
�h޶I����DW(Th���1/��6F�G#�/��O��9����c`�#l���(0�ͯ6��{ӷ���F��Y~��^��òj�xԚ��
Aav��oկ�D�^#B����q�@�If�'p�RGܙ��1���X�,$�(��d�r�E�!�q%����^s��Nv����/�Ś}�m�>�/b����\|�TPC��[��M�D�@֥-�T�������a�sԲ�XE��p�У9��	��(
��ո�D�	(�����۬+%��ş�نv�L�� ��M�V\��0���=P@�c�E�kǻ��W�"y%�S�P�*u'�/���V p�g�=�����u�~gF�gmW�nf����oY3�*Bd��j�5r��&Jɺ�b�	0��JP��d<h2c]�~���$z �-��I�1<Ħ(*�Pe�L��HBRf��L?����cb}�9����ې;��L�@�'�x1��4n#�n�Z�'���ز���uրr��"Ð Û���3�)�_����m�ä�#lW#l�L�f6�u�;��*��`{�l�V����QDZ�6@��.�o3��t�<�j/�v-��qŵ��I���9�ix��F�P7�q��ϴ`yn�8�o��ʔp����G�)/�!�Y��y�&7����p4�M�X��d��[o���㾙R~WO:��qA��$�%�v���L��W�#������s)�����TI�'w��1���r�1t|���w�E��-,D��k�V�;�Mgi�����`F��VMs��%�,�[$�>�l�(e|�.0t��;�9P�,���>�wǙ:?�Irs�}�|����f�妓B?l�D�Oʧ������#$���]�V�D��/;���T��LS��Y���#FiL�2�e跂6�H^e��l$��{��/t����nYM��͖���W�,�H�+�Ii�g/�<JM9[5�\I�
@U�%��O��:�:d@~[�&����8j�*<�R�h��=440NY{$g ���v!zuEt��+�o���_�u�=�y5p��(o��� X��Y�"�%����xo��4���{м`����rn6G@ҕ�S���*�?Q�?;�i���N����Q^�L���޵k�݆����`B�9�M�'�q�äRwu^>�.�d��I~Ɗ�ra�i� w�ۻꕬ�򘨨�'g�OM)�������O�<��fj�q�+)���/��7�O�@guL��~[�ר�EN�+�ʼ��bu����1b>�����1�L�I4`�^đ>�>����-R1_�%�Π���^�[ի������>��������n��� ��S�n�"����Nkǥ�],2C�e��n��<�?�o*I��z�������J�a\�t�y���X��Q���Rv�E�aV�P�;����7Rq�Du�:��g�
A����)o�k��+��Q�y�ƥךYa=�1�buJ��� cb�Ӝ_�i�63�y���D��x~4�����ۂ<�*ǿ8	�.kY�	~ޛ�@&&F07 Ƀ%�]�k�!�M�8�b.ꅆ���hB�"N�9!�.՜�`V�.�R)�.0#��79���ʿ:��	���}�+��c�ƶt�;k0Pg6�p���Q �ph�yh�<!d[%o�����Y砹�?���P%&�g�H�_�y?ĮYp�ѸRm!���g�����F��jd��"WU�c.�����)����\_~��r�Ro4���6�S[���:�֭�����������t-��h��aAC>F�^����'���
bJP�pSM[Ӊ�E�ZJ��������I�N�	�A1qȔ�8
�v_$禋h<8�ȴ���v���5*5�(��0�+o��}o�(?]<y�Y޸a�)-�	4�$�p�a
�Iq	R1ֳ����P�J�p!�1�W4U�`��)���Q�~��.�dI��ޡj�[�{-�aJsW�����'Cw�FP0u≋@����D��0;�k���^�����R���3g;�rO/����?6\�|�9����BY]��_;!$����7�t}�x��;�Sx���0�����Or����/����8�#��i�����GU��4�U�/��d�-����m�Ҩ�7@�����% ��p_X\�ZlI�>�_O�i�3G�i(a�'����Lx�M,��H̱��-Ї�ۏ}��d] YL��IPT�� �kG&T�d���b��Cm{v��[�~�UD�?��H�6� ;�'?7aS���[�n���iQ��~�n,쒖��S����=$S���ND AQ�J,����<˒��"y*��Vp3�S�V<'���:��W`��Een���<S�,�0��Uu`=Nw럟�h%�e.�9��VHM�nM�n�*���}���ݻ�ȘU��tkvTr
ez����om���)E�.4�gv��l��(a)$q�Q�w��>�����\1t0���w��~	~B²���M�nߏ�i>>�+���w��Gy�����nk�E���K+���/5�^�G�}���j�t�#9��񝌎D`���lG���k����QJ8iC��ҿ�	��W>|^��ܿ�8;o'aA5�h�#�M���&���x��W�b@��� 0��uY6�"��h�����z�W���(�2u�!N6�fQD/��5qL��.�xoy�C�O��Q���aB�<����V@�
��@+L�f�R��RE�/`���OӄJ؍<������5y�J_h�U��9��3�u�%a��$7��z9���IZ�a��#+�n�][`��ۤt%���=&Dj���^��i�����c��^C���a ��2�~����%�:梕<��W-�w�C"����N��Pb��`������Ԇrd�t�{�`���si!����[.)�P*׈�Gȳ3	@G8�n<�Т����#�b ���Xk���z3+)!ć\X��3c��W����]�	������u�k�Y���b�v����/�"	
˳ ��<�-J����fE�UK�:�Ʌ��p�\�w�ϬԐ�_�R]fP"�F�|"��q�:\��>�� �a�$��EǢ��/*�I��=�K�]�!ǹ?*�(���n����������r="m�-T��!�IE�jB�Nᆤ��S3=n�d�٢���*���	�^�Ը�WrO�(M*ܝw��-�ܮ;���jy��p��Wh��eB���$����S�H���}ߵV��p�[_���!|�(r��Ϛ��N�#��?�Ae�഍Z���v��@''�#�:Gdm�XV(����������z����������g�R	I����(}������L�<�J�����x�Ť8��:�y����i��s�M\��\�i�R�o�T���d�35z�.@
b�<��+�Ցwe�}Z�*���-���a�	�l��y�Y͟�[:��u�ゑ§|���Jz��s,�	��Rg�eS���q�!��Fu��ʹ7�]��3ǝ����:�-C�u V��R{�vә�����taTj7��V��	ka�/���26*ǌ������%��7��.SZG���@���]�Ύ�/!�4�cc�%׽n_yn(�v�rpg�;��PVk�9�3S��j��7�yd��S8�NQmюE��'��y���H��s����v�/���X����b�v{��-|SSK��jR��B��G~	(�T���sR"�&���/H�=�^ӄkhـM5Cމ�3���Na44/��A�9<[ʐN"��� X0A��/�0���6��z=x!]���5�(
S%6����r^��]v�z��Ъұ������Ҥs=���>me�U�Nh�J�"�������?5`J~�$@}Z�C��T�����q_��C�����Zń�"��:���݋�/�io�J!o��d��8|�H\�B���e/�u�$�D܏��o���?=N��=��F"๟�#R�Ẅ�m�9[�tj/y/w�'�ISϘ�����\iػ�Ur�D�}D����R `p�0�L5���b�ѷ%{<|@IfJ��1s �-�qk��P��d���2d�ɭ2.�Gf��5-���S�o6r`���K���ݩ�׬|���,Ƚ*���e*g�X=k�ҞM��Q郄q�ܤ��P3j���R��8�0�f�z��q�M�mo��J����'û͢H�*�Y�i�J`��w�����Wmޜ%k�Y�� �zj�`�m����et� W�NP�-�z�������/����9��7yC$!�$T��c|y��n��N�*1Lb��a��^��w1l��6�������	�u�ѫ,)۪z6�٧�5΢�o�T�KD4�U���{ż�կ�yS��Y��X�f�#�Y6���Ӕ���1*j-o�;�^��L.�!|�[x{����Z�H��'�E/�\��������ՃF�7\7l&H"���O�:1E�wj�8�|X#W5u:|)Y�c�@�ɩ�GK��R��N!��"&�)��sR+�5}j�reY,�;nc.���K�NQ������ׂ"�/z���֟z�$ZSc��q�Cq�~�筭��7�B�D.m���#7��Ϥ����y}������P�&���3��cK��յ���2��aTN�Sk]����6���xV��DQj�uC���X��z?��;u?�q��ʆ�z�+`���*iљ�e�#>S�5��`�������*|j��r�W� f��o@M�������t$0�*0�#n �A`e�	��,�5���ϠX�j��Ftի�?��`�	D ��t��凯&�4"i�v;��Rr�L�N��q������������
%����Ҧ�xT-�Ⱥ�z�C�e�hv1@��Ɔ/}K�L�Ng��c����a��o�+���s�Ԥ��y/^C�g�����+}ò=ϣ����b%:�������iͮ��9{��隞]����#I{�Sq�g�(E��/�M�)��2#۵�C�0�����1q�[�{��5_��̶�I��Uo� G���є���Ub8��c���I���T�1��0v�o8�i+��x��H���"@�n���b�}VT6�������A#���/'(x6ɡ5b!
�Y	&�s
9YnԽ%�C�w��� �ҙ�6Nս�*Ajp�r�m�!��h]��Y?��2�����q���[d����[�C�"�>���ܰ&(���������b �ޓ:S�0�n����%�.K���)��&AE4�s��x<�+����>�'G����r��Y�~��|4^+9^ȴ:��`@��^��(��?N�X#���p	��qTbj���m,h�� ����HB34B���Y���b�`�IJۼo�F�ם��b353�:%�\�1�ܰd��d�� �J��k��A��HRZ��RH���D�S@ϺQ����5������vVl^�Ee��g�k�ܟ��ӏ�CW���Fm��~�������wW�Mv