��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�o��ȃ|s�Pq��Ty��AG/�M5�ɑm�.]4��2��(�i�a�P%����%!n}I>ǯB��QM��k�v��G&rA������C`�����Lt�<�-e�X�T��t��*����!!��ڥ�<2�OjK��0Tp{���!S��"��>��h�{�Y+X+#��.>]���o���zH3�~Ǜ��,6`?eJ��A�(J���gAs/����;��C����Q���f�#��:�{Σl��P���I���FG���5�����mSH�M���y��܏���5@�օ y��~ViD{��^L22��b^�k����vb��#�ͺE����>��<��d�5
�*�W�1^�������q?g!N� ,z�7��7]Js����9|f�3���5u���Pd��{ܾ�p+gT�5���s��!�Q�['�������&�-Q����?g�#�e7;�1p�i�V7�c���m�.��'��A�f��r�bB_�����~�������䅀hs�w���o/ƞ:�|dQ �q��q���r)OTﲫ�Qp�^��Zh��8�����=ZJ�R&=u){���-f�F��M��7��_�4�z���N��/��$��������;���S�m��B����5:�.2�G�2i��0}b���� �ʮ3����OS������\�|�mǚ���K�*-�}^���H ���dP������WH�67�GtvZޗ�p�H�e�/Fȴ"���p�e��+��؍'`��!������}��/�"���C�� TP)�d���
�92�roV81:������޻:+����(��;�D��ݬZ�:3����V^q��S�Gj(���w��ӭ�z��MU�K�o�L%iR�	�m�>c̿���]o�H�����?E��Ff_��㪹}MÚ�E�	<s�k���sՂVX��\T�?�	�ϳ��-�����7�A�1�ḗf"W�L�:ulu��;$g�4�[s'�]�d���9� �\g���'�|�D��s�^�/f������,��I�(7���f��m�����dPl��Q�1���xɭ�VM�#zow{2���^5K!�hJjC������ږj�E��� &���� ��zR�z�C�!��-��K>��0cM�K-���S��bmv���[ݢ5�7~�@9�,�O^����F�7C7��^�$e\*Y�ɪR�j �3��lV���H5i�>�C��bC������4�")aνE4ǭ`Wz����-�1��4+q)�O�c←BRW��>�r����H&n��w�-(%ʜZ�����R�L|/�&�rě��|KT�`I��?٧��X�^2�е4���4ѣ$B�bT0D���u<�ɜI���.ϨIvo9y���Ӻ�q-��!����J�*��!�+�D��@rN�lt-��#F�8���!�;�B�t�;���{mh2.VE#x?VP�BF�x>X֘��ZcF��g��bV�<H/����v8EO]^�"�nI���52��$ٯ~e1���A��n� �I|��I��Ե�G���92LZ�4��c��c���l��\B��
�Ӽ�Z~���Wv�gB_�C��KȎ"D���{O`Xab��*Zp⏃�����,�$b`6��Z�G���c��'��8Q��z�����ݯB��w��&���Hp����3��n!�X'F�7��Q;u�"�7h�b�ň%]��œB�N�E��6է��.��mk�LPl��غ���Ǔg���j֤90������n���v\�Ta��<(% �4d�nD����휢ȼR�´Ɇ�h
��*�um(Y��Ȟ�Nֹ�� ��׉�q?/��[�B����F�ʎ�����n�d�mP��e�׃孿��f?�����]��,'����;T���z8(V%��)ޡ�Y]��'����YgG�LCI�E��-t>�,ů��pK��A�^I�9�5��Y�
't(�!�W�X�n\��b��yA�%h���ԙ�y�H�~c�� ���HP�Iʙj"�FY>�5�A���51f��k�Sq����Y"�=��'1�қ*`�61���=���'���ʰ#-���tz� �	�9.�i��L�������1�.��m�Ѐ_�|y9U����@��E��_z�_zN�����_D߽+�����#�c�/�P��`{�C��<C�� 4%.�S<�ݒ�뽁^䓓�[����W=�}]���G�*Mn��Y�ų�������qb�7�Mr5 ��ޙn���j>M:۹NĎ�`��>�:Lkc�i�^]6+� ~.���9�J��O���wt��u^�Q�|�i�4y5l��p��Vڣ?$[ϡ[=�Y텉�R�˺g�m��9}|.p@{ʆ�*[�X
�^�p8��$\`��GB?�UX��p�~�������K���
�G_4R�:q��>F%?�$�I�����PV����n��@d�A���pC5Yǯz�j�S�<��^�$3����v"�2�v0����j[X��Mx|�xC�9PcR}R�:�F��5�G�D���pxW
1f&
`g�z9�w�Iq�j¹~ �՗M��.N{N���0����S���i.�vn����r�M�Ôa���hB�_�G_n�`F�IC����*{�/ ��;"��^X����_Nj���B�X���&��A�V�Xj�2���4�r���g1Tx��H�+�b��ei���C��+���iK��c��Ѡ{J�vl��^y�U��~ͯ9,�Lf�sS��qݲ���np�L�������n���8�~��NKF�7�E��";����YV�dW�:*����=����C�$����B���EV�ZE$,j�1���'��M�i�R0���#�33˃���7����=P=C�^R���)�g�����!!2w�γf5�L8ӄ�N?�P\�%ۢ,v�P%�O�.���XeSdˑ���ބ�j������pW0V|�L;U������%��B�<jk��wi�o49��}� �G��7:%T�u��6�o�6&��l��)]?5Yr<�P�;Q��[�e�s�xM�-�	̉V�Q�&\�V �Go��a�0P�gC���.�_%T��Щ(���$���-�7�Q��B�&rɡ�1-�(�E�')k�f��p�Ѳ��P��������o��ҏRb6�O���Lw���'��P��u�W��tZ��.iC+*���]�F�����H��L�&>Ӓ���N���ck���/�&[����e���k���"�ؐVZ�C�`��@|�����"T��r`&S�KDЂ@��K�y8'���-8��9�w�o]����k/���,�yؔ:8#1E5p�yO�7|9Y0�q�!�>tL#P�D��I�}h}��#"������t��6�ܠᳰnw�j�� �+S�pj{9���bS�˘�no��	��4�T¹�-2ވ�X�YGyI>!=K�C�Awf)tJ�XW؁Kk�����2�hu�
����O�4�
	ȯ�Ze\������Ϗ�}�S��ŉT��?�\$��ս�}�F��lG Z��_��g�x)�P��I�.\K���}���If�GrOj�����fܐ�n4��e%^hn~�9�*��2�I9��Ѹy�����^my5�ʅ�]�B}2m�um&�v���ejE����3?'\��Pk0(eu��e`\���������r�\�Ig����y.WN�bpb�/�zq|[�F�������d �M��&��X�ݕ���~�,�
�M>�1Y)�дG��wVB�y0oV�j\�Ι\|0�hu��P냤�f8�9ι���P{h�s��^q�t�J�H2�	N"����,U��5�Т̗ ��q�z
}'��a%�$�9�A($6����Nbq�P �\#D��hfA�������~��+�Y��e��"���W��-,۰D4�~����]k���`���礇7G�{��5��ҁ�%p6��h� 5��^�f���9�߆h�U��a�[3aj���dl���qАE++2��E��<��v#}�/���"����i:�g0M��/��ਯt����4�v9R�Y���6����1��)��c���W��/�E���������b�g6M�⦣��ܷ'�e[�̬����ҷy�(:��g�mܛI69�bRP���f#��͓6�
N0E�e��z����¡�S�:{����h�x۱Q:�gT�hN�gZg�zw�E�*���S\�������1xK��n��V]�n���(���eG���z��	��]����Dmg�X!=.@ bX�3�_��_ĳ�ф�E��s|/�߬P�nLi߾�d�W�����߷{T��������f����f��[��UCx�5j2]M�|���y���K�v�v�� ���Z7a�F�5e���Ca�NJÃ�Y��q������M��4f�P)Xp���<�5d�J�3�N�t3v,a��p�\m�>/��/U]���ݟ�nh��k�ug��m����Ē��ʰi|�^ ����5�杓��)����(���'���)}d~��a��b
��2����T@�%5��5�8O>��: y��~C���g�*Ռ.���W�Rav��Fa�ŉ�������$�?�k2�)�A�Z�@p"ɰ�E6�2#K��Wp�H�z↰\�_x����Xà
F�Z�iOZ�&TY�9mQ�v�f��f����:+���e��<C�%�z�g�����d���h���{>�En#D�?��f��J�b�|K=�q�hG3ٮ��+���8�x�P��[���`�����H|x>J�
+r�%������D��v�1�lw���F��7^����b}�N�ɦk���۴����K���!���zc)FY�Q\�5���E�x$p��͓���#�u�ls����
���`N��hJ��0�i�`G�(�Gr~����o�a��$z�<D>k�g��*���@�(�ހV��F=��|K>�=�%�s�kƞS7�wU�q�S�����i/]��0:���V�(z�iU�g@�c��(�z�?�s:�DtsIX�$�GP���%�C��?�VL����&��B��gx"���&)�:��o��gU��� #���>z�\�K��NA���ڪ	x��u���+,ܑ���(>YM?"Q�N������Wa�\���tC�NS�/u��n�~|e,;�)���iW�]DIB��v<IԦP�%��q�^5Y�}j�-�;K�LU���|��K������)q��%����b^\���������H2&M�B�䌰�Zg�k<���Q�J��� �{R`sN�׳�I���C�t�6&u*�Z�B�C�V��8w��tsCJg�Ns�ʥ'%������L͚���C4@�eqށ�iCN%�ֲy���e�D�K���ԾSa�b��#��2����֗-)�&��4	=s���k#F>s�o�2uI�{��0yz���I��g9M�������Jv�3�_��?R�j��<�y���9�?79p���� v�}uɞ~!z�.4�����0J='�D�kx��y/��\��3������/�#2�0�e-��d�%rW5l��]�T�!����e�=i�aE<�cK�|�A[�����qH}��m���zr+I u����?��f*r���0��zޅ���tZBAi�� �e���G��u��y��U��� ��<��j�6�?J��yC����j@�Q�n\����m�2�*�F<F����m!q�`Шw�[����k��5JaJ�|�����Vd@	���k�'���g��bmf.�X��1�*��D�2O|n�\����cFÈi�H+^:�#d�F�%]p�"Y�,&\�������
,ذL����j�c1dK�l��@�`��߬�F���40�,4I�h�н��
���L>�I�5�ݫt�����%5����/�E�4��|��H��;���	��O�F�<S�P��:��}ם��;p�NƐ,�<�8�5QDv���$sgk(,y����X�ٞ*9��?W����0�����_i�eo�e��Z
��Ò�*�����.�b� �B�o]�C,\��f|w~�)���ɸ'Ą,��[�c޴��W)*r��8Ě�l�ە2��ͪ%���89@#֠Zl��0���)�:�O.h����Zet�Y��*�f��w�4�1��Oԕ��KJ����Iے �Mؽ�zL�ݎ�r�I�S�ؚ>�P T׷�9_�#�r��MhOP@o�����r���v�r�x�+�LU��J���c�4��t�4=&�v�1���9 �ƕ�������ŉe�+�Z��m�����R�:uQ^�`��88��"yI�d��ㅴ΅�F��{��oK�k.�����ݯ�7J�mƮ�e_$��j�� ��寘?܈��7�5<�g}�l�H�ưN��X�����[��k�R�2�Ҳ(r���,f���+�x��	�ԭ?�{ӊ�4����:ׁ!����Ȕ:G&_M�u<(�n�ya�G�^������R���I���r0N}�%+:i�H��W��Eu���q-�3�x�F�x
(�LL�:�Z� �D�T�����q�eǛ�
���@�������pJ\�5z|t����g��=� �P]���� �xE�ˣP0�8xҟ�����5�l�9>���"���l5�ߌⰣJ�ʂDCт�p�L���s+�����si��������'	|�gb��^��(��9D����0i)^���%��{�I���L�Z�We������F��d���k��
"��dH�̧\Տ������c����Z�s��|��{�#�%b�v�x\\����M������0à�sS��
`�/
ڈ� Av���/5����->�Vu[���z{����X�.m������ �#�1۾�կ��.��L���D��lY�ģl�YV�h���*׈���3J��6�b���r��ʀ����
��� ��V,0�������t�Ѭ�v�v��>1@$&�j���񥛽q��������]ջ�86#��-4!��L���AS��c;w�+���kG����*�AXG.��P2�!�:��=ȁv�&?���E:�"�2O��oK*���H�''l�	�7<r\_n�Yj�J�W�'P铧��SڋN��V9f/����N�g�$J�G�U�>{H{��^�rjtZ�l��f�J�[�+s��)-|,���_2���;A&Ar�x����l-x�<~N��z	�!��	�ϙc�Z�W�1XM	�/�̴]Y:����檽�&\�R��~�qI���56��(
V|���8_~ٻ*z���� ���dݞz]��h�����h)��h	abu�z����H��1��&狞���7�~Sb]G���(��L��'r� G�@`G|
T_��x��ct��68��x@�o��'P~۬����_�y���I,y�_[l�HZ����"'�If�Y��!���� �*WNoi��o/�F�%�r������ �I",��.��;�����WB@�Ƹ)q�~<���-�4�^r8Ǐ����ӡ�/��n�.d�gB��������&��냂A-+�7:� ��xY�"�/ܭ$��@R?]�D���C�%I�즔�gO�֕e�����䒱h�R�ٶ�7��� %�н>Ê?���K"��}B�ݯ:��09�/花,\\�~q��n�\cٲ#σ�"B����s�Ŏ�!�<P�nex��Q�����fdxW�C�NlLI����f�mb �ko�`�q�- XG��kI�5`�__zWl�X�o\ug�]�kֶƱ�\4�9����!�`@t=�[:���pme{���7ɲu3�������0�������Egr��ɱ<e��_��|+P%��\�����ޟ�3�)��.����|���>2����&�̳�(�5�[��O˟)�
l�מi���tg�x��|�����y}��4�td�-����F��� X*��%�f�<re30���,���eo2��%�R��yƞ�K�z����4����K;��EPگ�ʤ��IY���C���:�$���RA�(h��R�=���ߠ���\�d�c�\�����<&)p�s��������������5�DJXC[|��`����M��}'y'��jW��Ys�I�˂�y-�Wjl���M�~�"X���Z��giKZ�[�ߺ._�o�̚��Gi��N�iUۈq��zA�K�zVK_PS]%۲)����CA��!������>�w1���ͅ�D{�f���%#Ѐ(Q�d	X#غ��+��rf�JuPN䄰����|���̞V(�$Bzn$W�L`�a�Ōl�����t<c,wK�MKjp�@���G������,�H�"ן���(xd�!�����O�а�	��\gњ콉�G�a�sO��b��a��:|YM&��@��e��� 턠Qy,b{]���(���pEۊ��Gxw��ͯ��w����:�f1�'1��?���Ҳĥ�����TΪ���-��`4gJy��c����� �|oI�[`�H�G�=�/�W����U5�^�y)+�ƹ���B5�w�^)�B6��cd�w�8�wD(�BZS�e<����\׎��+~U&�����10�_Ф9,�J���ƭGO\�����5j�}�-��rdJh������M�a�^�t9��e?z�/�($gƤ3�-�u,UmY���*�X����OG�|<��@H���Jy<�O�QZ�=�&7�6�O�L�
���G�ڲ�{嵿%ɍv������i��X]5�ʶW~��X��B���I���Й�%;,��BAdVm�B@<���ySua������]���!���N!��"vF��ڮ��E�>�8��g�>�F�s�?�ݔ�����Ef;bdު�2��tE�}�D���1����-(_�-o�=�-�I��|Γ���#�|x��\c��Qlׄ5>��h�IP���e�O�L���e��h��'HW����	���р�c�G��q�'�;��l�3��ȺZ���%�p͉rdO�����s�W�w�M�����] �9}�d���]�V��7��f �կr]!��%�U]�ddC"sp��/��7α��-9{vo�/BE�e���^���É�=J���ڽ^I-\]c6��6(.U�sN6��U��^��P�&�?�we��o~n�u]���P��le�/��^E�@�?߼���"Ps-0��UUu�����/�'+L��5���#�[b�%�æV|�y<�єݶ��`��К�*��g0i��7|13���2"\�3��>�X�XW���7b8�h�2���	�s��VM����{b�a��uC��(S!�ۇ�|H{0��4���
ܮ��/k/�3q�gIȪ�E�6?f�����ل���Z�`�a��ma���Z}dܔ�����f8�Z3�>D�#��G�s�櫄z�T��������-�^@��oG��ܧb��n�$`���d�!�Բ��!i���'B��N��&�qH��0#GR+�	��������!Fr�����+�D��\��`��^?�b1���I�ףr��<+��Вd)�?�}S�}��޽�Y��w�#S�I�@E�ݙ�I���<k�1$M��Sf������h��d:8Em߳�֏3��?,�\��Q^":�F2��9�R[%�ōc)S#0�Wk����`x����Mo�u�S�j�VL3Aȸ2���P��a[��;}�=�M��F�L9�GQ�����gYG�$=���^?E2�<5��?&��ά��#)5��ZV�>�&�F����pBRtU����ח�j��|q��q�-dϓ/�[�W~>����V�Vg	�a,���a�~�÷�n)Hv8a᧪�6����[�y�ަ��E��r-�lcb���5\|�*�_w�ʕ�����ڦ���y����,��&̨e���2��]D�\���ivd�@n09�0�-5��/��s����·M#(�u��}+���)�U�.V�=Y�W��r�|Ҿp�&e�2P)���2�b�_�	WE�a:G����"sX�y�Vu�mb�y�����ŦĎ��i���K��L�����6c�@+/�a#�:'ߥ*i�°A52�#v���,fA�̫G�1eޡ�}�J�����$f73DH�#
ތK3R��/�3-)f�̢I%�Dt)���O��1Q�P��Mף���&=j��zc��F0L}��ʉ��!F���� �7��IWqW��^
8ꃕ�6�?�)��g��a�~K��*�=�_eL����ǉUR���աXڡͩ>�(OO����'."�k%�Jz,ٶ���O�7܇70��wɛ���k���h����1�S�"��<!J��%��Lj��'֎��#� I�����x�kEz+	�|��}K���dBnA�7UF� OB���@��u t@��5�59��lw\K*p�{�	4^7����m�rac�:��@K�9 C�gXY�J�|'�?"-�vm�7 ��lmj�T�X!qE�~�t�+�G�����L�i�Fe�2�1I�{����6&�ɝ�5����Rl=c�+aviB�����Y��t s)ӇAC�z�;֚�K�����WsVP� ��Ė��H�ҲuQ�3�L(�O�T�ܨ.*ؘ�O|o�JƇ�Y����$��y�����-�%<m�ܯ�踯�䚆�ߔ��&�h'�S��T�٘�� �/m��� <�\��6�Z��<���ݪ8>�Ky�B =�g/�״x��E���5bE֮'-�%�pW$�P�'����!��	�I�+fϙV���ۛ��uGs��/ȧ�[t?����y�V�C�.�!���m���C��4p���F�z��YAn�g�R3-���l�0���ՍjS/�A;�� "�f����]"���1�h�0�p�$\�3W�t�(�����нY���rIgWݠR.s>3bPYQbNe~){<G�xX4.�H��@�Iy�N�߾UsI���Y��3ӵ`��R��+
��2���ss��aE좟��<M��:cla����ig
:�م6��%S�ߌ\�yW6;�.^����Z{��rɑ�E��n?LՄ�)Eɀsr�-��e[%X%����GA
QL#�i[6P���W��h�����d�H����|�a+�����ds0��?�F�l��ˠ^��d�l׀���T
	�eR6�3��Ёѩ��E��2�����i�4��^�kZ�C�G3��癏m���Q4�A��$f�q�F}�#��o��Y��Ug�#v��\��fw��z<�%�h.�e�����[�K��6ݭ�S�ir�Op4I���1���R_pCW�"�.,,O�R�-yV{����O�	z#L6G��n�T4~dS�6M�ѱ,�ɕ���T^ �w��G�jW/|�/��k�S}��Ƴ}C�2���r^��0�kǉ
��uՊ4��ի�G��@�ﵦ�KM�8�����'��dV�����^&� @�~�Zr��	�N&�Or���4v��KA9L^"�	q���� ���i�ֻ��]6���4�%��#; �D�N�EaR�Hix#K�@̇�Ë��*�z���0|ͷ;w�}�#m�o1��7�K��
z����^�hZ�)-�+t젵C{7%�h<��+P"ߢ�w`�6N�*b�î�=��acdK�)w�
,����TS�K?�<5���2
g���HV<��\d_�%�C����m�m-�;��uDp��,��K�]'��i����@���"�Ҡ�J��b*Q�A�討�A#9QP�sQ+Hjc�W������ֲ�A[��#��@\ �%P���W�ͣ��B�f��F�����H���:�嗸�G��O����o�Z1Rw�x�ă��<��L;$[$lUd������&R�ձΠӞ8�&Z�2�Mr�2�,tȬ�ѩa��Ǒ�Z�����f�c��o���*�v{�x��<�x������x�&�sqN~	U�rXB��B��;�%,=td���v_5��P���I/��[q�{���v��\v�K�X���U��[CQJ�_ߠw�g�50��탒�5V�M�nLo��_aK�ˣ��I����?���L�%D�AR��j�=� �gz�=�Iq!����IAS7|���w��p��z6y状�S�Ӳ�X�����CMe�H���<���ЌU�Y��u��u�˰iZ����Н

�󊚼1�u���`�u/��_��"J1ι�y�-��]��a��B?��:e��`Q��K8>^-�	>�ŏ�QS�	� ��`0���v�S�� L�������}�9	׳��j���@�p�퓇�3~3�D|p�I���c.��]���qffx-�n2�J��<H�(H=�:l�w^I���is�]�k)���/�ܬ���;�_'�N/�Q�ĵ��pR�~Ho�y���%��<��%]itmMT�K�-[m�{�Mn��Jaj^�V�Ư�ͮ�se(��a`Zmr��?tI�/+�u�\(����L.g���TL=��r���X���_�M^L>�;��T ����g��u�S��^O�x4�)w����d�����#)�$d�Hi9�O�����*�y���d'!7{�t��T�C>_����_�X :���mFp��m�|<�Ґ$a��k&�z��b���[<�[`l�����Z�3�J��o{l�.c��Y榛��)���M��