��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ��N��������*�%�rXwl`��|�1�EQd��Lqސ���(����;�tό�"E�7��e����A��.:E�״�p���]���/�h���������ʰg������wz\o2����:N��L�^�ҵ�j�]��8�G�Y-NT�!v�.�7	8���R�TY1$���vCtIíH~F���i�é�p}4�*,u�z#wՁ��Z���x��4pYQ�22����J
�<��LY��&؎E@K�8�+�VW�?�h�(�J�]"� �0U
B���Cc��}o���{e@��U��S�
�c�G0|幖�4��K!�Y_���0�'�#��8�c�Cg�.#���NWO�|Nc_t���]��̧vrt`KX��\`��J1XmL��$F�Fy1;�t,�(�o���@���|w�me��(��FgPm&���܀��Β�����~$��.>-4���d^ ��$W�t�;4R^��Z��%27yÿ�_�r�T�<2.��������� ��~�����-{���vHG�rsTQ&�Lv\,s���[I�Ó�:?g�J���W}��G��E�M�ra�Lhd�:[�R8�f)*(��\t��躻5�j�Ρi&��:����� �{_���\����v�ͯ05�~��S_~f�L�T{[N�oΒ��� �ф9)5n3'%�δ,�H�(l?�2��]⦻$GYNwU�.��_��6��A|��h�u.q�)��a9e�)UvO�=|�ˀ3}���"�= nN�-Q|���nW��~��#S=�¬��ֿaE�����R����(�;����\!H�_�:��=Z`�������^�C��&
O;Q�����q6ԏ��e��5;�-H��:z!j�������`*=?������Q1� �4H����ȟ�=��(p����B/y��<~����/��H�`k��l���1�����f2Ga���<��
�dx�Ҥ�v�T�,��C�{�_�s�����,����BN4���'�I��d �+���gAi��Y��&�q<aQ�"�)#��E	���[�o�v�
������6��;�����> {�����H��_U��[^e��Mg���D��ҵuC����{��w�Q|�*����T ;���y_�/X�#-}�?�٣�AJ@���W�7�Ycp�ѽ���Y�Ӭ<�48���\֛��[:u���uXh�Mԙ�#�q&mF�������CE����7f����yS����Ym�V�ɘ�7ؽ��v�d�<zg��0PT�|0�G��ojt���̎z���3��Ȧ�֪_%&Q���f5�*�f'$�K��Ĩ�N����.g���"\bnk]ƾR�IT\J|������(��^�([	��ս=�Z�T�	4-�s���Y /ud��\E���lh�30#3���E.��?�j�ܭ5�pԙ9��m5���6��R��J3Ai�e����1
�	M�LЍ_��ЌW*w�iöe���̉��w]ɺ�
Ƨ���YPN���5���F�L�!���,&HzOu����x����0>_�P�$��8rgӧ��n�
����V@���<g+�X���!���(��J�=�������L�^��q�nyEsU>���Bɾq��	�"��B2�o��t+!Z@��͡_}=@s�X���᏷1��P��R��ʀm��2 �ڒ,P��z�������w|�\��*���TI.m�yĺ ���T��T���$A�u�g*�*�z���������d
m�N@)c�󧜙)��w���e����1�C憛�i��|HA���|�F~H4~���$f�'4��Q�@HA�B̏)� %fP�:3���w���Ab?��ҝ0�����۷X<Ҵ�R	A����߻t�&@������#l�+��T�V�y� 䆡|�\���e4��ؽ�����T1���\�@��o���L��h�aw���#�[�$ �����|���r*6O�~z������[\���$��:�:��y8/X��S
Ⱥ�p0)��d����8��d��LwR!<�+�`ɾ��ĳ]H��?�L�Ũq�h�ޱT\��;"�Y��nR��E��W�"�m�EYk�'o%X��OF���cV@Xi��ZP��K�Bt�+�9s4���)vTn ŏqmU�C?���扙T5X����,V�(F��`�\0��4��w	&jݘ,Bxka�M��#��؍!EX[ꅀY��o�X����<�fY0��m@�̡�:%V@62��m��B��^�6-~���oߑa�
�6�]3d�.2�	d��c%MO��#�K@
XS�Y*�������#S����x�o]S�*�A�C&wY����n����A�E�)�,�����H�E��6�B%1�9��9�)N����eoy����Shk�]��L�;gd�t��jS2���c�1���>�,^��%w��F�f#��|���[�U��J�-w%z���J��xLL�����j�����XVd������ p�c��l��+����ܳ�T���v`8�	h4AW��A��B��$+�_3��c
��rd���Y95C?4����-�oTՈG2 �~�0@����\�I�(�%�b��0��.�m�S�N�.���g�ky�x�H��:M�GM�-�U(���򶽼/2H\q���#�Y5�ѦШ���u�oK?������p���]���[��RU��VN։ˁ�7��`\�����o�^o�]��S�)��4�k�a�[}GV��4��-��s����!wAj�C��<aXf��"rqYVhԨm�v0�d����#^�q<����Ac��ʪ+��܌�~K3a�9��� �e}ႁ���n���� �q���]x[+0@1�/[��+x�4<�5�K��-ot��ʯ��/��wŨ�m�WO�Ó�� ��$���p�v��l2#�a���M��=�[�4BY�2K~RD�c��	
���f
(���vi�o����/x�����4�ձ�2J-��$���<j��g*c�����=���r+oSjS�\�1���2[�d��L%C�h�������mG�,1��y��`���7�=gh�UI:@�KVɊ\+���Y������ڌ}傕R��1�5vh5������u�.]�4�h� j�̷�����M��N�����Q��I3"nH_e���c�
QB煤S��7�ϓG�t��WvdT�k�!@�7��"�riW�� 7�^q�\���Н.M��a�F�Գ_�����@�
��W_l=~��7�j΄BX�ަ!:��O��mܱ���7m9/)m���Qa�P��*4ϧ���Z&^»��\�r?ms�4f��ZY��6\^�c�c`̷E��ǅ!F��i�j_d��������πK������z"s�lT��7���΅e7�P���,/�^�'cp��ꥠ��d��I�93��,4g1��,x߫!���\��`8 4�҇hbs}��@3+��������-#�=��u�������.��M~EW>��M-� ]?�p�%B e%y�!��]P=�V��R�3m�9��1Pt� 5h3�z�~�i�� ����TL�a}k������<�{��ڒ�����P�,_S�'	����;x��*6�(�������r7�)ͱ\�e #gGy,��SO-��q[4��fE5��"�Q�H����K���70�j����K�G[�uK��ܲ��eS���uM%�VC%��7�!�W��`�x����óc�-�ϝ1]8X
�N��Y� �IGP�x��5�i��Ā1c>� y.���:$F���Bֱ<RP� ���@��mN�5��+0|s��O�:�	1��Х/�+̙�5e~Z  �0������G�R��_D����͊E�����ޓ�#D�x�<?#�c�yϹ�cΞd�'hVPŶ۪gO���	1���-��WB��PyX2���<�P=����,n鳍[`@��ӆGc����:�4jlY�{F���S<�G���"��*���w/o֍�ӻ��n���f~i%�%+�߇�������q��@/���MX1O,�?>��s�c��M�!����y�Ybhq��ވ�e~yl�ۺ������JN�G���Y5���򠂏2RxW��+J8#|CC��"ez�%1É��S��	�L���W]���I���v��e
��o����0JU(���cA�c�`�EuR���H'�n9���ˉmd��.,z�+�8`}����h.g�L��x�O0��\�f���,��<y
z^T�#��WY����&���wΎ �Q��'^��� ��ৃe�{������&��4ȷj@�8=Y>�J��Rj�����C���FX?�R+��C��'>Y
F«%�Q���P|�����׼Ӑ�ۤꨊ��ۮ8���4�]�D�Rx CMm���[�p{��8aAF
_��'�̯� Ϸ�M��X��$��e��nޑ�锜�Yww�o�79^��]P�����D:�����lJ'gi'���-TR�*aW�%|���T�i.w(u�N�nlj�����^Yj7_`b����׆����;h|3#���X0�Zv:�Y!dݿ�05?���]�[��#�������f,UQǻP���~�2�(����u�>���ߺ�rѲ�=��8�7Օ�_�Q�>��Է�"�*0\���`�B|�Am��h \���6����fk�pt�gn�������j�r��"�� �xC�xV��$��?>r��p�Jf�f�O9��+�����J��)lܡ����$�)�/��� ����Մ�3k�ڑ��lZ�|���Z�Y&'��;��\*���Z�e�NY��{~N^ӕ7K>��7��Ũ���	��4���P3��7w\f��;�"��@X�>��|�ޢtz����R���\_d2H����J��>S���tH��]t��5q�h���7+:^��Ԛ��'j7�<��%cx�SI�ʗ��KS�ш�R[^�~6����Π�E&��n����_
�b9�3�x���$�(�.$�Eb_������jA�z����H�d&h�EVj�v�7OX�͖C�].|�YB�i*�l
8�[�%.��#E�:��cb���C4�&�U��Ւ��O�c5)	�xW���m�*[&�Yrh&�2�à��u�e��37SВ0$�?����{�D��1�K�@��].���Rkh�b�Ғ��'S<t\8Ʊ~MƢV���d��C5��2.� 7J��f��H	��oN,k��T�6Pl8������V����jf��P�<�B^�*u5�&�	�;ks~�_��U&�Z�H�K�~@�:ǭ�L�y3Rs��ݘ�1�Ȳ#7,���,՟�yIMpL�[���(�# �W�@����^��$C���w�Pz�R�zSs������M�OE�� ���n眵��ľ�Hf�OK��9�~o
�} }B��)�,xc�#9 \�����^����yX�¸�3�t����y��: Kn`gd�Y��7^6��&�Qc?���������՟�*�6xut�0�!���ޛ�~P�,zA�c��-���ǐ�ˈ%y�ڐ=���@;{H�X����/�i�3�Scj��&��c�YW�zn?������W_u�Ϸ�F!{������L-�-�iF�r��F�:��H
QJ��tb
�%���m;���e����<YT�D�߶e��\>ޕZ�Dmʷ��?���c ��g�O?���0*��=�tM����5���n}H�.�U�,�W�w$B���Y��l��g�X�E�r��nJ��M[Pـ�c���`%�"��<Sֵ�A��Ϟ]�ZPt@� ��~$�d��	�2|Sd.�P��}��]W_b�s\%wn�5�$�A��wm[���Ca�U�y�K���̅�I[���l�������mH&Ƃ����[�B!�5MMN��'!7���� k�=��X�a���塗ŧ�)��uj*4�cr���"�в�n�u�b��1<v��Qs<� �NNKϯ�^2�)�M��o�o�ȼ�o[���gf��U�B���B��z�!$����5U�k��嗗�aH��c0�5C���'!�%����B���u	��=���s� GC.]�y��F���FS����-�c��ǷۇN1�>�F�,�u��ɐ�3��	���s�|1���Ns��Oq��|�ޅ��"F:2�.��C��21��R������o>���
�d�U��5Ip��0Ψ8{~}���4������̥���D'���_m�ց���,\�8H�v���7�o��Ƶ���#TG�&r���l"�}w!n��@�^(/�@�)�7yM����{� ��De�Ǻi)j�5���#9xz�4J��������g��H�� 4oW9OJ���z��֘7����O�Nx_�����q�L.�4��En3t䌦�
�7+��.�޲I�%+�{n#��x�ͺ�t�%��5.S��Υ~�j�; ���rs>ͪ���0&hcw�D�{��p��ÅK�u�_$R�]B�n%}N����MÊ�#2�k�ϖj��#i�����\��Zk�Y.���D5W��Ohv*�7s�S�
��f��f��W,����-EL�t��c���h����h���qKo� 6�U���2�j�^��MF�i��N;a�FMٌ,�@E R\�b1��|5&��Y4��r�Zà�k�u-c牊�=�ۈ����G��E�q�-ͳ	Rn��a}�\�{�ć����&�]W���撨rL<%0ٚC55<���R���^u�Cn�w�=�H����騩�7Cx9��FpV����]`鼺�ܖ�vF��c�-P�j���lX^�q�/����X�1���eޞ+o-Wqq<���QN�*R=�h94S�jI�~]͗�ĤP!x��Qi�n#� �U�����'I��A.ÅZ�_���u�$m�0҄��? �#�����g!����`�U���o��)n#}�.�@�xg�=�8��*���gJ=�|xN�>2Y��ZԱ]4Һ��Ē!iϥi4����N MM���	hS=���kI�7`��@k�g᭽�x���`8�����y:�f'&I���-3�c�m~t�Ϡ���3��i3��ǖrrpb8;�P�h�V<���Lӈ�����;��O��p�vH�j%�skӠS�?7��&����m������\TL�uĳ'��.e�>�7���9_ =%��`��r�|St �z�Bؽ,�����9�c��'���p͚�s�W#�js�1`��
��/&��קױ2��?�{�Yw�Q�Q�W�J:�����a[�
	���Z��U:.�)�1���_�H��|��y��/#���4J�927v���,��B���SUPm�2�1#�)up6��Z��0`� �bج�8pEgX�|�<�zA�U�>u� Hn~��%Z+��nV�� �숑s#2��g�;=U�i�"/�]�a����?��E���$�	3���2CbE��X���e�#�eV���V	 Ư5Xj�����aim�<[���_�����·��-	�.&WF�0N�#y�F�%��:_��V�0ӷf7Lu�x�Z���35&k4��~������� ���Y�EX�T'��MI)�&@��&Y}l����{� ����j�;R��L����Xq�V~�CЛ��4�F�4��ؠ�>7Q����K`���