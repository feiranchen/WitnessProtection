��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P:� Z` ��DJMS���Z{��N���^�=�C�;�H�P����h�<�V�Dqe?�'#��:�.�d�~\Rnd��~i*޸�!јe�h�Gca9��YX����B���#�V�,��<P�u�j��e�5�p$3���`�1)%LsӼ��ڌ��y�3�J���f��� Bb�^�qE�7ț��'�'\vz���9^����Q�IG�^m��C~�VB%>7.�Q�ݥ�4��\���y�tU3�8b�~���`�Ý��A�sSμ�\�� h��8`g�����>g�4���}�1xI�84%?����t����]v�j���6���a)�@ߣ���Թ^�Qa��X�X-Ly?��!P��@�PM����^#�q��g�ң�,@O�Z����2_�9���s��v�E���s\�I�b/m���m��/����I���	��׾M����)����9�)̶ă������߅���"��Ad]����$t��z�	�/�(�򕥲J����uo�5]O/������ܲ������6-����#ד��t�s(il`k�3e=�$fTai����@k$�J�)��[�'�z�*���_}�r�;�W[F���q�SY+�&�^Y�-y�\��iE�;l�C�XuQ𕾯�83�����
m���4��`�?�(���
r+X�%�c� n-��BK<���t�;��:�y�^�c�0��X��Pen���P2��g%\zHz�bk!t��N��;P�P�=�=��4�j�ؾ�f����4�71���ǵ����z��W戰i�j�l���4��u4p��§�krJ�P{���3���]�-����)[��s�7:^�ҝI�abb z6"�4�>���k�K��+3�u��|�k��EI�q���������1�=R��<Ў�8��7����v���l��ڲwZ LJ h��������� ����F�6�Q�`�i@0VG1���8f�����W$��Bg��h
��ٽ�KN4n��b.*Zhfj��,����%`07���a@������՚;�N`=j�@�/w蝠E��@P�8�ɧ�G&��w�:)���o�E�d�MF�Y�X#zM��pa?:=�*�7iA`��E���>�U-W�M�<�?�㋞�8P#T� �8��j��YՑ�\��Щڟ���s"D�"J^
n�o��c��.
(����X)�Lh�Ǵ��,�Ђ5���R	#�X�$��d-4��M�jZ���Ȃ��d��1�#�ZW-F�w��nMq�HVb�F
8���`¾�gw2?րq�F>�%��5rB7x�&hp�� ����^J���/aTO��a8�����G0�ugq5�c������̃�>�ʧ�J8jjN�	\������ߛ��:f]&�<�������.�l���`�$����x=�d�����L�O����X/'����^�j�(FG`ז×	\;�OV0%Y�Ļ��~wF5����dv�C �.�V�~S�"=�}w	�� 0��HH�24���U�ׯt���)B��2�&��m�7���nHؒ�U`�^��g�� K�n��}�/�ܲ5>�x���C�KJ,1�w³^H
rY�r3�G�K8xAёA8$����e�0�t�d�O�+n;�7�lX��]��e;�YƏ�{��ٍ��#˟x{y����S߶�ˮ���X�Ű
����9���ZH�vEB*�`�A�d%�h����Qk�a>\?9L�V~a��-d�jVR�N^.Q���q�����D���5A8���I����7i-���]�ٱҜ�V�d�s6�B��0��t4��˞zw�f���:lv;c���X�WT�����-1%�n#VI�q �ʓ�
!�d��=��)ho��|���|{	mAw׼p�׵����dz)%E}���#��FBn�0����7�����#�
�{�L[2�{{ǶaX�_`k4�t�e7��V��#{��"(�����e�t�L�d2ˮ1e�¦���@6��}�"�6Zh�f���3I����վٸ�pF�Q�]
����|D��<x�J��y�H� ��l�Υ��_�H1�]9�oRw&���E���>�7H�b�7U��k�`;~��V��RC�A���kk��s�y���+:S $�L��
�p�D���!N�sU	��5D˟V1僚-����O"���[�ۅm	[���FJ?�@���.��w=��m�\�ӔoN3�RA��ܑ5�L��n��CI⿨S���֋ܝ)��	�,�Y�P�X�2{�v��-J�׈�y��A��T��ZY�O��i�a�7������O��B�]c�f� ��:�ţ~���F{�v�0h\�v�)8����,��S�K�8��]#���=����_����35�j�y�y����p��N��%��;�O�s�c�Eׅ��O��b����ߤ����ՖV9*���r	�T��ާǟj�%N��7�5�l*e��r���k�F^�b,Y��	]/,B���4�V$��5"��<sC|j� �z^�I��)|���pd�1Gk��`���	�~�AM4�����U9/R�_�jT:Đ}	5U�fX��L�3�Ô�>{�Z4��x���؞	��^Ҏ���������~YgH���,Sk��].�ԝ5	��/{*@���3�{�1�E���:�i�X��{���[�dB����ʒ6uR)�Cw��$�t��V�4�ݫ�F8�?~	������n=�e��:G!��tO���9.�I�<��Ӕ�������J��3fǚ����Ē�+#n�
��깣z�z!!�7O���i�k^�'�v�ނ�����P<`Y�Sb&�S�����Dx$��X?g|���6e��!G�O+����%�U	��Ѿ�a}/�3~�������M�,�VM�t��=#k$Py!�#���/{��6���W�����!]�w>�=sc{� �[��(މ���I.֚�Кv��wÃ���}Wb��uf��>Q���GS"�������+}v���|��o�;��׸�[>rT����8��E�*mF.��=��y��6��.�d��U����Ŀ$�.���M~|�_i�ơ��B��`$p�?SvÅ�ߡ���u��1En7NXYWZ�Z�*��n�^���[��{|�6��ou���9kc�(���^���|�:%�LȔ~3��g��v����m.)��K�9)y%���C�P�a�\�.+ol���ºg�9}͢I�C7�>~'���"Q�iC����~�����m�!�L�x�K�A������fq8�A����������;�����@�s��\����^����}$�cٮ�k­LD���q?!;�~�U��g_��>���5
��Y[��6������J�S��3��pk���&;��@:o�lj�c8��RЧz�L������I0=Y
&�+� ��u��=���Pf��'��ow�Ġ|�4?n��8����m�w�ά�^	����LS��Qr��|I�F��@:���h}]��*W�02�^��']vw�uW�RsJ�-I�Ա
I�]1|ϝ��⅔�'Ϯ��歵��d�����u\�Q$���&���7����<������F��>F����������9����}����V�E�3u �{�a6neI�x�#ϻ|�/D��ۧh�S��L"���-�l;P�������P��Ci�ѻ���-�N���M����'�e�TJ��L��X@"�ƟC�W��۔��T!Wऄ��۟��Ke+�_��7�'�E&���F;Q�t�-����`�(�~��t��!j��r7�ٔ�>���RX� �H�6'�T��G��]I��M�ǒS����m^-C�~Ԋm|d!�C����J����5~�{y�;P [I^�����\V�ntL�����3��r!?qj�� zv-�x�
*��^好^D��I�~��Z��~¡�+§W$��5�<�T�/K �ؓӮ5�T6����W)E��xAzW/ �E�{l�+f\KH����X�9k8���/���*{���gY�K�@� ���'�=yZ����o>,|/D{���!bN�)
�����.G�3H��L�N�^�����[��%U��Q�B�ڛ���vڿ�b��b�l�#�~����� ߜ�a6T��-8p�$��!��0�| H�1�A�}ߝ&%^'��G���Cc{��z_ �MYOm����	�[����
U���d}�^ m�hm�mթO�<�=߼zQ��=�I��� F�Gɚ��,[S��`�09ta�Z��G�j�׸�A���Ǉ�o�~k��.'����� ��gfFa_�Z8t�S6��`�7�%%;�N� 8�{�xG�Xp�Ъ;C�l=\����Ȉ�daw_���#���Qxd9&5x�bp�@�qKu��=��I�:�)lC?W�'��Y�%(2?��S��xē�{\G�����9|����P�{��LWa&#��;b�6gh�exco��e��4.#m�c$%���g��������#h��s�<ak��F��^��uwNR����'*�y~izј����Gà{����aql��ê��~������޽����vO�օ�K3�;$�����Y��>1��/Ku����^���FĊ��Z?�0�쟠�׷��n	76�Ӏ圠�͢:��#D���ݽ��U�[���
������4��v.~?��	�F��*��bU�c��x�ub+�Ջ������H���ф��F���n+&a��s���B������L��a�G�(A'/��G�oGV�a�:3<+�lR��C���p�)��4I*S�q����#����&�R��쑽�NVge��N���Mf����3����V���ͳ����:u\r�Ü��L�~f���0����J�RR[�	�u١��zr[ź�Y�N��"B<5#��m-�I���)%R₪�l,����:���?J^�nu��P߾HG�8�2pH0�������bO��UrB�9��F��RQ��}�}An�ş���2_��5h_�6��6��EH�"��h������Fj��O5���b.]C^ɼ�(wm��A�z�}Ij�/���j'�m���Q-��X�)Η.����}J`���qE�1��ɼ�74MN�J��G�H��E��D��|�Ycu�����#l��a��qjv�:�f�C�Z�	���͒닽�A��x]·*�<���xQ��!�W�p?��_�=�34\8��<X��ma&��ѷH���%���=ev�ǒ�#�����8����I挄���1�]���D��R7*��Qѻ<[6l�mե��!3	�%_�)5�-�Q�dN��vLX�W<���ӻ�?Z
��0�}��E������d�.��xz%]�����V���:���j7�E�G�9�LP[�qˍ|d T�O�8���ٖQ����`~k�Mf�&�k}p2LL�y_�p�{r�`V2'U���B�o���[]�á����ܰ����bP����8�
p�?¤����$"hDM��V��������3��?��\��,۪x!G�<���A�K:�A���[t�4H�S��0-������^�x��s���n^0���3?F_^��"}��;G"c��#0��%�x4w�&�E��'rt�y��.nY��U��#{c[��+2p��d��G�
9�<O�W�I��^�%T���?����� Ƿc��e���fk�I]�ʮQ�4���-1X�8����z�Ņ�:fC�ct��<�Q^΋������{W��G�3�, /g75Wb��BP�ZV(�ƣ?o��˕;$T��x�3����h� ��0OM=&�'�4����"E�G޿QĘ�`�ߎ�2Ń������ј�B}� ۆ�o��WRv�$wN��5�Rg/r��)����b�5q�ƻ�C���j�9��3���=�6��n�oGc��.��%�x��J�U�#0=�/�}�2�k�{��)5Wb���^��nУ&��.��?�xå�w��
����J�G�+�*|rL�A�\d�b�ݰv+�J:�$d#���'� ��i�����j�~)a��<�� dk�g�7����?!㹕�{�����o���`�1���;S9_�l��|v��7�敺�!�#�~e�O~	:%^�]���.sm����C;YQ��lɠ6� ��N�߰�8�����k�*�o�+�(��n��%�`@9�p���˟����P��Ȣ�f`���+'������rN�l/��Ԉ��R�`k�?q��V�����&�~Zҵ��C0��+�UT�����bň���Ͷ�Mn�������l�LIϘ,l��D��t�D�b����*�d�ZԒ�����k�μ<�n����Ŀ"�q���Z(�}v��#��]