��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�g�����B9>z���SEޱ\��c�)�P٨V�LB^���l �g��V�P�U���,Dc�ך�9���}8$/��w'ڵ�=e}�h)��8�E�j����h��B�&P&rV�� ꊔ�3�4���Jb���at�$�V</(3�Վ�eˆT~=�Z�Y��C��1dWg"�y����vʖP�ɦe,S�O�5b54�0�TaqЅ�� ���Z㔹#i�p����!98���W�v��=���M}r�y_b?��Y��o�:�EH�im�Sc8x�J<��T����K:�q�E�F���9$�o��\��}��h�a�$R�b_ �5��\))��ؤT��*ڜ��~�Ѷ��%��b#�~�g<�����zp�1��&�s�Q��'f5�Տ��s�wѨ��ʬR�~�a�16nX@��rʨ��L���s��
�&�R��/+h׽�[�����2s��@t���>�#sFuY��vM��T��L��;�N���2sF���o���9ʾ�&�+3��zʅ���G��$��t���D�8xU���������]#ᰯ5�PZ��3��4�|rD�J����'�*���K��F>ܬ�(��pz��^��L��>b��m1Q�|S"�#�4i`D��L��wܥ��=[���'֊��t����kqg�_sX��d�b�$���/ס���3���fA//�l��3�A���|Dm��O*WI_>�
5���RT���`d����>*�7�A��P����Ҿ�Auk�qQ��4@�7I�7�5�8�T�۶�����sR����%?Z}v]�TaKMt����us���f����
Ά�%�umc�m�!1�W�dI_�oFA ?��t(5�����ğ�nSD;>��W����{�`� ;=��Z."��,����(0�=�?�F�!2"����A�#�D!���9�0)�����KL�WZqe�R�*<�'	�K�)5f��E~����~;ZRY4�׿l���S�al9��2��;�Ü](�1�:g��Ӓݓ��Nԥ�/܀��[�֕ǽ[j�=	ٲ� ��M��2V���Ce�o��RpV�
�Aׂ�v!�����,�&�	�7���a�#к�]�|�J����z�(*����S�(�˛�  �������IoNcY��O�q��j������@�6B`�}�g��Zv2�O�4m�=f���Bb%h��	����.L?�OE� �.5�y�
��BY/�g���,3�DZ�(쫆k���	����@�\@nY�j�4�����sI�v����yB1b	h�N��˻���*�C~e��`k6!����HB1)(�j��2}��@ؔ&N���jN^S1e�bY��L��LM
_Hl��x�%t�6�[aS��a�x]�687]�vJ~�|�K�6���72�� �BsX�^���Dk��z�l�[��"&��l�����fo&�C��<?s)�3D{��<Ⱥ2*XOfj`�w���N^�}���ݥ�+�.�vK�`���Y�>-���w:��Mj�?��{RY�D��	��A�t��Fn�O��������'H����G1��Wl���������w!P���,�*i�s맿 9�X2]���R��~p�l~e���4��0���������.I������U4��6���P�uI�A��՞ ����Tܵ53�ݻ�DV������F�oԁ����mƞ�%�8�uC���&��l����۶�Fk�I�놎�&q�+K��e�Ѽ���f����o��U�`��Ov� ����x����h�v���6Ԍ51���'��~�"%ӿBp��gB��3�f�<'�}?��\�lU�e�N�[t�+	�ꮛ��[��1ƿ �#9N���?T�o�Y2�X�O��j��D����sT�u�v� �+���X'�.|81��x�>�{�-5�[�S�~�G����$�~B�X��/Kx���Ķ�����H�q	�`shm��>������
 AZw�bl�Qa[��_�p��]U���A���������j�B]m/PC��Ҍ��PY�8X�'U�wuw)�[Q$��X��\8�w�1�Y�JO�T6���|�F����@�����B���K��aȬ�:L��Aq��햜\,��6j�X�� $�[��tX����D��A��Oa�q�.�j/\����Rb"��8\���KO4�������e��bF⏖�N����@���0ȏL��}���<t�qT���x�I]⥌ X�ަ$0�!n�;�qL�c���ϊ��ފQ!Q��������^�iC����&.�B�0���b�NǠ3���V�ѧ`�O�mUm����Ł��ݙ&`���xjRtێ�(�3����#�/�EV0;��1�r%�T,�����c����Y���iT2�B[A���5��̆���������M̢n�I��]cm�~��ZXd�2���"�xً	'�E��Tw�j�\+!˾&5dWM��JCb�ԃf]�&'ڂ��7��T�$��] ��ïN��N��T�o ^�3oa��nȯڶ��E���z�M!�i�[k��u���zK	G�����Vc���i�)	<[����>�%gyN	_\��bwO��S��Fp0�K�) =h�0B�ZQ��6��-%Y��=ֈT��@S
��^ZB�[Y̧<2���@ePg����NA�j�<�q��#���>ÉK��(��X��[LM���V�b�m�ԯ)Ė'}0�b�Dc��F�km���r���T�0zu�pnJ�.���4T��t�k]� �Z5����>c��e
����l�L�^,w7c�	���E��G��n��c;ټ�����g�+}Sχ�h����	4aVz֧	R��u�<2ϺʁO�xl)� u����e���i�8��w�A����~�BvDݵ`Gn�09e@�fׂ�DV���6��Q�%�:�����+K¢���A�������k�_���E�C���*G���%eU���6m�vV%��
�f�>|��|u-���nM�4�cW{�ƺ�/>E����0y|���E��1�e!\J�����ȁM��{��6����hS�x�U�G�l</�u��t��K~��O<��Ň楸$�ˑ�����d2�F"TL@!��g*xP������U��m��X���\Y�������}��51��l�Mu���䵓��l
����5^��]��D�mf�x3%�}{��E�T�'�yI��ռ��%Շ�,^�tmE�C�ma��XrR9����LDy����7�oa��L̓�iSsH������'��ǫB��K�A�5���3�O����k�K̮X�q���m"�y&��7� �D��ޗtZ5HL�����1���vji_�pBmz���J!�څ}+�!�qvТP