��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�K��w{�E<�BH�a������&�Jn�/I��hK0Jw8��|��^�,��wK'��348�S�mYw�ߏ5�u5MW���1�(�,24���,T�pmV��}T�jj�ܹI����F�k�}ݰe�Ss�����H<�m��k����Ԍ�~�D/dw��Yf��(��D���B́ ��P����aMO��CϠ�Z�A���m\D�S��J���̖�H��\�]��s��_���&�xNV�"�x�q�W����l,")�>�`��m�b� }�}��f;�'~yrtO�FJ��x\@�P��|8����0`*WlJ��(S���~�0o��/�PĠ�Q�2�2��.sn�$���c'�~�_q<�H�Z�uw2��y�;Wn�G$I��TǼ���Ɔ#$Sf����)�Cڦ,��tNT��xUC�|E��k:��+M9�i�A��ӡ�s�[F�z1��v2"7|���9 �W1c��l�"bŋIV��@��g�x�
|ʗ:�^�0��7�ڻ�¿���]b�6j�Hҿi<j�\=F�d[5OmjT�&q1H+�_�M5��!y���;ՁM�;U_�]�=?{��0���1.5��z��_�~U���S�Jk������b��E^IUA���~��WH��^��Ҳ08���^QE*�L[��Tw�*)�'|~"O���:�L�D!wI5����.~����ZN*FEp�Q�Qo�L�Է�+[���$SU��:�zi�/�<��љ�j��Y���hfc����G�{��9),
6��$�:L�".^kX�qqfi�$.��������Y���}Вs�+��8�\z�6�X\N/�0W�x3�0��	b�u	��Z8ښ
�.F:�*gu�"l@����=P�$z���&����¨�};�+z�%��X�T�JfP�f;#�oס��R:8�Y�&��	�QQ<�~�ޥh�kߡ�\s�~���2$�Y"u�`u0�[>e�	2�}���z��zT������S���(�����aJ�J�΀j��#�{\r5�g��]ִW\z���2��P�ѿ��{[�
F�p�Ib��kx�I�h��Kz���j��<�Z��	���)}ǣ�[Dy�KI!:�� @ ���p�	�����؟U.�8
	�l/t�ɯ��h{|���)�N�t���BO���Э=����f[+t�V���wA"�|n���A��od���k��\�n^�(�qM���n�c�%���^�эm�5���:�,n�b��NHH:��Kٟ�{wj")=�i�DԶ�g[N�g���v��E�MkR�43ʜ6�4�N�5)������C�Ekd��X��WL2i��DD�I�����sL �h�c:�D`"��k�c�0�k�A���c���ϳ�*w"�уn�W[��㏯~�G���%�h�Z�q4R�~�}?�P�Ԇ��o�!ok���u�ƻZH�/���FEB�����n��;4�1������f8DOfo�i�����ԑ `��p>\�;��Vb۲�6��$s��E4������k�c���&'.b����~t�׽dke~5�Pp+��^n㔁&I�!z��U�E�;�X�"\T�t	A�%�,ZpK�@�5{�X�E0�I������o��P�j ؃�5�4C�[[|��[��Q����aE�q1)���C���#��7�-�A50��$��^��z_�*bd[8��~����)=5���-]��?�؍�E�ۚ9tsDy}���]�@����W��r<�5ߍs4<��0�����V�,5��*<>_(�g8.�"v���r�YY�ȧ�x�{lg �߀v��0��#KB�H WM�����+i�l��&�<��(��JwZ��B�����ϱdU�I#�	̎C�-B��k��v8����7dM�+40�
�:�L��#��
*x�_H�R�QU�۹3�Am�OY�
O�v]�_�����	 ���l�$/V�n��s�?"Հ�982=�M�C�>�Y�d�Ui�04ANB�;�f�"�4Z�����Tp��*��X���7~?�������B2!�S���ؼޑZd��+��׵m<�^��CK�z�M�'�G;�$��W��H�9�R�H�Gϯ�@U<��Q,=�	�.ߗX6�,���Dg��[��S�����x{}��絵�D6&�8�;ʑ�E'Kt��.�=b�g���	[�k��i ��G��E��s��mK�\9�;����%=j�i�nG��t��]�ܻ��]S��F������,�#��T?��m����<���R���)�R�{��_����e�� �g.�
 N=��P�2�t��X�1K<�g�V�^�S�=t�g�������9oL��y|J���F|2�\�
,4U�f�V�"m��8m���>��"�Y��8v�CM����s����1y�Y!}���
���_C("���2��zx܋B�͜�V[N
S]�/ُ�n ��wʙqG�,e(���A���*jg�$��O�s���r��v�B���	�+��vq�(-����{>O����6I��Q��I��&GY$��ͭ�;ƞc�B�F�6���� �%��o{򯶛�3P+n���˦W�#�wg�G:�+��!��Q�{N.b�/�y[��(I*�g�3~\���OUDbr�T���"��qL%�9�荄ױ���3�Њ癹>���z<�.���Js����Wh�܋� ����)�C�E�@$|J����P	�g�tB�D�0�wb�P|,� �G���Nk9.b��xWH�߬6��S��Z� ̟��f@�DV΍�B~ZyQ����� ?�E��d��
���.'�s�x�?�q?�ߡ ��Ҿ�2���x~蕤^#����b���^=??r��&��=��-἟��{�T��٬�u�eɅ�+��]Z�A��'�¹9/���
�(�v�ch��Ӱ����Y_4f�^e$hf���Z><8^)�%j�k��^��qy��m���U4j/䎏>0g�bhI����8�z�$}-%h�zIB����ٔ��D�H��0e�X�QOi�;�oJ	T{��B������(���e'<.J|~�*`�3��Y��Lh3�;x�i?d�t�)��=V��':/��_��jZg��B��ſS�(����]��FcX�� !ǭ�	��Seiuϖ�~Oq06�氶ݟ
�TKX��f�n�����&Î�� ��6s*�cA�5�ĪB-�� ]EC/�&Wc�P�3Ca �2����ˇ���kӅ5dL�5.,��Џy�58 ���	ɽc�q�Y>c�j��y�>j�qP�S@���)pRP�~�dH6S�������B�/������̕Ï�S�h�06_��ȼ����
���q��� �o��;M^q�T��\N�z��F������p�~7^X5N�5�}�� �z~vâ?�z��;�� �������:P3łÉ��K�Y���M��G�Z������w�[�d�c��v����"X��z�:0��b%M��P��ե���Ryga�mŻ�/�.�LZ�P��u6��=\�]��"r�AB��� ��ɸ,�������,�ŚK�t)�|�zh��&��~L�6��`$Ni# /�S?�YD���`��XG�?B�g ���n�+�Il��C�yL�'�;�N�L=����|+�&�L_g�N�j�����٩$A��QDf�Y�4�+�ׂ�|���S��P���^�Ԏ��!��*�E�eא|D�%֟z6��^/�̪��eEq*�Kԡ�fk��?��}Yz[%g���0�n��OM������~��&� �sꇳp2,�ܞ���1��b��	ߨ�`'
-tݐ�?I�3��p�=lϡiV�G e�xB� /�J��9���)T|�ST/^吊��{57O¹�=��"�VM� :�2���M���gxl_�%�$��c�=q��xN=���w;0�8��pΖ &I�Ŭ
�䕉I�</z�|.i�<$7e9n1N���{������h�d+m�G5s��cev<>��j���UW�TQ;(�4(%"�3��C�Ppr���y$�i��I���%�
>/�X ))v��@�Q��\���6�0�Q4���)d�{�.2�����'HT��6��0�lC;~y1J2�&G'�r���̤|�+ju0�cm���	�{L*�;g���}��xq�.;�[�op,��05�y���=>��!/��]κ�0?~�3yO�4�7��q��
0�aq5{�P>�O�Db����y.)�ez���'D�t]�4���]���m@����M��̭�ٜ�k�*?�l.�ϻ�J�%�hy���ۢE��x��7ﶂL�M����_hP�i�S��fll���"5Wj$S\|,��4P��,}m�����Y��S��a�"�%y��w9�f��t��Gjڹ2�J�H�=�l��3�>��}���N�~��s�)f<Ք8�NY+�ڍ
^�P�m���.)�᝖Y��!����Tn�}�
ٰvyL�zLKVz�_@���c�1��Gf�	
_� ��d� �jn��/�!J�T�Z3O6RkfmxfJfBݨ\â��j�����->�O�@@�_�;m��\�-���o�]-,~��O��w�u��zt�͎x�~HL�����|4�ӻ��)��zn3�����/�Fz)Ns�����)�H�o Z#�ܟ�C�Gi)ߒ��^N��{�j�q�$YDJy��%�$Yc�5�q�S9�8DP�y����5�T���L	���k�L`Z�VF�Tѵ4�{k��X$��Z���u]p�*�2[I�K`��k;����)/�߄J7�^[�fܮբe J���.�0񑬽��tϟJ��I�2�P�/<����5�3П�y��nW�b\��Ƨ�c	<�6LT�Z�#pV�5
2��w�5�8� �O?�S~4��-��R���f��Z��A!S1t��w�R����0�60�_�#���<Όmv��W�u"�l�m��(Iz�ʓqQ�s_�����ɜ@+���⤞���&�T���ܙ+0������c�f�p�p�����LT�I����� ����EV�o2� z��R�,`�뱣,3�>��Y�9ܑID��
� &�k�篨�bvx��'����oyw�w:p��ƿHTq��V4��I���j��XT��r�7K��i�<��̋��(p��͋�>#^��H�|�a�ç
j<�Po��t�9B3T�d�N�n��N5� ;�)ͧ-�,�W<)���b��05�%��t���	�D��Y����-3�])6I�c1��FSɢE]���/C��\R�ⶅ��6��7�4CG)("U�$�'�f���FY�2]����;��d�aj.�[\T�ʔ�d��J��g�	�w�+D�NF��f�i:�E��留�0j�"�/��xٔ�t[ͣE�c-/HzRy,�T��G���������/�M_1S���N��	�F�󯇿}����9�]�竊&]����arv���"��tGǋY��'1�T˼ِ�'���Lqyݤ�ȵ���!�V�i��Y�2h�K�zW�;�\⫃�6M n��~Jq�8�Z��9�E��Q[Ŷ��V'�G�"<�$M�xr�EG	雜褻�i�[.��*� ��qRcϘD�pL?��me�E �+�>�X��g���H�w��j�������壁�(^�$K+#6�/8e��_��S��X�eɞb�W}��V�:���?�J'���
�1��2�ǆ�E�M�XD�%��?����*khr=2;AꃢP�����Ō�z{�*����5����v,�#���GR8��,6��e@΍�'������^�IfRŪyf.���&�7�,Cfc��Z�b���w�����[Z�%'h��ˆt�I�:u.3�3↣=���ה�v�Nd��Jg�}�%�c㘿^��gtr�z�"n�jq%h���,{B�t����a�}R�u>ڟ
q�"ඁ�ƣ��/��يc�w�(�I�pF�[,Vd�iX=��y�|~��u����|�7��