��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX����q:�}��d-3$��_Qǀeo�b I�jA����|���ߞ�	 �-	!昕��k2?|�$jE`}��ч��Γ�<w��m��r�͛/�,��?w|�@(W��!���S>\�o�����ʆ:|KŎ���^?�L�S��\@��M��/|$�]��'�l}���~Ky�{92q���Sy�����U����⯎Z�=z��=>gj�6P'�a��T>������3�t�@������3ό:�+��C�k;�`G�|ݢ��e�;�j��3�/F�����c��y~��0�|��rVj�%U���L �0K�m����J;�s�x��{G��4ʹ�<�\�L�k$%am\�GؔҊA��"�Z��"�n���}2U��(�΢X��W(���y�??L�X������Л��	��	=h69�4����i�`��k��!L�N��x�9(b?��r�~�L��(5>k������t�7D5T��*��c���A] ɉ��E��;㳧B3��ͻՊ��������>����t����?gw�a��!��|��q��q� ?`��Lg鉁������T"�Q$�����1��g�Î�&�¬�@�?�3��X�`�/B��̸�����7?L��_���V�[#�F_k��:%����,�`��Z^\�<��}�}�CKDG&:�ȑ�v�ߛ�ot4�@�<�k�lQ��@���ݜ����h��w�T�BY��kAgRI��$p��6�M����ä���E�0�� ���_�Rb]5�Rj����z�Q��}$K�sZ\�� �=L�>������G���j�V�Lx�^�ӛ4͑1.�U׸�R)�F3�x����
�?�	\#��1��^�IW���&vt����B}�.'�������� P��Ns��7a}�ܴ��H�l	H=��y��"`q�M+������ fsL�g�~��V���e|>Lj�*@7���;2u#K2�kj�~ɆCӎ|���E�D��N��v������|}v���]���Y��5�V��[�I������xv�\�ɳg�)$W�GjkXv����]�w��������!X+LX�FW�U�M�h�����b1k�v�\��,֎��9�2a�k:>X�\(���^��}
�:Ye�/֭gb����v�Iƃz�������iG��ֶs��a&`�K�7���fR
?Ԋ�}n��5������S�-m8��� �i�D�Zz��b&�^-B�1atP"2���Ŵ�t��� k47�j�mD�\�Wq-p�=贕v�&��S�FS�Ħz}�b.#�N9Tp/"���ދ��֚b��X��>�R�8|2�$�5��se����#��Tp��#�9`[M��a���e��c�&T1-�BB�4�>B7r�ǽ��Sl�>O���
‍&�.�uYӽz8!ܜGH/E^�����z���u�-��r�*ſ
����r���L�o|�.�H�}���t�`^��=���j1�0�I��H#�Gdl2����댓hA'p�AD�2�<ߜ6�����Z�����ھ`�l|��p�w�[I�H�����{L�=�/[pԴ� �i��]W\�	��ڠ-��������A!�
��w	L�p�٘�C��`E�ž�?�l,�Φy����.� E��!��=�Z�=H�~�8�:�a��L��ճ+���p瓌 ^U�y}�]{*2⻺�qB1e/�:͵��%I�6͓��Vh3A�
H��mt����?�+@s�_�����拡T�3��1s��]�Ǆ��V'��\�g+�]�ϣPk��I�� ��Փ�jb޶���.�>�6�Y��iO��y2=Jk_>�̖2Gz�Hq�'����'���3�^e�}��gu�1Cn�;��"�w��3�n�~�`����j{}�ǆ?�R������#N���S2B��)���"�����Od��\���P,� �DS���	� ���zV�5<��Ǝ�hW�V�M�ر틺5z�g�����
�?�XaFf����~ޚ#��Q���o��n�|����sp��n�JJ��,GVn]d�>a���}]�`JI�M�P�v���K蜚��-������W��:~��4���d�ё�$|$F���8}������TwR��Kq�] J��Vg��m�*#�(�K��k�fN& �����Δ�\d-�/܉��3P�Cl!�6%|j��䧥�����Ggo�X �-�*ѫ��о(�6���<N�P����E?4L"w�ȸ��A��&"L/1.�bgjZ-��ʛ��xq��Dl�a�A�Ů=R 
)���(>�k�Y�y�~O��1��V�-g9y�����?t���p��G�P3�{�|�� �e���5V����.HJ�ݤ^A{e'w_�9�u�������!(=n�?��i�8)ۂ�ū/凈���j[��HYYo��KV$C.����oO�n]���:�H�A�T6π�?c��o�Q��ՈZ^�Q� )�$)����U������ʓ s
NWU�,>���)���	�wp'?+�3R�vڤ)�H�0�2��S������10�����?�_)��UO��(+�DL�+k��.��{`s	'!�Ɗ:,����w�O܋)���T��G�)����.W��6��b-]�_�����:L��fZ�A��w�X��q�� u?;�_J/3��(Ⲛg��k�<y��a�/����S�=2���x�` ��h.�N\��,��x�	�,�%���(G �x�|VƇ	�ׇ��\6�7�A���&_0��C}�qU��<c#��_�ƀ��7�~3p���D�b���Y?t=J��S�����ۧ7c��������9�Ѝ���L���n�מ��w�MV�W�[�����=�Ll������[�>���~�_�H�_�����9���^��Q9��K!�	n/W��?��#���bt��8�M�sG�� V�����	�&��Ǳ�E���o0��s�n
�\�wesf-�OX�*�3�t���u�>Z��#AN���+{�_� �d��CA���A���O���Yհ�|���A�-�֍n�{.�@�L�A�|��7J� ���{	Z�>�{�E<�`�L�I��1��R3^��(�%��^Ά������*=���m��*��?gq�����a�(�i����ȳw��r�E��#�%��:���M��H��_���V��缠��DA�[�����[n�,ժ���P�b0@�;����-�����A�`�}f�s{��w-0�"V��恵���fy�U�x��`2N����r��p����y&
a���I����5�Ӽ#�9�;Ws#�0JT��(��4�n��@v�%�����z����r��x� h��~蝂۹�}����B���v�{� ���@�`���k��2Z�?�rh��ğ�"0�8�!	��q*S�8&�'癥S��%��6�S��iv��#�?U{��9ݤ+�T��?��E<�t�^^���*���J�Ao�=��]�\X�b�`�%_ �m��(�z�j�|?����2K�p�{�,5�{DCb�lE0�t��:�?(h�2yP|�:����R����[�ml�		&��D{�9E��_��T��^6�'TS��|��P�W�🃵�.G��E�	vO�D�L�/��=�"+Ƈ�x9���{
�鬣�����s�i�o��� �^��S�Y0r6	��6��O�[R�ݹ<aI��c"��f��P���&��_����� ��b�JQfC�h��F"sU�����:���Ju3������e����f��eM2�y�t�k!�����y�g#�{�`\���0a���rm�U7.iPl�mҠ�]�:ǛlJ<h��n�ց��[�s���8�*��T�T���`̪��
eF�x�(Z-I	�v���ȍβ~9����2y =�yGg2���26�\��>lu*�]��F�Ȏ��CV�����@N�����*���=;���pE�'�)�p@\eD�(�&�����n:��W�1���Y�|�UZ��>�>�P���������KE�X�Ə�Ó�}Ʃ��(�˘
1��,�ؖ/�X��'!�i��>�(KϷ8M��i�#|�O21	�{��������_�KUY(Z{D�n�6�û{�I������#�[F��k����棽'?�O(>E��%0�qpɤ�*��:pɚ������3�+�0����?�RI��Φҷ��h��7	� ��"�.���>n%5E`��r�łyi���1ڤ��#���uz^yR�φӢ�3H����]���I�Z���b_�^�x�E��\�^�/�b>[��;��ƁF�$���� 
� 4a9��jg>
I��T�������UOo�n�s}�S�m���T1���_�'�g�\Sr{��a�ȱ���������?{�H��W�RFm����@i��V�[�j,c�E@!U7r�&��� �&���)l)�-�Xz�Ɏ��@	py���p� ����+8Ɔ,]�"��������cp̈��{��;p�� ;����ꥪ�����-���j����l;�ǖ����׫�A�P	j���V�b���t4�Q��;���
�"��oF}�
}3ȰV�r�T��`�d��!��l<6�ۜQ�?E�:��������5E��Q*�I3FC��	J4�E9�k����a;t'sPj��Bo86YC�ui)3�O��I��>�3:z��]�K_�i��l;,�0��"��)��ѤN#�{k.�[�Y:����� �g�A��%1�q[Ӗ�#w����x���#�O
61��H�\���'t�IЬ6�v��<
�3�7P+Н��ך,�%{Z]n@�"��?�3�'j�Z](L���s��+`{K�N�!0f�׶��s�n�e/N�t���0�֕@��_���e.K�G��_�+�_}�_�I��?F�6�B0����,"�U[�w]�l�;��:粊����|x��	tt�����.�wz�d�'���X�$l�Q�5%4j@_[o��m�+��Yl(;�."f"V�(������®�&	k��S�̻U��I�j�5����qʙ�xl3;,��@\���S`����Gx{��żL?�T�ɨ0���p�<8�f�ҩ��tW�n��v���8]2���J:�d����d���B̦@��#D�i���\i���,Sş$��x�'��1�)����\w��Ic7�������iߙZ���W�g�M��Vz��(éR b�ruq\4��J�?��o����ѐEM�P�+��<�!4��.�V�k��M�.�Nd�diaطt-R�P+�#��aU��LR#�X�'M> ��z�!]���q���T7�=$�a�*�n�����,��m~RN�{rg�f���_Dw�k��h�\��a��}kBɺ�[:�G�#2��ψQ<z��%������ѩio��Q\���T��T���|\ ~B:q�CKz�!Eսv�x��C]�$�S�e#%Lύ��-9�ku��	,0۶ϝ�M��P�4˒��꬈o���;��t@����d�ʸl�-q��Z�|��<`
��T`�}�C�xaS's��1X�XZ��=��&N�����y�ɕlu*�	���Q�]ȩ�����d�ej���j��RLzڂ�Y�c]��>�����6�Ti�	���9�FB���٨�����@����.�pGEr�l��v��&��*��A�� cl�?����Š��5Bđ��'Ą�Iג 5I�i
���#��VpS+o ���K	ȟ�7x��YD��pm02�����'�e���]c,�N�8���!FQ#��KC�Ƥ�ƨC�֊�V6��-��J���0�е*��tm�j��D��;Xe���`���r #�������%�R ދv����)iIؤ�����B��q���<�2�� FO��1��g ��f�X�VX�[2�#����+u\��JFU��.�&����B ���\\#qŐ3�&w[!��N���h%xg"/7ؚ���ߣ��Mf�E𳁞�a��f�A��98\�7nQ2�,�c��dD�d�SF�y�UJR��$�0*�*�^� ��]�����s�?I����y�Q5z:�af��&������i�����b�gF!U`-?Y���P��p^	�8� ht���U��4�,�
X���6ʲX�{��	��&ց��|��Ԧ���KD����H���[I�?��ή�~x��g^�����Vz 	�qP�8z�ʶ�Pfii�]r�x	"Td2�YП�,n[���p>�����A�Q&cb� ) ��dK����k�k`�?Rڈa�}!r��s�<��,������Vm� X�YbC/�8R���Ȕ\ҙ��@��8��e�"�����
=:*dɔar�s����ѻ���â��y�
��`�j����3&�*�I&e0W=�d���p���ҧ��;�q��z�KȒt#B�|I�t��ˮ�ýj�2*�W�4�#�%c��+j1�pb\A�ϙw���	�=5�I>A�}���S!���:��R�S������� �m8`��"���u�ٔ縭���qÂ�܅/�����������W�5"�|
ؽW9�h���=+�t��I����z���D�úV�-�!��y����'ON�bش2�ME��� 3mg��������7�zC�9)<3���L��&Zb����k3�k	���<D�/���#�5i��ŏ���T ^�HF�m����K��-�D�\:��vf7���qw������������nca�������_̕���F���p��G�>��:��:P����F��P�{P�w7�)�sWRະ��4��V�w)\�ܫ�|6D��*<������w��p��D�d>�O��s�[4������,�O8,�Q�>�S�<�,͡g�(�s�^�Ya�t�}��	\OG��<�������o���%��/�CIٜ���{�֎�I~��[ �HQ�PGθ�_EG%P�`�D�$���q�rW	Ǚ����HTX�l�9�*�)ʾ�r+�T
��T�;Z�˺� �[�]�@�����-�8hJ�Q�֎Y���������aY��<[����ˑ-��L(����J�_U�hl�v���Α���;>w_/������T����{C�DPX�-m ܘ,�A*}z�V{np<�?���$9��X*s�V�=���V���_9"��� ��~��'�&��d. ,��Ѷ$�H��Y����l�ʿ���r��
$wΉ&I�r1�n:A��V��S���a��b@����&w_aYc�y��4�Qk�砅�G�-��9�Q�F�s�/�%�	֒����O6e0�9Z���.�8�uQ��� {�~��㿶}h��<�p���y�/��5�=�����#����:�I6)A�Ҽ]��<��{�x }�;�p���	� RY��G�V�^��pl�|y/7

^��{��N��7���͹G�Z���!	��66]�g9��}��������7�����y�r�(�琡��=߲$�a7b a�sز��~��h]g�k��D<`�Wz��"08�����b�]M Ӌ��Y�|�ޔ�dh�P6!�ڽ\��d����P7�X0'Ь�&��A���\٫�~j���2:hf���|j�(-vf͑a!����X�U I5I~�P��]N;)Vƕ7�!V�q?��c��n��p|��Ut]���c�`�;-*���Ӄr��H��41��
�h):h������9<P���|�[' �O�9�B�|�btQ�_"dٿԌ���U�O����D��n�Q�=��	>�0
O2,*�K��uU!@ �9�m G�\��.�ٙʸY�÷3����$++�����l��o?������$���[�B����/�ڿ��#,���1�(`6^R�`��t8T���א_g�ȭ������~�z��	- �	9�Xq�r�,7��<���MV'.c
(�u��X�|�?��^��}1����/��i���q�����͗�9p�c���q/��-���\�匱嫡�Xt��V��x���m9QS5��2C��0վ*���*���h פ��ީ'���Wo����B=ɼTْ3�) r�Ӳ��(|[�L4�i��Ȩ$�[�4�l180���$U����Y��T���eY\��j���i���s/�.̠x׀�����M(|��J�@ZFM
��-�~�0x؉֣��g�W4�N�P�wL�r�<<ш�YŊG.��k�%	�1eF`��
۴��}�;���c�1��c��$D�L��>C@��|����i	��+5��ҳ3B�� }�"^�;v��\��ڥ�D����>��A	�q�~����<l��ۨ�?۝10�<7�����ˈ��(�:�D�8�� ��os���� ����1�7�n`9��6\�L�ሥ�4sġ��)��8�����5��6���G0n%k���1�B8d�G���vƮ=�ɞ���^�4��K.sM�Җ���cS�_��`�T)6���;�&��Z��BY���׷SV�&N�TK�-�hV�q��[��Δ�ł��-�;F(�ކ��%�4�ɝ\D���]�㬙"�z��]�{��'���Q`{ga||mH��#7�L>8��0+::Y�6k_1jW�^vlg�E�zN�?-���4�����δ���}���Ќ����8+ċ?mL��V!�X���h9��1�k�������*8yU�p�-w������,��À2���%q�+ �r�{Ѳ�w�cta����{4��y,P����Q���<l���OE�?4j�)fl�<��J@��� �
��������D�N�E��6}kzn�����ت����*x�p���;T�vkbR�0�@�+^@�z�O��{������$���d2f{7?�����U��|a#W��E,!��@{��
*nϺ8q�O��cp�Cd6��I�߇����N�A�]Nh�3��3��8J���gUS�EDL(��!U0AaT���(����N~��O��i7Kq�&��������_���G���{4�ο�=��.�����`�wG����T8�u ��� T�P�:���v�4Vq{R��'�j�u���"�iO�s��P^����C�(�M�i���hjȚ3B&¢J�x��]o����	�'o�m�G�kp_X<Sn���R�?m;?0޺UK$%�� �$�p�NP�X����Ż��)[���[vE��vpe�/��������R8��[@rn�h��f�2r������lU��&�Tns��?�������}�ֶ(p���a&��g�\D��w]��m�h���k(��7���E[j��+J��e��v˒_��TS|Sj��wE"_\4a�7��0���j@^������T�y�nhڿ����8kH�)�}�����1��1jgh7ɥo��K�Y4��k/��Zm��JM�ww[>~����u�2b���w⣂�aw�[�%�Y�I4������,8�	�`!�Z �i���C7QS��7~�vY	6�$#�GL��Z7R>ꮉdZg�)Z�P��@�F"J��Ϸ���0C~QNnw��wDz���>)�TyD40�x�q׸E\�5�ġ?r��J�&��L����-ѕ�9��5�Q9�V�3�(����|�nK8�*�?�QV^=�#��II�y^:��׶j���d<"O|���M������[�>��&�����^���p t��
���!f�QT����V��{~��r�Z{�Ax��,��m���7V� 1���F���g!K=��g��Rָ�y�m�tP|��P^	�W !�	��n65+gO���&~O_>��j^T\N���,J܍���W�I�[��,!G�&��@Uw��t�{�-bр��7%A�t�V��h%�E`��P~��j���~f���E�ņ|K���=����s�e�N���+%����Q�5�.1ݨ`��7ԽB*�R9�~�����4:՘���_��OŒ<���I�����~�
[��|I��m��'��-�j�1�[?������9,����#ɶz���Z���jo����O��3�Ǻ�[Q][?�L��{|4�����<�6��K[�X�GRE�[�}�fz'c�n�����e�sEo���H��Vg�,�ɐ�ô���͉��~������֪�=�׾���ޠ�V�5���ywr��37FcلҒ&?!�ǭ��
!'�kp�7��G��GqHd��]�[+8QZ���-,��j+�U/0��n�X3�7�/���X�{��q��ff���.�1��u�$���r�h��r�[���b��]��ߒ��J�l�s+	�k�{�n�d��:�E�	�oE7��9o�d�E�\�� ��i�r�:�sº��C��M����X�&�I�ʷ�%��;���
�c-�����wP؞?t�XA��v� ر�	ې��d�P�ò��O��?y\6����g��x`��N�kS�	�8�OvT���CP`��Zv�vV�v�Ҳ۰��/��G���'94m����V'�a�6M-�w�I3fP3����}L���d�Fʔ�Lץk�q��)�g㫕�o6]7��fX��2��7��g�%�އlT��V������� ��Ɇ6yHW�K���*�#t�,�-�LHH-��XV���wZ��-r���������Éc�G�4���Gb�o�7��d������~2b�i�����ޕ��XfHD=�4�4<��ț�C�~����y�}�+H1��*+�3�(�Q|��Qϯ���hT�:p��	>����/�_|l��MR�U,g��i�)ȣ��ӥ��V�H��yC���1�#8�hǶ� l���D�ͩڰ�N���t���Ҳ�c��h U'|�U��I�-�Y(UO��ē��rp&��a����L$_Ƅ���� �u�^ HO�3�g��֩�gӞ_M���X+{�<�F�`H	1ģp��9D����A�{�/�g��`Z}�ᠭq��ɵ#�TijԤ�tU�R��[�ߧ�����=����>q\�s�c�8`�$;�JG�S:aE/y?|oܤ��{���A�0� _A�7�h[( ÐT��)s<��,yfTMrQ�.
N�A���%}(ux,�8�D��(g��޺xJ�E<��e�&����|h�7���V�n�ߪ͊$t�.�')�y#l�����9$�-ڦ��8�;c9'���A�-a7������J)K� )ٍ�|<���M��q�	��G��S:>����b�X?�nS��IP'�#���2���Z�����w7>����rѨ�q'�_P�h)\e�`���̈>����F��L�i����6q�O��!�E�y�g����Q�(6�pݣn[v��U4ܠ8��ɉ
R����Ke�4
ڣ1:)\*咜!&N��ȯ�|�1��B�e��P��Ƭ�4�E,u��2-�*������a/�7�\W&b.����k�D����[�b�S$���-�3���EQ�A�nXgZ�0m�$�I��L+cd�A��jC������5q�p�nŏ��|YTJ�R�'Q�?֗ �J��x�f�F?�����F�׀�!�=�7C��m��FC~Ο.|��ƕ����9r,�4�:CO�����~V/F���ȱ�Z#�O�P��~I����Pީ��?1��<XpUr�#�lH�N�Du����Њ��Y&��W�� �[W(�9x�=L"��3���w��F�P�d~�WP��������$qS�t!f��^W��%���.�mP�]m��f��\��&a!�W�n��l�i� ؠ�� �D�J��k�<�����z��9�Q�癩A#���UY�t&�����ƭL1�D���J3ѡ�k&qX���]ý�Cڋtp��x��H�I�� zd�i����f��2�Ѻ8�;b-�i��գ�`Nr���ₔ�ċt�o�R䞤�|/�H���V�W��yz<O�ްE�XCz|��.I���+ 3�Pb�DL@
�4�B�����ے��*]Jqm�G�_;:e���P���4�dk��m�2;̞�x�[���-��5�7+*��z�92%m�u1�j�=ZACuAV1�w��T���M?�1�О�;9��1-'������m��|`�|ص���v�-��N0��'a�z꬝�G�,ߨ��]!Jھ�\bEZK����W�b5˃4<�? ����8��Ak�݉)��`��~�u�I`��^����uP�+��kG1����Y���W�i�^9���@�)��[#\,gS���N�!�@�l�]���Ŷ���%��R�����婓.j�Q^gg¤�rv�H�u���A8F4� t�=#3��jX�0jd���)r	�p*P��~i�/�~z��`���f+gRy'J�aR�6)����oT|j"%�����NJ.��N��Z��Q��ۃ��6G�\8C���#�Ze@8��z~��˃��]�A�y�����S�Y����Z��
��~ޅK�R��Q��g{�����SM�5���*��ǟ��
�_{-i��T����O���*
�/zh�����,�(�;��>��l��</��Q�Yu��Ԉv�)�Bt����!'�[A��L�loS2\z�/���]�vx��<�C����9[�)
�7��B3?��3���q]���ٻ9��1/��ɢ�����nJ�'Z�%4f-a�w~5"�<ƭ�@�Z��c��d{N��..= �<2�}n��EJ�c������僟��	@b�����E��&sGH�-���*�}=�����)�+�\e[�
�}J5�*I���ˁ4��h����0��/�K�e�wy�Y�Z�O �;?�oT;�,z*?��4���fL�Zz�`@�1��Ò�<�TŰ�nCG�zT�Z�ZO�=o_fqL�Z2�n�e�q�a�VO���g����a?Xj]X�M���qG��1eU����wꈃ�l�8�V����e���5$"�+����\�]��b=���� ��+x35������wb~�v.c�`�A���[�x~������L�ؗ�{��V!��%}o�C7ɝ�?�j�0����&�%"�$��oAyj���8� �rM:���6G�֖��*�n@W�4�����oca�0eL�Q�Y�du!���w�}�7.�;M9o8Q�O'Q��S4uA��QP��ޅ�Lp�i��4���l�S��'��GKJ�K����:ܿ՚|"޴)ri�����Ubs%g���L,b �@���D�����N>]R�����|�7ke���|�A��ˇ�����d����S;�ެ+�������lF���mVe砘S��(��;��'s,B0�Y(�d�!f�*ˢ�h��j�E'��7'�6���e�a~�yk���#���$npfRV��l���P�$$=ݎ�[)�	50h�^'ϊ�\��Y�Z�D��(E��o���R����ӏ�vq�K�,ޙ~%�����A�w�"�ix��2
7qI�c��p ��ꥡ|�����Wm��w?����긲���*�[���O�����#?F��$H[������S��j����+�0cT���vq�.��=�S\��UQ�	J�"��Z����G]��aE)�/� ������ι�����f�8]H˷���+�|�U~g�I� jr���M��(�{�T	=}�@�<���������~PA���^s�ֻb���-0�E���L2R�Σ��[���ںJL��	7u��<ց�cχ�LmZ��Gx�F�b" �oπ�w�0Ό��c�s��,�fلV���iC#�<&ȡ�'�G��O����M��	���� ����4J�������]�{��D����~K(мv����S@5�M���s��a�s�x��O ��`�S���F��C��C�;�=��%hf{D�-�v'��J�w�i�$�k����!���[d��'�xzR־N��<��W؇v��u;�F����������fF-YgВ^Vŵ	Џ��ҝ�� P�
�<Qy5 ;؎�Cc���yY�`�ng���ERQDQ�e8V#]�6S�cWI1^����d�������ՃS�n1j���S
�hm��mqM��X�d��7޽IS^k?�0a��Ӧ���v��-�A×'n��Cq��10�e�3��í�!؛ZS���7�U�~��j�^��u��wG!U>NE=,��yqa�*�<�]��p�[��X��Hӯ���}�E"��t��F���a�)BX��2g�=����j���J�p�J�)�fd^>��m��#���.������17�8;��E�Eh�ڭ��D:u�t	cT�����S�x��+g,���=���gU�*�-g��`��M�B	����h@�T�n�;Ej�-"G5��E��7VT���4� Ei��@�c.P����h����_[G���n�~@���\��<�t�w׷�m4^6	�O�]�
��XW�,ʐ.�d��@�:lx�v�gqo'����6�:cEX`:aڦ�M$�m�ʡ"�U��=u�y��NJk���)3�:�s�Ձğ�A��`,:�ُ�����M���Ԙ��8�Ls!J8�? I����<g����&�M6�3A��Ř��� ��o�T�{i����TF���R�/P힘�o�y��5���ۮM��%+v��� �������R�4����h�u� ;s�2�{U��4!4W��R\#�2X� 
d̏�8Փ˦]�ӊ���pT9�z�@�F�R��E0��EC  =�f5�_�}7x?�X�3��^{�I�������7d��3J�+s��M���.N$��9�n�
mFa�y��VG'��b�0�xЗ5E�����i�[�H�=�uI�),[���r�:C�T��ñz�&zg�_|l{ӄR�����Q���g�H���򒀬���I���#�+$Ll)yL08�^ ��Jq=��C J�rP�-�$��"��(:v!��j��8���	J���y�[ҙ���5��۩A���VX짺��aS���w&�LL�;�*=�'�m��P<�����ϻp���Ai��V������2n˅����t�ɂ�Z�)
���;�@���L"6*�B�)�zZ?�\����Q��h ���b����O���%�F�U�w)�_@Z'��VS�R���1������.Q`U;��TXG�AX�d����}WQS�����U�T�b��-V\�w�1�(�����s�+�4R����A�&1|�l-2�y��x饀�U�W�1��d-�)QM��:}j��(D�$"�ډ]��<��x���=�R����>�|��	v៝��9}o�͈�׉u#|柟	?�z2-���;�!��KDo��5��W��^�ؙ�h��C��b����i���>4��Yx�{�9�7a����b�14�*�A��0��ð�l�-9�%�m~�H���I���S�{��f4���BZ�XQ��N9���#�0�8�N�ZR�&�9�>�c[I�ETz�h�K�������t@��%ؒW:Ԩ���_W������R�l�L��S
�׽N(6���n7ǐ��K��m̺��M�+?���Z{���gc.|=J�|K�ùā  j�b��=/5�4�B�^)�v��T�$kN�|Eu2I�8
���*5�C���RT#`_���ϒ�����0����=�w�X�]F9�S?yfWl�2��2T�gV��y�R�Bf�J����ѱܒ���F�i�`O[r�l| ��h��������U�����^O���֤bu�����'	���(�߮�j+�]
�I枟]y���{���<m�1���hŪ�Y�����]������嘠Z�e��wFl��*��_�-5�,��[;��
�p+�����v�#n��GHET)�R���4�Q��$��u4aW�����GA��\~�	&�sK�Uq�'T�/�׃����������1�����*r2~(RI0Ȳ�8�9Dc�̫N]Z,eQ��$��\G��i�b�vJ�=�Ҡ����$�*��mz���* A	��zcS8�I�͊���h)"�\O�.������ �0/���N��J\p\��1_��' �@:��;&��B4zi�h�jJt��iw��bBy�8$>sZ<�z;��1����zܿ����>\���q�M*����rgj	�������=�f�8��~�3t�v��rW~�\�W/NO�Q\��4�H6%`6�|�:/;y�."�v4�<�Bw���=�c���<����$F?1��7wx��˜�o����μ��݁BX$E��	o�Run����Hs��1����l�ݼ�J7,g����FO�=���.�DRZ���N�N۬��U@��	HXW{���[���66|��{��&��*�$@=X_<����FXCc�s��HöU
�c�aOMw�Y�;�̮��91|UL���ϝ�������M.�hl��ʞ��M����S�2�H��dx�`�]�S�E
�IU)�~6��W����!�)�#gKi���G,]ݼ�G�P�=QE0;r�lonH�
�v� ���9Dnϕ���S���_�jSs��$.��:ט�'
H	��9�d��W�q,r�!5e�ͧ2j����H��y��E�s���u��n�8��pX��,��[K�Yd�Ys�,n�����y�\o����q'+�[�`��?��4���L��x��|M*m#�G|�6@�0q�h^M]�Z�����`�ɓa�4&<��?��{-���M'x>��IP(�@*����"x@u9�d>���"��憎2l��W�]'a�~���b�Ա�<W~0��&C�O�T�_dw�}��FZ'������l~�S[
���Ӈ�.�
��6=,
����а��O�Ȟ�_+&Kȟ9*���f����nyЅ���ω�N�K���Э�(���ى+Ƥk��E����jɴ�r�f&�5f:(�;�/�ǧ�3��7��"w�m�f,����%\ܻ:h�����:�Ǖ���y�m�����i�&p�Efzyǡu?�jd�����{�o�"KH�;Wt�VRj�o��)9jJ۱�!��B����@��(<cg T���Sn��ő:���<�:�#S�G��DN@��^/��=ZXKv+��U�Z�_~��L�lT�w�Jo��
���SE.6����^̷7�+��`�Ԍ�=V���Τ�X�����o�J��A\S�1�NU�����<!ުy����o��N#f�ܫ�����e��V�����8{c����)�ʂJƥk��vT��˧]	���_w�����oؤUĵ�T��E�tԫ�hɋZ�~��o�
9��*��K�H�� �hm���i4�1W����Dܯ<�Z�����K�� �Q�̀��Bc�K*�E6��!}r[�$+8UK�FV�h���G�(������x��xI�3�`�L(u�U�y_�%�KPQ�mbI��dn��(������lIo!H���m� glm~-��۶�cM*5v�7&̧���4]�/�i��[�h̻����t�j�g1d_#�~!a��l���ĕ�'����YVX���۫�7~�Ԅ��v�a��	���M?1���Z-�օtc��Nqڼi�K�w3�lSh�0;G�Ե����m85-`�_���v|�"�d0w	Fyo��Dw�̪��^��X�o�p��An�7���c�h*eR��X� �>�tƯE�0a��t��#�V�9����ȷ{���H���r��%i��r�� ��������g��	8�vw��w�ϱ�+����y�P��
���6�x����E�u�a"���[d��H��uP�4տ�w$��	eb |��֟ځ��\]��K�J�X�W$��'�K��e��	����Q�|٩'�����(�L�i�}G:�M���P�i�J�%�N�]��z��{N�6����J�-�,����d��t��Z��R��d�M~�.FА�P�d����9�BX���;��A�c���mv��l�vL>��ҮX�x��H˞Y��QY�0�%H.0L�"F�<d��,;��V�kS#1�,�$�h�=V�>1$��x��3����/b�����i�y&��D
vT� A9m�	,� ����P�܇�2R.���Vu�'��T��1�X�z5�V^m�܌�=G��P{�뙱��l���LC�߷?��&#����W�L�Ja��m2L*�K�ʿG�Ҟ�S�N;ʌ�Z* ��������<�ge��[?:�2Rw��v���.�9�_���$�a��G�
��ͺ��m��2��k�5�6��Q�?,K��(qs�x紡b��Yh6]ֲA��j�bd�}3�f$�[�x��Y����'_����=��x���_<��U�n��=,�=�!��fvF�a�#:~i�![lN:�� E���d��N_Vi��גG����������D]����'��'��FHMG�>lE����0�G�9��@)��F��FK��&��ԛW=�Db0�$��T�/^>�^��PV8�~kרz�N��3�O��>R�R��i����~��oDRh�ZJKda���e�'%���^V2d*^*�k}�Ty�Ғ��/���$�Z? ��G��v���}�~YI{�m��FT��^/��I7�$���w��\@�/'�?�hAV�?=x�����]o�=ŏ�>�<z�g�>Pre2
��������׷J���Rz�w�X��F��P�kL��f�0�D����ȵA�����'d��v5:0
3d��η�Rn^#p�${�|
�S�5W�Yp)-�إ���|(������}�m�\������B�0�y@�;�{���!AJ����Ԍ�2J6;~�%��Ϸ/��F��9ț/bҋ��P�A�W����L����N����T����2s4ϫǰ{bQD,5.��8�8�#��}��N��Kz�Mx�s�N�%/؀:�N�)	�&��6<�@Hz𨨠m�O ��{;[��fX��\��� �敪=�u�#Ʈ�;���4�,�L^�E�"(�*���0�����ҽ�M��ɜ��adj�h79l�s�l���"?���˙�E���'��ű9�ߣ�Z=n� e�f- �����D#jƻ:{�WB�G6��`��=�ף~��V���!>I�S���=��j�]	�?6pZ��g8*v�``����OEpB)�DW��$W�h��U<�[֌�Jjƙ��|�He�۝��!}�{ۏ��m�z���j�ZJ�����cz���f8���&	���b�Ek���%d_�����k�V��LW ��07�m�S�����(���N��[�\�uZpرXlʢ��	!\����dX"�g�i;1�ؙq,����)�ZIa;R��@�W�d�Z<�ߧxv)> ��x��g��T�~C��Ɂ�X4R2�O�=$���$8l����V�b�L�lIy`,Y�������W��O[v�Ao���qT,�8���#��]S.�0q]4:�+u���'x(�oV�L�_��� �&l�S1[&�����diӜ��]H�b&��T�sZ�W��Y.�@�f8/���R!��"�-^��X��`H�DZ>�"o�}K׵/��v�%���I��`*�ueH��d.�"-�&���3�_Zٝ<��S/5/o����zP��b ��X���gH�@m21s������0�{�J3���C�Mɿ��V.O����d��ܠ.['�N���̗���(��K����s��3;EB�s�j�I���4���^\�^��c:?W�2ǥU��5���������'����{�G�[*��\5�P�H� ]0]vgH���b���3��!G!�;J�9@�l.�c�]W5�R��M����?=��j�)R	7)2Rw^dNr��@�]{���-k�^��|����I��~7,���Z���Y��2I���:��s���༯-����ӟ�G�}1��������>� ����q�*�����ck��(
����!�\OX��C����e�Ⱦ>�� ��S�:�?k�n���!�)zqCO���>p�7r�Umc�C�Ü���gORD��a�w}f�'����M�H�'�4aX^)������tNT:�X��^f��P�$���G|�?���m��4/�5�,��1��{�M�o��tc/�yD9��ݝ�>H��<�]�n����}zY�l�G��X��4Xc���T-R�{�Op�QX�5v���f��X� u�y�v'W�s�n��e�^��^j���kd��%'y&p�,?=;�B�)��mh�d�J�P����E� -�E���TMZM���	&x^�q������'*RT���6.��U��Դ�R]e�q�����2��H�&t0y�6�nU ��WH���͐�) P/~�9AJΈ�9P���Ë)a#��h�'�Y�u���f�o�S�&����rl(�q�uo�Q��uF?���h�F�/��#��h�K���Dhf�6$t�૎Cr�>r������7hu���r]M���z�b'm���a��8�ї��Z�@�9�2�#Z	@C���%�¸H�
��s��B�"Pj|	���SM�i���QU�b�!<9�@�V}�ݻD�Ub�8=�)z;���ͯ�*�,�!�[j�n9)�t(�`�i���6a�ʵt�ۡ��S��&W!���m���pb�b���+O��mT�}�]���S��n���4�aÄC��������N���ӱ1A��t��?o�-���R,��Oz9���"��ŜAMz��I�-_�Z�+�	���|o�o�T�Q�?�Jg �7FE��_yJMd�d7uQ��9\h�n��~�
���(E��=P'��">�>s�p8�r�E�<�Gq�Ṫbq7����J�g�d����z�fP���,V
&B�+�r,��2����R�i)Y���ʦ���5$��l��x���s4��d�5���PC��B�E� �utVz��k��_%�������!~��e�C�e����\������-
2�&_���!�h_�h} �L�6RQ�����[nEń������r�iSw�W���j�l�}�@pc��@%2˨�j�娠���^���2��v�:�,l}>HF9ДF��.���l|�	KUXCO��j�"EAs]JOÝ�o,�V��t��魯��� �XUlFT]'��A�\�c��(�sݳ�Y��uS�a�Rm��J���(�m^nEr�T���1a��o	�o0�2V'�*�.�]�q�`�� ���*iKO�2/.ϊ����΂K��60ns��~\���:��cX<���_�;�2 �(X�B>�V�.vFG��Cn�c���-��#����?չV�
@�Ez�a�����9 j�)LjT3�S�;���Ą�#&�8q?�+2l�Fs�x�c���mxyU��-n:}=X��rp�l:}n��v�=��8��/ĥ���9�8�Ʀ�6:��^��º��Y_��{=�{>��2%g��������U��9:B-2�t~�K���\�~+m�g�h�t�a��eZ6���#Ë�{���.`��	���M�d���`+�|z^'��!s��4���OQ}��G���}�Z�_̍.��s�p3z,'�0?����ȅ��	v]9"��K�������W^[5��Jo�g]�(����;�G#//�0k����o˗Q�ҏ����'�ZJ?�i�k�;3>����mD��q�ǣٺ�ιlz���6lH&��g_q�L;�3>�S~�p�D ]�F�ȷ����t�Kl����ے*�S�e��7���c�o������߷��V����4�a��{𣏕�"uūnx�s�CC�aBI[\��Q��_H���w��剑����Q`	���v�JYi���{�}�1j�*/yo�bƫO6�5�rS޻�9�+��FC�ʭ}ݗ(F-� ��@z=g	R�7F��p�D���S�eb�U$��W��|�!�K��F��0is0�8��Q^�
>������F�r6����`=y r�r__7m������eՖ�d)+����+=�o���S��c���7]� �e���#`�FY�c��cy<iȬ��tm�m�Dƽ�60����&w~Sn�$�:[�Tjd��?5��}}�w|>6���M	�G]C�G�����#�d9~��,Afe�W��n�q��Y�mC���[�O��c[B�'���O^|\}0IV~,�5�Ǝ�OP/��8d�K}B͉��*s�|������Rү�v��D�\�x��3*����3Gn�rQ�u)���ѧ�y%g�_4E�5��8�5%[��*�����X������vp�o��>&Ķ$ć�J=�}؍e!��V�BQ�R�_�5$_�.�_h7.� ��8p{��\������x�9��2ʚ��<���s������>QR�M�϶1���/V�;J�<���v �-[^)Jy�ïȓ�m���Awq�]�͕c��w����m�;`y���J�����Z7�zo�iK�G�����-���2�f���1�Ϻ�!��2)��;��Rt⽒�0��?{Zt��6���*�������N�G��v}Cg%��,/Kw���е��ѭ�2A���1 �O�E�)��'ߣ�0Q�y����zsQ����*��:3�^�F�����iF����MT���k֊�X��ئQ�B�"�����2aoL?���Ť8oF�Eb�F;��H�������/�����W�]��XR�Ǐ�s�RE�ckGߥ���e+��a���hd�u]��O�� /�n���2Dx���'�l���ۡ�.�.�LW�۔Bk#b��ڱ�����9�E�+��Q�U}��9��zk�lᤧ��y�pv�lJ�vvW�g ��<�p�o}Og���ȕ�fJ*)D�v���x�V%�v��'������!!N�,徇ZTPЏ�6VxA��y�t
cڿ�gI�w(;W"./�M(�騷9���Ywu}R��VM2�lr�u�9���/�T��ʻM�ю��yV��E�I�V�v�j��d�$E�}����ԙ����Bq+��ʬ�(���G�fDJb��!��$ZB��=��.D��7�nR
����8g�#y��9j����0������� �9�2��xtT�>����� +k���v�j�KH��{�R>%��>y2��E�4[��
�Y
�(�(�pP��X1IW�:&��禥��&�����~�͙�����n7��#N$�BX��A!�Mᒴ��si��F� � K�n�������
z�"�O֚9�?�3\Ю3�����_;>�����?c��%� `��E���eL �p��ῧ*�L�Sv9�+��i��q�͹�9$a����+o�U#��E6w/fn�$�l�a��H��v�coh��:�����44�ňכ~@�D҄��V���*�Z���ɀ��#D\��1�[ë�E���8t<�c!�`:�.R<���I57��o� 0�IB��ɪ������x�i#v�N�4��f2Y:�"��Q�8I��><L�t�?���yy�B���+q�[E��F?"�J^㐦�4��D<A�~Ӽh��IUq,̶v��;�Egv��;����2�����cRCH���y���s�Ց�|�u������ŖAtn�4��0�2��l���6%0Tp�g�! �����aA�5�� و��o�ԫ�
���E2�*��`��`�t��|��`;�^B ���	F��?�+�c�슥��T�֡��[���e�V�Mˬs<^��i],"�z��i[�+*`
A%Ms�Hћ��Ksa��(�&�br�AC����k9�u3{��TX����� S;7�-]n'69���Ad5�D�u��i��]P�U1"�Y�e�e�Z�t5�rI�.Mh�������X/o�s��<�9ݫ��e������b��U��`������}w�8�� wYm��QB1���o�{n�]�7��=�1�V]_m'�M����ཝdG�]qn�
kS`�&߁�a�u��Կ�Dk�h���,�a�ax�3� ۊ��ӆ�_���'�/{;���Ւ8w���Ix>�'Gɬ��sOU"|�~�.��{N��>����0{b#2�G`kp�n�n�:����L�YW�˼q:Vb���t���q�P���F�[���m�@��K����WUF��I�)�/s ��~SuSM�H�$��(�i|�MB����~8&ee���l����;�e�e��O�����p�G��nhj�vV�v%(�\�M��{�]6u�f�p����kO>���y��s��k��G@!��V�t�d���E��:���:�D�4ʅ߆j����T�T ��[Y>��X�
0{�$B.D<Ǆ%L��c�H����i'��
^p\�=�Y�m��y�FZ�ʷ9Z+<]�T�4'D��)H��<?��+��;�9+7g��ඛQ��#
g=�=�,��"wL-��+���TO�۷<Y$?#�fj�%ψ���,7�o�0��Ea�Ѝ�xU��3,�/�v&�PYս�BCR��4���̂�N����܃�?�2x�-�����r����@���W��1-maz�Y���1B����@ �-���҇M��@B� Nw*_�8�~��i[Kc:�&�gg'}����}��)� �*��ӤB��Z�l�L�o��T��q�n��9'��4��E��D.i5�H({�,d�X��F� ��O�n0<�^�����G�+�Atrh��9�<IKQl�Q!�w[��bD��dd~����pO�"w!k�.�>efҖ�k/���D�*�;*��'w��.���d(����O�\�WL��P5��������P�f(%��?k��h�X�&I�/3�k�zL�c6�\	�tɉ�l=���*�	D�e�_��ձ�A�Y��N5a�����Kz�4+k�N��Нvɡ��-�mm�O��X������5i�ȶd5+	��"��5�6^�Rb�WM�X���F����JȢ�K6����)̆���nHZ���X������]��%����fFgў��U��8�}� ���3�'�?%�a��_��t�ɵ��y�^���CM�5���`f�l\e�"j^�ò�5�z<[�:C��P@a{���w���������!���vG�bq�,���Z�cN�{���x�{.�mB5so�y��ͅ�O�m��V9���X�zf�R�dW�H
U�u��|Ct׮��*p
a ��n�)5���
�.�H�2E�n��R��d+>�,��<WvT�<��ۨǕS�C�m��n���n;0[{�/8��V�\�,��y�>tvTA���G�vRj�	��P ��bD��R��92T̉.;qK	CE!(�/��%c�ï����mӸt=������>vZeN�-@mG�xs�s��sO��j���׬8�Iߘ�H����?�Kf-�}�d�Nj����W�����JU�������(h�r݃7��?�e�QLR=xz�y��x�rFnî��ڍ �H����N�8C��?-��ڿDi@�������ۺM����}0�x"���\^�+��*�9���W�\�v�nH�ۛ�#:�B,r����4,S��̭4ٽA�P#j&�.�3|M9xLY�� ?)��hΎCy+%�&_^�LJ����pXhP8)���K��Dڝ��c'�*	EvFc�/M@eU��~Ok���e���I��w����?x�_�娈2�c��)�\��Y�W����w��|��������	= ���L:ð���ܜI��Us���
�� he��l����5b@5:J��^�]��n$F�.4��I5A��j���ױ���sf��UO+��QRM�U0-B^��т�����/5$v�e��Ui�N� ��}C}��$�m�JV�O�����w20�D������l2w�}N���o�o��A��R4�"�t�=�����I˾�V$�5H��h���]�>n�<	9��{�Ȥ����|�>)��j=��AX�FMK�j��`�_�2�x��[�Y$f�@�*- ��JjH=���JYVۿ�}*u9r�=����V^*��'@{L�_��pSב��0��d:\�Ո�Ә4���lFo�Ȝ�P�ͪ��)��E ��e	V����9�g����ߧu (�� ¤4Y߾�!b�P�s	�`:	*4T/�`��E�-B�0�?
4âs��^0�5�u;�t���%3�W��8�a��;xS���,�	�կ7U����&�J���*�=����~������+O���ys$�p��k��"����M�H$p������ ���4P�1<Hds�"�6����87^r��Λfy,ZRZT��:�7�m�wPЂ����{���������P�Y�+m��Z�|<E�0S��n\jca9SaWN�v��|s�d|y�G�^�J����[��.B��W'��kATJ��8:Š��N��55�RА��\NU��c��@ӯxb�݊�_'�-�ET��d׶8���7eZ3p�����[�M�'r;t]��̗�]:!b��X��R�V4�H
1��ɱGˌ/���s#�i�#]�� -<34?��{�@�1�]�e҅q�C��+eD2�2�B�S�Y_��
��*ڱq�vJ�TI�^9j��Z:�<�;�VkV�+��/*eI��̛;G�Əm}{�D�ag�==�I�>jϛ��I?�Ă���UWC���,�G�&v^I�L�QN�dŔ��б2|���@	����(��
��u�{h��wzE�3���΋�Ȅ��S G]hv(���C�:I]��Y�9[���O�jWw�>�g�Y�5�HS�1<��K�
�N
���w3�Q؜��\�q!��	HM5��{~�l�s��#�$�����@	�5���.3j����dk�84��yt���D�e���5<Nğ2��Vf">�{���K�i�T��Z��Y�ߪ:ՉwR0)�z>k�r��z�*��PYp=�(<FP����Zk/�'�We4�D6��|�.GJS�{�Mܧ���4��kߘ��@���y`�Y���7����f�����El/�V�7y�P"����u-A��霬b�\�Rn-!(��S��IlX���}?'����<�����K�`K���SW��L��i�-��̖AG2�S����E5��+�� ���5W�L�:�eIZ9�:5���h��x��`����S���@�c��T�P0���0�=2V��r��2|-������=�5�Fe�4�l-��+��_�WX�.⪵f����6r���C`Ro����s��i�;I�x��Uq�ne�Ħ�R�N���jrn��0��#1�ت��O�t��T��Fp8���o� A+T ����-o޴���-m��↏)`w;���`�f�����D��ˇ2��T����zXj,�JV�� ��Y��Xb��N�d8�~Y�2��ҁ�N�ɵ�Tw�#��1�Y��N�����N�
	o�K;��:��M�m�K/Ff�Ӿ�O���Z�DGv�:��n�홲M����hk�k.�,��듄�h!�ގ0�oW��腓/�)�C�
?m)��%�w��f�"w�xF׉[P���)q=5��x��aM��)@���1ͅ�Hv+G`��޺5����4�:J|27�b��KV�h��r�$w��bBs:<�������jD��eF:�D����>G�Ż���
rLܦ�u���q\����P��"��:𕼕��['Xl���&��=�/�P-�