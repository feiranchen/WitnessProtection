��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0P�
��T��[i�*�s�S�,�
ӧq�}�ߥ&CE#����l��m'�4S��8�M/�_mB�/�P�њg�s��7���*�D
�ZOƠ�Z ,<�Z���/� �<ĵ`	oZ�a9 [�4u���fƊ��,�b�p������27mm�J}FgՕ������,>�W��,(K�D=�J�Av�W��̍�0o��G:��� n���iScw�i�Y�e�X�����C�E���o�$����F��/�[΄��(Ɂ��8r�Y�!��x[���?tG<�L0�#{-a��� ���2�DF��V|ح�#�=b3f,��r�@�x ·ק
ɏ��k=��Z(����@��`ʜ7d��$~<��w�.��i8�#�Ų�{<Y��!�b��� ����O��ބ�%\�7�4�$�m���t���Ӝ�Nz����;|TJ�4��A+-��ȭh��\��e1]bU��F����K��%�Y&*�7"��c��8V�7$Wk����W&|�eŞ@��8E1 ��O��Kз���wɝ@:�>�A��q'�VJ0�5�V���aCu�_^/��s.�t�Mz3��=,�8#gfFǈ&e�#�C�� U���HrA>�=�a?�ZP��]�)�}B|&|�_�a��
1�x#N���!��ⶃ��3��U��,0��������@��7�������S1�a�F�|��{�Ŀ΁�l��=���Z@@?�N�
cS��x�e�V5ul$�8�,�*�ӗdf���-�X���� %��)��ArB�[�k���2ءb$Ǒ�"�Kr_ި^�Bn�G�@xXS�>K�8
~̾�|��/�s��I���r�X!�PBnr߭��?��?�	 ?n#������݇39�&Ϯ�dP��`����[�1���("jJ^PGM0 Z�m�8�<����@�����4�.��I�2���,�a�:d�B�E^���ׂB.5[���f�����.�s�����xv:�U����0>����L]��^�Z��5� �8I���R֟�[ݦ{����"��y��)�$�E֍*x�G�_�,��M�"�³g�����r��>A�])i?�E�Q��?��8#j���xJ6���Q��>�~շTALc�8D~�uo�~�\�A����tu Az�F��@��Gc���w���$�_���j�΅�����/�腷���U4f�7��ɺ�S0��VF��U�N�:̣o����"��7�o��A:Oh����z�"�����F��Ӡ���CW�c�`�>�s���Q5����G{���[�'՘�Ql�ӹ�19xB���o�Ƌ�����I7��(��E��I���I74�h3�� �k�a�y;1��:AD��?&0G�0�V��*2�v�i�~Q�O"�s��K"%�Cft�n؏P GL��)�y�3-���8��5�(���	E]_�Z�?m�&rK.Ȕ節�0�v�����<l|�8W)�%;�c�����M�de:=����ڢ�5 �.�z��>F��t���Z#YT� {ߍ۴�n�.(F�T�-�Mm���n}I�~�{�s�>@�q����<�����rژ�:Q��oZ��T'���O`�d�gM�R�k�e��K�gɖ��ɟ�i~��^��O<�5e�Q��7J�эx��rk�����۬rs�^rJ�N����D���kH�-���e��s �~���>A��i���~|�| J\�|�ӳ��e��b�
���NqB�	�:+��U�e��c�jj�$�%�o�1��Kf1�O�W5���m�7y�Lr���g�&0r>��?��K��ϱ}&Ym�s�w|dU�W��_&.&��8�N�{�=kz(�������7d�*�!"�)q�5&f$�����Pg�Ԝ���܍� B��Z�n?3�m3:/g ���}pr���i��PN�j�]QV�5mʋ�_n/�j�����\?�狇8
t�;?��a ���4��}o���Z��#�k70��5��5�@H>p	�H]���'gn�]/����Aa-sA��fܔw.���W.�+�̘g��!�	�����{���[��)�"�[Y9�.�~�y��O��m	�^R ���:�.�mq�H����m��,�+�a�/��$K'v�H�ÿ:�&�E��䍎/���!#ف� ��E>��������HS��Vʻ*m��ұ�Cp��P�=LR]_@M�����]�ĀQ�r���ٕ@I��k���D)�!��P��tu��Z����	�+��}�"cH�i�jV�/S��Ya���r��կQ����	��6}_�&�-	��c��'��V����(���/f-QN�@@�~c��(��HsXUǯX+�a�NK��,�D�G\�j՚[�|5\�.|�	�W�� ˮʩd&�._��"����m6s*m~٫oF�� ���.�#�[�S�A�*��e��D��K(@���j�I�����~��^�8>�:V����g�=��nm���]��d�@>J�m�g����G�{���|��?�;"�S�<7hS4|�0m�pu߯Il�Fe�̄̡ӿ���QJ����M[j�'p�W���������֟�2g�K�9�A�gu�K�����3�]b�/S�õ�mo��2����9?�������A]�E�V��n��p�PlІ�u1��l��X���Ō>o:������
LM/���$�����唴�0֣&<�����N�YWԊG�t)wk� ���P�\�7eO���r�V�U��ԓ���MQ��}�4��o-�_[��S8n#��R�d���Y��᷹n^�3����4����M'-�ѹӇ�ϴz9��:)ؒ���;K�c��9�!霵:}dV��Yq�`���%Bא'|�ډz��'�;�*wmz��������`�!1�/��ҥ�.�G"Y5
�$1�Q�����<e4ti���� rɴ&b��nAh�j��D���k)�
=�}�l���Y9H��p\�#5���.�T�6��Ͽ���x���R��Xr���(�h�k��Q�����־>/M괆p�;�l�F�r8$��3�6�e��\�S}��5� `9���Y�E��8c��"��Z�$��}t�<�.�:�30��`f�?k��ʻ+̆W�K���/i�
��@����I?��}�+a�|ʗ��{�F�EO�
�!�r�6C�}��