��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����S��$tF���e�}�Ꮇ
	����ÀǙ��<�f�Vģp3�&�O��E^6����
� ���%ap�W�֘��Ib:�������ф�h"���I	�JD]�K�A�/�#���K}񃒂�Ib���v��'c�s8�����vվ�9�Z���ݦ�g���􇜃�����zp-I��C���E�l{\�#s��X��Վ�՜W!�HY�Ʒ�!�W�.�$O�YN�����b��H,S+��q���7Q�kK������Ǩĝ���=%Q��Y�
9�%@C5~Q��:�r�OD��ľ�x6�X4�0Gu[��aEs*���-��ñVKdL7��S�'u�7���Y,�����`#�l�;F�q<j��0����G�<���65���)���H��䆎EB�D����8h���k���(P�c���%�������Q�4e�ך�?ٻ������N�ˌ?Z[�u���'f1̀7�K3Հ��'�Vz��MySp��:š�N�����d��l�mv�cb�o�U ��ዒx	ۣ��	H�&��(���Q����6��}P[�5Tko��^
��n	0�"?��7j+�� {����n��9I�:$��(sA�Up���Ϙ8?��:�@��Lڌ�}�N{�&�W�xc���#>5t�1����Kd��(H��J������]�Pp�sX�*����.6�(g3�cq�k�nދ<_>��x�~V�=��G�fdkF���T
6�-���5+��+,D|}k�b@�"�!��yB����T�U��Z�G��H���;K�4&͞����kݓ���%j���,u�޴�n������(\�pf-j���J��D��tH���w�8,���-8��+���j�<@��E���@�Ѥ(�$%l�L�
��G��,p'�G_JÝ�� ���\��1�5�h�ж���V�õ�q���{�aԷ�%ݮwڪ>����d&� ����GS���i$��`KK��VF�M�m����:��n7|Q��6�j[�����gܔ7��moȚ8�M_�0���_���Ҧ����dZ�^O�1�W�@}�Y��6{q���z�|ZI+lcOX4RI��Em0R�~�D�@�g�{5� �c��]�Tu�"�����F޷c�Ϫ2����e-^��H����Ƴm����%�3~�p��`>�o�V���e>#-	}I����s��D1s�3;padw,�KGb�sC�l*6��dr��b���|�>t�Ϝ�� ai8�, m](�'f$��D��7=��Z��E4���{��kU��D��07N\�p�E��Lb] 9+0ї0��?CiǬ�y�@���D���#�<��l��и�|��8�gSkN��*T�ˇ����N��)sc�P�{蛿��6�="��`�kO�Km^p�#YǞ1�(���2�-���^�_1b���۟�??[%��Vx�l]L`q�נ������Sk���E;�9�r�T�U�u�f�UZ[D�&�)0�J�7uKT
:�;�=��덛+�Pڗ�7i�*0+0Wc��}��g�*VȞ�g[|�q�މ������D�`�Tf0O+.�v�)��d\�q��z@N{H�i	F�a�[^r�u<�"�NN�ZG;���鈍�A)|ҡb���q/E
����dF�@ǁ��2#��9W���7��_��/���ӂY�X�߹9W���,�v����k����}Ϧ+v�8ڦ��ŴQ�L�B���o ��;���0k�k7�\�^�8J�>د�����_�WdA7օX�ʊ81�cI�,Â�2f�z�� E����yT����uRaZ��z�MoK��ΔF�d0��B_����D�
���]^>�@�������s tM)nP�YT���;550v�����Z�I��Z�h�a���m����i�5V�i�t'b:�P�wJQ��U��G���1K��dO�x��K�!��iǽv�)�Կ<	�w���5�O�u�=g\�!g���O�c���~n���	?����;�{ Yo6��*
k���Z��{GIȉ�@��k��q��t~��m�^��_�8��f�VZ/�5��u�+;�1�"X��Ø�|�����f�����KEH�e�LI_^��X�J!�g�\^&�*.��;Y�=��d�#7�Y��'6#&1f����\���9C�.YI�ڄx,�Q.��
B�ˆҸ���z[q�p��M� S���$�j�P�,��.VT�y����yfF����U�?!�$b��@άa��wl�b���U*���Q��ho�	6i�V�1(7���A
~���R�8Sz��=ǻ�aK�`��4*����GA��o|߶�S�K{�T���֚*�N����a(���L���H<0m8�&��4%�F�M9F;�U����s���ח;�OJ�= ���޵?��Pw�HY�`�m��'�R>$J�Vu�CB�aEi�?Y�ٱUä�g�#fQ��t��6IW.�R���/�x��Y����RN{�`F���։7}��m���o��T�L5a&3�o��g��~2t�������Tz�4���G6 @����'�׃f�tQ�kX[w�r�-����XQ���S�h� ��$�鵜H֥s����D�1�29E�v,�:\��Bv׷��ڃ�w 6�F	�3-��P[ףb��ShE^9Ϙ
�������33i
m��%������N�u �|�g܋��a�#����4��{��6��������ՕJaٚiZ����I �}�V��}L?#����>:�"��|�T���[r�d; �#�?��M1o]+Bohz^�J�����B�&�UNh� x�zw��YF@@Q��I�ҁ�+�VPG<��XQ�3Íi2=`�$��R��C`�&K��Dc�$�*�c�:�K�Lǳ'jDt@�?�C� ����fn�:J�c�@�{�V������v@�I,>&
� =��>�+�ΚG�SWY�>J�YW>�8U�!�@� c���IZ��U���x+�������7ڴ�]N'��h�������)HjG�W��0��81�C�G���
�v&Z���-���+~�z	^\���K�{����z|�D>\�JP��~<0$pi��:7�7��V��oJr�A7���QF�Uz�����x�A��̋�U��Ϸ�+����s�>c��� )1�G����n�6�[x�z��:a����.�uO��*�?��ݎ�?��N�λ�)����/X4����S& ���+?A(�o���C>�oZ�����m����9��X�݇}�� @%Y�n	�Y���Gj�ܭ�3톶�!q�x�W4޳�z$�P�~S>�?���v�C�D[<mۉ����ە��O�t��-z��㒤 �����=���)sJ����,�(xN����u�T���^�_��c�w�I,m˫��x3��\��/��N�]�t�iCE����H��[�(�ףx�!�{v(T��S��
��<眷��ʲ�be�֫�5/�<��T�}���櫎�U]�����y�Y�ه��/�*�e�S����@�j"{��ۓ5U���ҝ�k1��=���M���E����P��b�נo/���t|#� �������[u&�¨�����f'�˼�i�2������B���%�s�	�������HJ�#J��XA�����o
8������,�[��3W�>xt���;9%A��{���Z-��y�U������[�2�q���\��j<u��>,[��sq~3�%,�޺M�.^����	��!�Fj4�AO�9�¶���s��Q~{� #�!l�����h
�p�.���;���D�b!�D�k[+!ڰ7���)��{�8~���*C��`��ƹqq���2�Ư�Oc:�O��K�k\l������15���H>���rh��ޓ&�U���;����ס��L/�*�s~����w�8G��ޫ��v|�.��h^nIm�Ǽ��`�6��[hG��Fq8vM�g56�r���E0�D
��}>e]#5Li�tqA+D�T���$,1�XG�t{+��S�_��Ay�`SX3�����6��y����t
G�l��.X��dv�	=������$�{���h[���{1&ra�V�B��u2
̒�iNk����7E�����Y�z�Q�t=5kٯ�Oq�K ����F/�o�!M�w���*�j��+L�������g-E2�M�gRb�s*��M�+�Mb���>1����X�R���Ƣu�Im���Н`P��
�eu���4Qx���@�5� ��Uۥ��̜�W��e�ͦ��U��mdycH��~4��h����Pi��5�Lu�*=/~U�,����]54��ь�ʮ���N�я���j���p���V`�F��.z����%ڬ���b���/O����h�\����K�ؒ�t�����)�<K�Pjmy�T6o�<'츾��+.�
o[X�Rl�r�Jzw ���(�gf�q56��Θ⺰_�Po���Y��2�Ի��`���EoL�l������5�UBێ�b����'b�5w���{��p�#]��	��:u]&7�v|qd������v���`��LXϹB�5�e���K��G4�1
�#���2�jq0��K�v���)cXa�>̭T��L淶BGtKg��K5�C�zv7�j6�hۧM��.��+Q;�]�l	RKO�~���F~�/cX-	��>9BR�Ώ@��v�|�i�U� ���h$��9sXsė��G�17�X^s�F��o�vy5R��)��W6�����r�U���&���mb�g� Z��fy��a�;��N*muL\���"�>�6��5O��6-�-��hW?@7���CQ-W�?���/�%y2<���ʤ�i!�ڎ1�%ݽ���p��y:m�L�K��=IlCJ.���a�%s�-ҜM��_2��%AOTM�a"\�DoDc`�؊�0g����E)I&�,�O��� �[�]ѓ-���OkeKL4m�:y�~��>հ�9�s�м�6��P:cƁ�7�sF@����رF���dw���?��N�����O7����<�������ΰ�0_����_����G����	o�EC�S	�\�h'&��tCG&C�odH��YkQ�d1�
���л�iw��x�)�I2���Iy�X��9�φ�T��IG�IY�keCe�[V��3ǀy��0u`%Q�#.�@��3�,ޫ�ws�P\1���`�XɅ� n$��уNULBG�tP�y
����	���X��W�pxn���� ��`	�M|'�:r
>`�̥OZ�Y��ۉ;�Ή�P��n�c'��Ms��6ɼE؝��Zk�~�%�T�:�:�^Ev���w���)j�u��)E���{w��B��>�����6S�@� ���e�U�����G�-!^͝nL`oD�)�����}8�;�4�p��\Βw#�VՉ/����E
�&�HBb���J5x;��D�������Ě9)k� ���"��k�f(�g�K<!�>��T8b��ns���_+��5c�g�q�fY6�38m�θPX��ۈ��/f���y�nY�J���y���wk~�+	0I4,J�<R,���!�J����۲�P =B<�c�m��Q�vj\�Q-Y�����-�M��Ā�� Q������({_�xp|����7�O+��"ȡ�˩CC.z>��˰]�5-��,�U���Ozq�$ck�R]���Z_����ʋd�5/|V�h{(�0���
n}�]�t�P_�cS?��s�7��~>��|F0	�~�+m��y��~p�n�6P��#?��H�m���{����]Ƿu;��AU�i�*�Ld�9čD9�������y����@͟麡��t��-�;�m;s�������{L��Ӎ�3��G�e誛��c3Z���F�9y��*�,�u�P�X�]���U��;]���)o�J�S����w@�KK��v�G�0�ɸ�zb�_jV��7�]�a�l�4�Ȓ��^��\0�����Ç�M�L�2Y�Bv��*~��ϟ(���j����`���+�XE��;N�1$�E+tm��삲÷%�s$�^�K��h5��n�v��A��5>�b���=Ő��@G��ߏ�m��S4n�ۉ�-��������i2��$T�昄�3&� 0&R�~E~�9 Ԩ�+5�*�Te�-�;VfE �N��0���Y�����i���h[@�[ o����l4+�)��BS[�T��w<7�ړv	�-,�1&�R�8J�7ג��Z.4��Bh��[Ϥ���P�!��]�NQf�����EYd�l�f�/W��� ]J��M�t-�iF�E7Jr�5�*2�5j�Fg�Ҩ�!��B��.d����<۵$W��mE�2��(1fؤ����Ӷ�Dc������0q�8<�Zk2���'����ѥ�Nz�к"�K[�@Zs2?�+���U��XT.��/�p�����B�W��o:�G�����ɟ��tS��6���^]~��ê�8Tk')�#D��Y�$�S��'�������$�c��Q�+��L��l薄C6y�5h�S�;�vD4*?�iN��>.i�"d�r,����&3�����gr���ۢ��_@/Λ�)��4�g]�J����-�vf���E�B^���x�\�a��G�w����+��F�'i4��m;��3�!��f��.7hf(�K�:��d�K��עEOAN�/0C+���b���F9���i�~��h��N�� ���J<�;�脎�YE;~�_3��l��X?<�zU�� YĒ=��8	jXJ�|l��*rs�@DTSL4�� oqSC	����� �4ix�����i���[I�]�ނnm�5Xz��[U?n���u'�{���$�:�1)�9n�ȩ��|?�>h�j�r��@贘Ö
m�&��e�=��-��<fz����x��4G�+�Ze����R���_3�������ֽ$��z�1:�Q��3���~$�Ve�;X�&���<�c�^+��#ּ6�BB%yYN��e��y����(K~�IRB�f5g�,s�������/���,�A"�]42���9�3,���n���m��.�H��`�%dR�?�uD�
�A&+Q���6�\��&RRW	�`M�j�m�>k�����+N<�n�����"z��UL��S��S��� ��
�&6R��Q����t����p�LN�6D�p�����n7L��/�~��Sא�!p��jL*�6�6Пe=��7��a�+Qa�����qsf��'�u�v�'��g.�Ҏ�4�d�4���ʫ�.�C~5��*1���w��!6�����/ry�����"������j����C�F�fY����-�f�^�֖���4�R/�s̏�$��%vp�-�]��.���U�R�4B���X��x�C��&)��B��*JR��R�I�6��KY�ld=l6��D�#��*+j8��w�}���Ͱ�	����l����8���J/��K�����\d��Vğ�����p��ʨ�~�X�>i:���f"D�r{���*�m�3:�����c%���6M"}%�fƂ���H{ژ��ڋ���F0��n��x~.��LX>��|�i��Potvm�C��l����l̇ōZj�Hd�,�e���Q1�x��f'��b�i��>��A#=��u�q�-^m�k�;�'�r�V�-�W��h��f/�X���$ցR�Xe���(��&���.�EJ�0���;Tϗ9?�n��Q�R�-[��_7�$g��ɇ�ej���l����'��O�f^'d{(t��7rl��J��
k��'K�������
p����7�G�k]�/"��J���x<$}夈O�O��2�?�9,/��C�S��=�YH��I	�X$1���d�[Q*k��A����Բe�D��˴ڟk#�н���W��;#Ѽ��+W����	�0����`o*N����]��*b��98��ԇ�����2�Gg�m��±i�t�Fi�Ke�U�QNF������A8D��z�f�b�Xk��Qq��n.���,�i���u y}�~���
�Yϙ������_"�����#G����)dv����~�O��a���c��:���,�߉)�9J�օJ�ajE5L4���g��V֙ �����v������cQu}�]�� 3�]����`֜{�}rE��N�l��@Ts�s��7����Ƌ�˼��].���s�ϵD+�E%�N��;��)a�d0�f�L��{�ìR�|���lL5r��`�#�Z�;���E���F�����%e�@��-ZY`>�o��o��&#�$~�h�38�k��7-����pf.�/��Yv�L�{��!7[|ڷ�k��g:��gŢ�T�c��fB�#�� ~�"yPk�um>� %�gLa]����G��7-���>�)eF���]I�㔬�"h�m�Tҽ�YK'�.�����/���Rj�P>ҟ'u�r�ɥ�1 �ю��؄��o7�8��z^����
e�ֺ�� 0��Qqf6����F#�+g��R�|g \�efK�h~���~�cC8������Bl
���v:d���{�E�K���+B�/տ�W������2�4o��}�>�u[Nл�[I�ˬ�?���f��-�	�Q�}לs�bkF�
��%�J�_�D���J���dh�]aN]� ��첱:C"!B<x�F���8$���j�h
����m��Y� F^8��gJ$R~�hj���+D3�n+�gCk�q@S�{?��%����-��ϩ8���v���R䞯���N�\�����[�����.�y�q�B��:���@�L��M�6�������̅�H{.p
QX{��'{"�ԧ����	k{�C���"eÑd�T�V�O����h���A_ꪡ ����5���@������Ȕｼ�d���_a^��/�vJ���H��<�]��>�9[���������ʽP�h�����s֬J 8����k��LH�dUj�I����Y��ML#��L;�h�O�,+��?�?�!�>˙Vn��9�p#( ���Ұ��)�W�er:t��FX��AH؛ȋ��Y�yTZ�@3�Ln0��Q��~�4�t2���d���ﾼC��c�i�@rS"V&��\V�!�d��1�:1s_ǅa�i_��K��pg��Yɢ��D,..��t�B!
�:4�j�sUs���}��IʾSg]1�A�m
���Ջ�G���[�'U�f��ά^�6y�<П޲!��,���i�JmVi���{w虷��I�{ޣ"�z[o�:X�.�&*��O��V<�?5��[����ʼҷ-�}���:�	}b�P��$t5�@�`�];;D�i����(��~�I_�+�,#�t�ݝ%��c��!�A���*��/�8��0xRx���#���8�[*Ƃ,�q�>�(�k�2b��g�2��[��%�����&>Ï��~8|�1u|3�ᇹ�-3'�gy���w�f�d���A[���޸4$�|]�;}+6p�&�L�H9�(Mت�:~�8+;�Q%�L&U��z��7���x+^-zj�'D_`�ɮ�4�x�	�Ά�p}8� 	u�H=�h�O	���mH�Tlݚ˘ӑVWI�<��5%4�[l����7�c�tC#�g?lQ��p���WHUI^8����f�';u��'��XnK�v����6�g^&���|5Y���Z��[��Т��+����2,C�t�%�e�ɷ�yD�� �h�}P=�H�������Q�%��td(�/�x@������|�ڲ��cn=�DD�L��$ֲ�E���D=�� �*����!]Ng1v�79u(�Q�\A(	 _\Y6��Vd� ��>%�^�e\y�z8�� �L2�~^�g�9�d#�D�x�X��B�a`k2nX�-���^gI��V�����2�]���˓�cڮ���r<��QX�hnV������I�|�H�_���N�[��6��"�j���С̯�.��s8pt:	8a����}��J��D{q�c�v��|�U������W��O^�-�DV.8�+i�
!I�!�4V�'��{`ٝ�����Bء�連`�t6.��@
�{v����*��96@jWTkd�'}�3���~�J-�#5�>�?�>Fx2��X��z1g���c7����v@�s7�
�k����
�<>���Q������>������[�D8I�%��@0����]���ܼ}����r*k�JK��E�x̮�LQ�w5�4b~6i��lIꉶ�,�Dq�x��dx=����oQA~MZZ:������l��ɇ��CQ�Iq(��J�����1�g�1�0�X.�(wM#{Q���;��[���-�d�]<`椏Z&�GE�|.�	(�r��'�^��F�a��h�.�BB���}�x��i���Ae<��`	��w8oF�1F���!<��� y_	���t��$�y�L��cϦ���h)fڏ	ם�$���A��6�Ӧ�6�Q�Q��>(r����\�#KMxZ�~o�ܣ�8�-B3�G˟�+�9���I�Uq����la�����f`v����\���&˯���F�d$��ؤ�m}�����M{=�ϸ�Z�ly�ξ	���Id�Q'-&<
*��f�2T��:6�%�ا�P�4���B�#ɞ� ��O]Q�_=ީ�IO����epHx4,W�b�����4�~��B��N��K���cUU��MHh+�{b���'�m��(����V�{s��>5���{���n_�]s-|��L�������yQ#������]~n,8O�z�&G�U��9�aƻ���};�L⼇�ػ�����mj���[�"��)D�����u��I�S�����*��m�x�?E�:3?���[Z9�t_^��2�d������(��#�7 ��,
������a�bk��-(���EGb��h0J��x��t���-0���Vr��V�I�d3|.����4mStG��&i��caC�}p�r��^7��K�jf�G�֮�