��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX���6��E�&���D�.��;ӫ��oT}8V��=/H���o=��nr
uYWM5�h�PGL~�-�������p��0��^51�&��/�E��l1%� �FC���21��=���������3�"��3����u��L�ad��W�&��֎��:-���mZRV;Kq	�Ϣ����F�c¦
��%#���R~U��P���q��D�@`�^�K͏�{��
����H�Hy����Ƒ����1����:r��k�6s��!b^�WBkq}��sm�'�:s����Etv���1m\�^��e&�˭~�SO�S|�Y�h,����/�ʫ8}ti��`���P]j�|ufم�t;�=e� *U��|��|#d��L��C�2��v
ܵ��I���Z��={�i����ALk���I��!W2ͅ�{��_�g���[z����[$��Q�_����C�E�A�ՓҚ�Yn3m�\C��>{$g�l��Iv���g����В��+�؊�?��=
��F��?��-��c՛�����Yl�����|x0;�˹�D�V2�^�2��Y�n���`�F��2i���qm�6]ش0��a��u7m���7/�
�����\�+��gq���ᛯ��{�b*Ҏgņ_;����^�/�XD���U��wr�����}�m�/�����T��(���l8��s��P�|��ǂ�ǋ�_+vy����.��vE�0��p�Ge�h�!�O����J|���#��{�Je}��MiK�����"����2�p�sB�ӡ&�E
�
Ɔ����o��6yB?jeB�@u~$��-1�Ǐ�������)ܪ��h�N1��*�P�!��@�/�H֠F)y./��E�as6AS�Gx�gܟ�bOiϢB�<��B���h�U�¿(�m&��4b�I2{Ul�f�bM�;md:��"{�Я���@d�v�E�:n"/�|]�~�П��Z�@�
X���A�g�*��.�8���h��Ӑ<`���XV_�J��g�Uyp['�[:�>�O�'M&�� �
�&��i�7�~:눐�<ScByL��\�p���$���SP�UZ"R�!��O��w�W�/i�V�>�+s��a� �_>��1�^�O�'E՚<��@k�EUt�Ѧ��g_�O(�АGB�`�q����&���[�E��A��M_�׷v�l�S�<���z�����2����/�.������2��n�
"�� ��@:3h`F�J��#�F���[G *��Bb1�����u�~ϡ,r����dTl���D���y"��&��L��0?�s-32���n"W85h̿ď����~c�N��%�py�҅���]��v�G�k1Ά_lN/�yo�΋�W���gf!�!�t(#�'�8�3 P��ւ�u��[Q��
M%�����_�?��)�tp+��nΔ!����A���lz3$��� �jb��ҥeT��L���ྯ�L@Mk�i3u^L�>)$\�>y3y�(�g l���C`�K/�O����B�J�^�dn4����!����J8�(b��-:5�\:��X��˧�dɤl�e�"#��+-kz�^��Jy�u�	�U�L��l~��6G���K�;1J:���#�����!ʺ�5��ħ�*�є�0W�|�6�䐓���]�
D���yԟ�F&�ufF�k���=��]2S�0�/g��G	3��T�	-g~�<�}<��D����*0�ȏ~KGJ��������L��C���þ��7�%#�/�9o/�����B�-Q1��1��͝��M� �0��Z�j��fK_2�h�B/L�R������t��t�LO�/GuS�Ӣ��������b�(s��5^ў��U�K�G�����Ip�ߋVˆ����A�T���5э8]$�"�O�$�#:����
V�O���t2]���_9Ji��.x�e��'�g�[g�ju��\��7,�چm<�� ��O�,��kP�w��<EE$a`���T�;X��>7LJ�	7rT�6�-���V[%7I+@���G�#I�e׸����Z[]&g �JR>�M�V���43�������NU�|���%
XQ�D�����Q������'uw�Όm.{!�n��t[Z��HI����X�8��]��y��Y8*��)�چ�@��ow���:��*r]�KOl���RA�em�kC���9%Y'AgM��J.ڐ4��l��Օ���1�e��XԮ=�7FRK(�&s�ҭ��)���nJq5 !�֧,�Ԩ�Th�y�� -��9���wYηSZi���K�"9��6����^�^H�0�*Gl�5p&-��q�����P����rU��1D�eRB��9X|���~H��d+
m	[,�}�����ۂ��B���Ie��>�u�)?�K�����ަ��rʫ>Ϲ8�mrI������,�t�T�]K�ve���^�YB��� �${ć��=���=���m�������-�E�9�r�b�g�^5�֯26�O �EG���[��Z���ɿ��F"ˇ%~d��Q��{1�~�����Id���lE���r[^��b��0�r��ԋX��Y$�ݢ��#}f�v����-n	a����rc�uZ^a܅������`�GN��dv!�8$*�Y�����\|�G�wO��x�������~z������z���o�U�7��C/o�tC3���퐕u�n�!���;m<��I�1�Mۦ�2����R���VC)p�Pg�4Tk��[-�Br�dc p��Q:�UR|����b�0�.�X���Z��,q�4�C��~�����
i��k�w���1�t��7�[�����i��<p�4�"*��X�eHW���.�0��L��[����> xW{��kQ1�ñ]Ϲ�&�a�"ٓ��a��i������'�~�FOܻs�`Z�.�d'1h�,�f���B6Oݭ̩ v��I��n�Rm�H�r}|#�4�<,�"i��X�3D�:�86�+��:�p}<݅n̎H@�^ڧۃ�S�H��.�2�z�G�n%�bM.N3s��u�Ӷ��3`9!��-��$����۟:�<���	3�ސ^Y߲X��6Q&�.�X�F�_i�Xx�`S'r���RT��x�OO�w^3}�]��#��MCՎ4�Vዩ�`n'��I��o(����G��<o� 4�,H�o/(3��cr��`�W,���_�1d���mMn�ZK�ɘ+nץ�JԮz&׍5�0?M��EKƫJ�jy����#D�ϛ�UY�}]��b�gbL$?,;M�rx�j
����oB Mq���EXv+Z�k�=�Y&�^��	� ��ӄ/��>��ў�h��e
�n��Y�͵�Ĵ̽4�b
��lsg��[�3e�
��xA��n;5�Es��Ӓ-=��JuCQ(nB���lM�'T� -r�k�"Y?��p��g�������C��/;+X��C��<@y�jAµK�I��͠�F�+eMiKWug��b�<#S�nݗ��捶Ր'�gu��:9&�����~�\�am�j�b��b@`���o)X�ڭU�͑{�=>D�:��ܿJ^�rkY�P�3|ݽ���#zɓ���+�>�I!�Dļ؁J�iy*(����A�rI=��'�;>�+��1�
˶h��4���<+VZ���C��<�7�PҴ`]ZH��Md���a�=�ֳ�n��-�yyy$����}rؕ����ⰸh��/�TQ1��l��2OYKϭ�&&U�� �2��I�w71���ծ�d�0?&�J��e���/X�/�B�?=�5���ew>sV���7@|������S@ I�<PT2��G8�b�!J�`�X-�̤Y8,k�����ˬ�]��s��:�?lD��[e�֟�!0�8�)���>G7�J�}�G�z&��.�kH����΂.�j�+�d��p]K��r�5"�1�t:r���q�od�ґ�l�����ǚԆ��pR��g�c�~�,'�8Ŕ�-�0���~Ҟ�p2q�:��93+ݜ�V�zS�O1�������1��+��C-��z��L���M�OƓ�XH�fEI��6�d�;�`�L^�^�ɔ]�{6fBE�����o������\��k�<"W����7�߸�C�ϳC�t��A��i+�uA��=��� )L�ϻ ���]^�]�4�ٷ}�l��j��W�������rhkc4��0�$	6�Ar�@��_͠Z��%-���	>�ǒ{��V��ڶւ��o�n�SP���r�	���m�usG��{�!m8L�j�ÔX�mIaмۙ�(�V��6ΔC96Rܙt�x�h�����]�f>�$H�z��ڳE�Г��p�(�y�5��k]���� $�:��I�F�C	<�S�D��Q1����K��J"�"H�x�VGW����0|@\䐏_����5�q�Q+����D�P�,�7�,�c_9� T7����p-w�[hcW�����V��u|�3\,�����mRtj��R#o��ly�� s�Aٯ��w�$*z�J�%wZ*G`�uox|J��Q�h�XWR4��=�9���ղ�9�ŚcS�8�����a�u���?��J}7����8fC%T�VCÀ�`�d����u��$�P�rC�VK 0����g�b�=Ql�2����.,��f.d�f٠]���ݻ��#"�����m�ש��l���F�Zʘ�!�+�v���K;�:�h�HO��I���ײ�
h �2���N���W���s�?� pw� ]P�5Ad��(�;���p�G�tb2���>���h�P�ifj��~2�bHy��2��.�{����$�����
tѽ7"k8��S'3�$��V&$ט��-o^�\�%4y*SH�Ѱj��#/�o)�a�z�Է��!����)~X\@W+��Ȩ��~^���ޟC��${^�K;A:5F/�!c����V�C^�U�Ëx6y�Z�^����#f
�����f��G�eV��^����d^\*x6�ӯ3�Z����M��1�xw�/�"Ϝ~�
��Q���^;bzL��-Iɫ�b����,+7/��K}��Fؐ�Ic|�溁���h$ę�18���4�6�&��XjZ��Tlpi�=f�®�b�q��$֣��?o� ;'��0|}5�`��Ztxuf������%��F"�a��X��gj����]R�������L�N�目��Ap*��EL4#j�70E�xR/_䙥&؜/Q��P'�C8�#�M��E�y��?�!�z4>��ؓ�4[4P�'�4t̭��Sqސ�@�BeO{�RuY������pa��M]��*��ӟ�I���F�m���h!Le��I�1���]�F�|B���]h�Ԍ�/��C��iebK����*e�s�/X�'.S܂����M�l�N����ѷ�Fz8�4���Z���^T�����".P՞�Q�L`��dg�-�q�L�u��s� ��g�F�RKD�nf!�o���&�h}:��&�2�P��V$���d8��~�o�"����W��wE�ΘҙaI�s)-B������3�۟>�O�.W�u�B�DY��o�U�\���;�$l�{̥"�<	_�Lz����A�KvX~��W)�9��t�8o*�*�jk�C�������͆�ju���8�5f��`�(��V���D��f��n�v���	RRx��`WK0z��8+���>N*�$a�C���׭%�gN9ہ�cX�Hd�����s�#�d����G�����_�3QL����L�2 U��-��cJ�g�]��Q�p�-M�;�ې/�+����c��f���3��B�Z��ab�XVk���aZ.�Lv39�<"J�(��_*p��x���#\�&IЋ���(�Rf�{�����|B�r �*nB6�	�AMԸY�/ڳ6�C�S���c��Rv�0�RͻE���Xő��J#o���EPB�1gE�W�Y����$�M��~����l����͎�A�� ]��n�/�M�4Z�#�E�I��7[�7��7/`vKߩ�=U|J-��A����F��Zq�vx7���Ȅ�Ft�.�o�T���{����� 7��=�$Eer��:9/3.ä�@�/'�����*~��WY	�w,�gB}l���������0���0�V/�UPX(�f�Z_�wɩ�7��V�-���U�|ny���V�/Ms���m�v�ݓ�W˴y�l�'��w):�qV��9p'F�k�\7�!H���bIk�J|�oꐁd(�Nf����$w�4�z�����F�-(�p�c{)M�~��!�/�D�%Ç�8�q%�nز�%��J�E�jِJ����༃Z�
��цa�`(`(F2j>SS�c5�d���NpSr�� �ꍋE>c��'%�2�o�q�qK�0ո!f9G�$:�C/�1-���9�7�g�[�^`��w�[�`e���[�Zà�T��[�b�59�UW^�\��q?.1z��ϛɍ���L���X!mi�e��,�
h�A�:-�P���4B|�%��輫&v�WC]q��#h���E�?>Uk���,P����C/#<TQ��p�Y��a=�R���]���Օ�uP����]�7�����,Ŷ�G�������A{
څ3���kUF�-��|˽e��emn���S?��6�	lB���;~���3H���}J�S@��½1�~6g���0��y<��|��T��9�SB���:"��z�w�/\��x`K��z��\{.��<!��5�A���c��%nK �c��UD��ol�u�hi�Ib2:��|'��e	�CڋӹJ�p�Fݑ�]i�0�����i��mq4�� C9,����_��PiW�w���AG�X>�ׇ�5_�C����<�Ɓ�����LX�A+^��Z |С�h[��Ό�&PZc<Db�Q;��vz�0�j�E �?����X�`D���\��7�~��G�Sr���V<X������D�&�U3�b4����\�7�3�/P���ja$x�|-��N����	�K��V��?�>����,D��C��7{x�t�Qs]%ߝ":�B����"}��%���3��LTCa"�V"P׏�2�u��Mpaa_@�n!J\�U��$m�aۙ�r8�Z�T��|�ZtM�����76�b������o;�/�����d�]�/��Y�b�r<���г�&Q�Q�������ǗU��j�ٙ��M�$r$s3�2�FG6~k̴;�,���2xa,?�"���M��\~�<�A�����>G��
�B���uS�,F8/����|� ��AKs�����Z��� �3�j$�'��[�kG}���[u�|���R�Q'w77�����9R��%�ӡ�~BG�#�$Z0�B%A���Z���dE$��h�(κ�`��8I&b����o�f_���~[u^ݭ��FLB�
� �sC�X��RQn��~�*��dVApxsꩧbR �{�'	'H��1�R��X���5+.���ֶEq�n�0#��s�d��a���*Wc�EΪ� �|�ۊ��[���7�|:M���Ŵl�N�k{���*d2b����h���H�ϭ���C��0��g�_s��d�p��}�pF&��`D+��*�uj�˵��?qH�U��)t��]��=��u���.���4��x>��և*Ni9r�:J.��Lt��#F�	)�)�m���)v��d�]�[���&�|&�aמ(S�Hv�k7.|�h���Z�r��=��5�ҸZ��*`��O�3�Ѽ\>�ah0f�?!�[�rւ%��f�
��$;�I�v7X^���u�8��DgrK�
�@u�@~Rf���6S��!�&�i�c:��AU�����	�T]�0�U�r���$���~����(�B��x�T��r��Ɗ<�o-1経�u��z�~=�lQ�j�%x���i� ̢V U��n<λo��"=9��I��h �z�W�GW ,�,	&=gnY�(\��F���Nz�l�i�[d��$f�a�f&T��� �9$�B�C��v=3�$@#xNI.��6�6vd����X{�y��@�id���3I�5��~q]����zQ�6c���c������:F�\:��L/��v�	K��|�[��6�Xܢs}0��|ɼ����0�!��>�Ux��n�R��y�H�ޯu��MZ�q�s��_cam$����􏞮tyh��q}�*y R����XQ�Άf�tS���t8���BV��ʽ�Z����Zs	d��uD��¶�#��IW��	� ,.���"�}�^[�bqe,J�B��נ/Yp��'��Pg�Vh��>�J��Yg1WV���eGU�#꟦��	]�Mٖ.�u�菩e���g��7y�+��?�(�V�O/&��Ei֐]7�&5#���ncfH�"��I?���Ra��U���vw�itI���W�k�*��4�#�GB9�h�� 07��G��xC�8�\��;BI���b��ywSbFK	��*�F��"ś����^�V�A��F�H}�;&�����LD)v�4�*�=�P	{:ԵK��g h>(�xV8`g
������t%&�%�?�����Yh߸�'�?=�3��ށ��h��2$޹I�,����å�����Zg�D8ҫ���pU�*x�,�����Ԣ0���_μ��a)xӋ����⬹/�g���d�zs���Y��܄کE.��AY��fX2��mw����l�Z(-��g�-� ңڿ� X�1p�4I]��E��F�� 	��^��w��������W�C�`��{0�o�:�W���,sm�c��V�e���x8o����)�-b�K�K����)R�i�:�I���)g�H�eaD���2œ#_���;Q��ԭB�S�����[��T��,o���~���K��НڠJ��w��IVM��w	$h�7��!�,�1 ċϤzy��&�XF��i�3��_�8���?s��oƿ%��L��	n���`N﯐�,H����r���fApa��}?�`o��Q�����i:�!��1�/'��:�X���iO�m��`X�9g~���"���;.ѻޔ\��jn%�.��|]�������>PX_�%k;���0i���&�F��<A3Jz�����1�sۀk+qL�@�ԈL�H�����y'/���<Y��d1�� N�u#�H!��38�\9~�޿���7(�'p�3!�8Fm����
B��J�Cv��I~aȬ%��dd�ڐ zq�,$��_��SF�U�
����뙲w-Fb��UP�M�g�M�
=WV�Eu�iɇ9�"^��w���_��!�+.^?�[���c���{��*�~��_ٙɿGdBY�\�2b$fj�n,�BU��n!f�o]���	�k+o5 �W֯T�k�X]&�J<_p"�Bc�u<}Bě�|�u�D��0Dwq툕�K\Y�����>�ρdnP]�hƇ��C?�^�ׇ�v�P��j5x����Fk��0���P��m����p�	�1������ϴU�H�y)f��p����O����ݴ���)��WǮM���W;��i����q���B�FI��M0���Iķ�)	�V<�䋸`�H�2��0](}bLJ���&�����a�}7�����ٸ%�܏LO��O�?���c2�z=�)��2����/!�N �v�����aF�`f$�gI@Z��H3Ku����?U:Y�T��pX�)O�M�un�6 =��#�F�9`��H���ע���\_��,�A�bq=K��ؔ>?s,�;z#���H��{ar�<�q��9ha���@�������*�K�(���8�0pɡ�g����t)Q>�`u֩� ��M#�Ը���aC��!�x��>���a:��V���^���y;'��-�+S4o�>�dSDY��&��غW��3�*w=RX��9H��n9���{�iP�?|�ĝV!�N�l�I:8��vk=�1�JDT�ZdDkv������!Ę(*�P�z�]A���U#8�P�"����B�E�8W�{ny���E�S������y<v?dqDi$�qw��w*��x�/,ߐ#�T�Y�vxJF� 칚�?����39�J�D�ɑ��j�?�8�σ��
$�޽�F�B!�Ov��i���er��o�}n�ӆd��n��b�^�/���R���g�iЮ�y���8XN-�I�W��<�]顥wG^<?�b���a���P-�zz�A-����ν�+�A�_V��,�:2����D1)�Z{�5<_�ְ<��
&!O�@�>�%BToU^򭗱��F���Ley!l��%�]��C,'SSt�#�ZdU)y�qԹ�>�=�G��>�Ma�Ӯ
\�pd	s2�g��xV�N4v���G����S���b�b��Z(C���뱯��(��lJ���21;V%g�;[��%�db��(�a����[��3d�h6���mf\F9����
G撏�:y�E@��e�o� Жd�u�y��9:�\;���WP	�)M��\�O��_�����?F(S!�$�����K���xߝ�i�#���Y�<�so��N�@��	�]���2��z�ε`�@�Qu�O�>׻#��)[�����X"�U	�mt|�Y)lu�IIT����z�/���bY����U�ԭ��	�\�/
~4	���Sۑ�g����U(7��3�Y)���`�
Av�(��"�J��w ��Q7�i�9��.Ȥ�˒R}��#�+�ߍ�U��<�.g�y������y�$T}�,*�	����í�����b�w׬��o�d�C��/v�Y�zn���f���h(6CK��8W��^�c�b�?Q�\~�X�M�k`;m��Ud��H��`�N2�qkD2P�V�w��j�;��e�1�)�v!4u���9f� uY�:�%�d�R�|�P��_N ��B	v�@J�!�Ni[u+�:�(S�/��4���ʳ[�U>�?�{����d
�
a%��ž������%�5P@i��4������p?Ib���5���`r�P~�J2u���Xx��lTS��A��B1�H����OX��u��#�H�wy�**i�z
���6�H����i=�O���YRC�][��`�I+��A����"��k�&µ�G*r��;om��"�o=|��1��`���&kv_�8L�5*���͇v�o�ܠ����_��W�����) 0*ZAo��}���ũL7���6���\Ȧ�֒����W��{-����$�޳��k;��,���(�$��P�m�Os"OV�H}$��ꌆ[�4�n������V��K`�MmUl��V��w���d{9k� _~��^�1�<�}iXK�E�WS��եH��ʱ$# ���=6���侓6em�N_���H�QM ?L�����e��̒Q=U��gZܾLſ�����F
���ݛ!*����Υ��A�j�N�M����wj���T1�MN)�i�!�C���Fj�3N� 5$�@?Z2�n����;���?*����gG�@t�V�S�˕��(�#�M9���A�o�����aQ�x�L�H�'W=
�Y�<�mO�Oꭥ��<������� �Ɍ���መ(���X׳�:��_��ˡ��W�=h���oQ�]t�ո�jC��~�G��e}���!¾�.Qv�m���=~�����"�%��GT��0& !l���_J�9}��]O�
Pc�VWf�[\�.S��(�\�8{0v8G����rurZ���Asf�0�� !Ϭ��x��ݍ����]�N8
�!��`ܭiMȰ���v��&Vu�K��,���r�S�x�\p~��>���B;�A>n��! SC+��M���k��b�� ��M|afҟ��6����.2q�9�h��Qr����֋/lר�8�5���u�g���-�*��1%a�6�38�f���_ͱ�$,���v����h#_O[�gO���Cn�rS/H�AGm�Q�j�hC9���捳=��(/�����鳐:��kWɶUZ�~b�ѓ'~���.7�$�Vc��u��ØI�hmf]��� +����(��}m�:�t�������M��� ��b��KQ�þ��J�s�02���Zڤ���`�����Ѭޢ֞w���ɛ&|���ŨFB��x)s,׈L�w4��]�9�_��oH��#��~���_M�?��]Z|�;�{E\W#���b�.UG�*�L�w''��	�;"K�����a���QW	d�}ͯ�VK�2�bk�3���"˰��r�w�BѬ��r������簅���
b�u��w���� �\��SN���S����I:ՆB�;����	[�tN�5�u�j}��1�O F,��q�p�M��P+�t"����A��G�VQV����t�f�h����.��?'���,:�y�d03y��7�y��|��
�����fŎ*6@��;1"_��9}�榏ʹ�1��o{�-�P��~�}:���kR�p���'�K9�lS���X��� �B�&�Đ�^$$��.����ѫ�P�&�tR[�g�-������s�kW�;\Ts�ӳ[���s��q�s����C�!W7���2� �� ���!)�H^�����ȃ2%���	���n�7�n� �},�9�v5�4 d	nM�n�I3��hkL���Vc��	��<r_��:LP�}��3)�4��G K6��a��l���j�<�Nt��C�VFW�Fȍ?��G6��D'̠7�Y���RK�
`/n�t<�?K�[��Z{����/�|��خ�eU=��.^6�=8���%u�T{,��������[�Q�ل��u/�D��ֵ%�d��5�2&�1�B2�����$E�����ZZţ!�=����Ư�H�0NJ�;�+��� H���̏�_m�]���ѐ;�bF����u]���w�ߋ���v��4O�X���ߩP`�T�e���[aహ_�(s����#ߒ�'��o�Ev�u4�B�`�E�S�-�0y�쬽=�$���ȓ��,��y�>)��¬���] qL��V���~B�����D�ωiqY	.)u�W"��j�@6����E� u�}��"ػ����~:Ѣ��m�Jf��C %�q֣pnD E�P�&�H���M�j�|�Q�c0ߕ�s>��m���]1S^<��ɻ�/VV�xm�s�{����1n麅w�!�{�P�[�dc{�7S|EgH 1��B�6�4q#����z��%{*f�I��I~��[�&d}�w��e�E34���L�.���+�X&��Y\p��\�T��#��[�}E�r��,��լ��fFڛϚ�wX��u�nL�cM�:(RjU���Cr� �'F��>����;fy#'�w��[=\Z�ɽ���+lf������f�"�sM��9R���yt��"�f�B!L^�I/ǻ�}	� ����Q�8�/\3���� {:�upa�. O�&G�y�/ɜi�[e&Z���Bҥ���i�y���G�`:�HsOxEV��Jj'2=���Q�I��F�z������r<��,�m��!���?8=�=n���x��Y��j8G���]ː ��6[n�pu�o]���h���
"��C0��h�F���q&�3�������0�aH
9�it@2�+V�mθ�P#)Y#�(�%ԏy�3��c:B����S�t����!w1�/p���6|LU�VG	&��~f�U�^@�]G`n	�#^<[�i?����t�U������Ŧ�l����O�=��ؠ�:]�^_�]�[��1�J�r�cd�dd�/U�}ؙ�!�|�Ȕ�J=�a��w�3�˫�J�%ۧzV�ph�����x�%��?%�\��@�����]���gmF9��	Ɛ����f���� T+�c�G_ �an�>����`c�Wct�jw�q,�j	eY����]��@�����l��+>�b���]\E�:��g�p�<}ӗ�E�Z^	��Ð�4ΕS�����c����#p�/|5�S2;3r�'8x�����c@ƯZ�숤V�F�˛������Sw_��>ַ�8�d���<ZFc�KP_b܊G�@N��ll�t^ϑ���b��H�&�����=f�`,�G~N2U���&u�'d�>8N�d�خ�������!��sTR?R#ڳY4bL��ʲs3yO�`v�Un��Ȗ�=_..�S8��)�w�c(|�Q�kr:�s������74%��A}Ǵ�أ(fbE��>�+_����N9�7)�		�$BvXzN~��fa)0����6p*��\9t
\|?1@p���(�At|���D�W��s��`	��u��p��k듃ȅ��_�np8�pu�v-xӋP T�܎B%��6�:E�d@��0�\��>���]�D\���)���e^���h
����lbsgMuR�Y����iI#�.��"qWI�8�S+���{R�SЗ,鳳	��m����,�jo͢����4r��)����Zc5I�~�,g��I����˕��>ʘ3�ᾟ���fɌ�:f��AA�XLF,���;� �s�닱�x�.X$��)��Q�N�4��Q��w5��aZ�F1TY�Ҭ��s���6;�acQ֬��g�?⻦��w��x�F@ ��R�?3"�Ŝ�kW-[�sn[N!R^9vV�`
C�e�{_��3�0�2+(��&����=q�}��oݽ�=E s����������I"����4����&6U�� G.�j~,��~?4�fo?�b��L���ie�*뻩"}�M�b�����OS�%z�����t2�J���(�1Ia�N�T3f�x��� 1�C��0���I��>&�<g^����YXκ�.���0�yY�����/��`�"��L`zH38���/��3��LK1�÷b�p�� D�"M����hږq��S����>���2C<���.�KL�1�?�]Ц���֫Ed���g�5wb(f^CR�D�p]�X�+C*�-��=W=	�VHp�g��#���2ߞ��M���T/ʃQS����)�;�!%�������H�ҵ4�P���w�h\�+�|�q����| oN�d������9�&�X>È4�=f������8����q�F-���'�U�%���J��?���]����<�n����d���Pb���>rz�?fvO���Y�����o,�����&^RM��b&*�rU�ܶ}���XVV��J$n���&:"���J?�v��	ST�Gi���M{T��!�,O�(�	5!@ӏo�=9����;�!�2Z�!H�rE٨[	�d�
�u~^������:ַ�}�xi&�� 1�����Xuuf����A�P��[A�Wz��F�n�8�g�0tM�@B"�SQi�+��`%H��#'��t��e�H6����)�W���z��y���4�Dp���[������e��d(n��!�V��b%m�B\�����F�d��h\�*���I����Ign���k�痏���a*�G�l�Ke��4�<����4���χ�W�7�:IA�{�P)|��D���58A���vrW�	��旗�;����Sߴ܍^.Le] 3���^s��"������vXc��7���KE��fN�Аf�O凿዗zS�8;�>��`&j���j1�Y�|��Ntx�Q��!"���='�x�-oR�7���L��?��ٹ:^Np����ѷ "dt8��I��8��y�-</��	.���8���v�╹6?�d��ɱ߈���>���=�׺O����Mu-8��7�Fz����q�/�[&
�O����*�|�ui�@����Ik��N(d[H����}T�E�K�.
ˑγ����Aw6G����#�.v�������m�j�숑�(x�U��DW,�R?B�ѣ3��,惉]�>by���O�Űv��4�Q���e����=��B���J��j�j��������*�8)�#�>XA���%�O����B�;����I����n�C�+��p��&���T,$�C'HWLd)N���[�u\	����Y�������xq' �N0?����Pn�T�TVxb������گ���P�ާ	T�t�G�&��4������v0�fd��C�<����&ˏAKl:�������I�����,���UH��;.� ϭ<rxŭ�A}x���O� #\��x){V�����3���������	` d5�R_�4A7�)�f�D���-�#�G����"��!�7oD��Bq#���cwB�@iw�}L��*s9�׹}���Je$��
ރ�쉕/����}��ߊ#��e"z&�rlC+���(#��޻��Im�'��w������%�Ԧl��x��:�y@�3Y���G;�!&�PG>��8�]B��89?\�P��-G���F��k�	iʾ�w#O�o��]R��3�3�z#n l��؎������{q�g�c�\�ʡ�'���08�S�w�.�'	��b��=�1�<��A��?��	�(�vvB�'V�i0o�@9X�T�WPR.>����DG�}z��̏&E��$��\��Մ���M��!Y"m'^�C��+ �����L��-��*J5�\�[�j2�x*\S'�#�uI�$E>^�����](�s��+���Z��������W�L��o���ͦ	g�$��*fI��>uT��3)R�X"�<^�4u�_#��{��!�A��!?CR�͋~�l|F������3���NE#HVe�x983Kvqho�Ն�<��QTW�C^�)!ݙ���d�V<od=Xkt�*`��}P��~���6ڤ�?��)����K���j�� �f���_�:�%��Ǳj���K�E�`a��9���|�z�Ҋs���nҳ` γ�B~�+�W��T .��ں1/�T$�/��J4&| �@V�p��L��]�[�WQJ<�b�C��J��8%Y��T���(��D�@��;��0�`׻�i�%u�?� >�B��P���Q�56��i���9o)��$��cr�R~���;���4b�F��/�����t���6ߛ�)�OzR��h�� eS6�h�Y�ˬ�b"Gi�.��D`o�,g2�A�'�>Z�\���]tNL�=��&�O����w���sB���o���-��S�"�����W�h����|�+��\5AY�ThZ�'���rEw�e�����U�\��|�CN��2tR�8ӹ۷%��i^������ځ1��u�I�>��wǠ�2AX��+�t�u����ۍ��'�T���z�.4�=�_���qD�Hj��x�n
v(�����껤������=��i2A��L�KN.c�,l�&^��O+��-����a4��,��٦��k�
`Ź ߗ������Y�wFO��ʂ]���9b� N��x@�x����e�\\	
R��"��N��HZ8�D�c���U4S��+j�������ƀߠ����#��;ߏ>�hp��U�ǇDs7͈����:O�iw��lEt����*��Nl�4HzS������a�M|"��(	��,��f��w�t�?=�w���ފ��l((�B�n��z����AH���eB�R؎��|���e����Wl+���\�rI�M��L\��-����$ <��i*F,���ݿ���b�C#��U����T�6�r��ݘY)��S��"��:>�����Is�/�Ax&}��������&A�'��G�4����;D.�)-��c��kS/��>ʝA��Ɓ�_d0�^|-�W�f�.h��/:���ڞF�LtE
��R�/�}���Db��T�f��e���2t_��-]8w�A��V3����o-B{�f�W�놎{��+f��*\�Go�����6���b݄�CB�\��)]Q����W�ڿVJ��r��ʌ J﬉�\�6ֿ`,�S�]<OyXފx�[~����س~J���Scavo+/?��v�v3p��
?��"J�J1a:���W�KP�ʷ�a!�ˆ��L�b����<����{��$�*���
�� U�*P�[������6^�/�≀�ʈ�T�H~+��z�'�Y�g�������.�_�� 7V���\#|���6��X�yvAe����/��b}�Q�:Nuy�^���O�K;E8
� d6��N=^���RF����l�8���fCn��#$X��'�SR����oގ�Dc;��O�=]'Tȩ�[aj-a���/~H����Ƹ.#Y�'O��%}}�v�Ct�5��S$Qt�Zs��.��8n�ȹx�Q��àQ�A���z.'#bD��A�t"y��M��`'��?��v5"���d�76l��ok�H=�E�,_.Ŭo�#�?����`�G�S��ӫ ��z[kr�2���	�Х;L�x ��Wc9��)��g�JXb�ʆ�Ʃ�"�� W5��K���������	��d����PO~�]܆�?)��h1%߬q�@HK2%)����f��.�h� �D���ζ�k��D�h�a�����.��zD���!�1�.r0<�e�Μ� <W��Py�hdh���jz|���.[�p�a�?ض���mcВx���L���"/GG	ם�\b��x��.%VQs��|��R.�ڢ�`������΀��O���F[�@Z�'=�$��p6�_��h���loC��W�|�����W#��?��1_�z��`�S�
DR��J?{iy~�ZA�je�OjbK�����(�	��ג�Y�A�[Ae�9q9bTǔ�P���O�1ڥ6jp�J7�����r��gI:U:!$/�[�Q����̎|C��:[�W2�~fP�8�%�#N�vi�� ��`:����ٛe}n����&.n�U��O���������)����c��F8��U�P��F�2d��m$(�nI��O�%�R�S* f7a�8E�E(���*�CW7G�k��j�����a�E{�L[$�YN8�$?袃g' ���%CH,n$4T��ly�2;�l���Y��xǦ}o�ܤ91�;1�}���KMC�LdU(֛�[#��L�1�~[�B����a*Z|��9x������V,	&(����B������*���r�~}���A](&'��< ���R��/��L�Hv_t�U��斛��n`t���H��/�Z�S�ПMO.��@bڒ�-�_{�귣�n��)�ѓ��_~mh���C��Bz.��	��+v0����#_���4�G��VM$\�W6	nY��_��@���\%����q;�����ϲ-�����ߙ@e��� hX�?y�yL����ҋ�����^9��X*��s��G�j�ë���: M�ɳ3k��������F��4F�#�W=ػ3�D���($�c���fZ�p.Fx��Y��������E�2�Zli�i����J���d"_�,�Q�C'��0��K�Ћ@�$�����&[�S�ו�D�r"N�%���o�(�	u�l�0r�'��41XG0���R�D`B*�?!p�ॎ�~���q�9�B�8CQ+��ʂ���7�H U�� ��o�w�z<���Z)07�*�̨-"���ҙP �1��9��b�5�$=ح���Ɔ`f�Ebڇ��z��X�'F�yӖfj�o�+�Õ���#�Fnb���ga�~7٭8#�#8#:��o���1i�vl�ҙ̢|���;)Z�6�{1�p�T8ͺ�����9�g>�ȒD��U2h@cF¬c�n91�&Q#��0�&���z� ��X���J��R��gvR���|�N�	�g�h�t�%����썎�q_#�yj*4�����5�{ph73��M8��u��9��g�ȸ���9��e�9�ݔ��k����螎�A\�V�������ظ�ݝQ���������X��XueI��h����p������$�Lx�7��p��0�������Ը=\����Y"Q��^:��#)����]�����1)�{���7v4��a�T��"?X&���Q�R�s��$���
!���a� l
5%|F!|篳�a��Z�U����gI�)�`�㮪	�`�(t(����Ц�b�����K4^yMP�6��`2+�E��B6LcV<��xo�P��G<�2��_�Qc G@���<�YO��B�]����_��x�P�>%�Ipr�Ư��Gvr��PXH���z]f�s�x����`*�k_�Q8%f�"ҞSm1�.��-��sC����7�(��M�7��rEw?��O�9�u��.��%,�$,p�_�O���Y+�����ԞI5xJ�ء�\��yA�j�̙�'r]�	l��`:>�i�a4*>V
�yBn���>>@ؒj~m�N�Ԥ?������;hݖaA��5�ԫ�̐���{��jO�	:2 �W�'4�z]�]���'2�:�	M�A[Z?HY�\�ZT��C����y��`�WjF�������tb�����Z�7籄�ފ��,z!���1�����'�6�=p"?SO��Ej�,�n�.�Z�Z���r�b��.jo��H�Et�$P�f�d"!s�o?2�qo	r����]��&a���?g��(�,a��?~�Av9aᐜ��&�Y�U'�4�x�V>i!j:\��	���-��Pi��^��Lcs��� Ûs|k�,�fH�W��vnk
��IfZp)/r���PoG��-��zW#����L>I��^,��_�,�w� $�Q����9�~Y�-|z�3Y���7��
a�'L}F������#oX(�v�8'X+��w��ǝ�w���do��@��9�O�ن�Z�>��o�	��e_�M�SO����� v�]-Qv�r�1|�^1h��ƨ��/�g��d 68 �#�L,pg���)�*M`�\�g;�9S��\�,���s�˅�7�:<��1l�t��ș]r��޶��P�R`����sW��h�ع��1�3�&�����̫���Kϡ3�l��m�J�2�t�{s��cl��M�'�V��
�o�|���o�X����&���O��f�c�o����'�&�A=�bG��nO&�4�X�k��cv�9��^iKC"��6�+���ޟK�9�&XU	sp��:������/�3�u��R%"���{Vb�H��%���@K��$��H ��W�m��uV�9�ېM��������/�K�!S�c��+/v�/�a�3����m�$�&�q��ϼFJ�����7b�ï�	�g�|ن	ކ!ՋP���%)o"hd�� �L��9.{�h|���'����w��;�3n�-��[�'��1u�!�1����P���~ίK�_m_�~W�:q�w�	�=���Z��;�T���2�N	�����e�q��{�F�tn��{�'���P�j��y���Z_�"qo��r�̬���\��|�7Bi���w:}x�5%^
���˭�)0��WmNt��3Ḻ��$�� ���v���h`"Y�so���'S �pR��s�`Ijg�ʢ��ބ����:�弻hg��&�5�Ĝ�H���0t˅s�F��a�	�~�4:��S�O��j馭�⤵p�s�d�B�1�
ZgA
�i�lQw�)�9.ǂ��=N
���L6KR԰2��Uȳy��	A�ԁ#	ެ��y�]�'?y�g&7��V�02�X4�~�ʳ�ȉ1YcW��B��r��_Y~/׺�� ��Af׾UN,@����wW
-ʯ�QX~�w]����M�U��t�B���Z�b��8��'T'M��V�{k˦��nN7CJ�(�s9,f� �P2�l�Y��u�̋��h������%;N�6%�t-h1_VCPLSŵ�g����-�\��L�B�m�|A (q�|D�:Jb�N��$	�s�6�����-(��\ܧ��Ge�X��m�z@��ف�U��u�{�����`j�K������8���p}ŧ� 	1�����-�K{q�3.�Q19i��R��ng����G�!�0)��x3��	����:���ν�v¤fک!d�DI'RN~��fW�l&ηY��Ah�*�Y����I�e��؉�+��3�cc�}s�rVY�~+�9�G)�<6�I��
�B�̆�m�!���I���ٰڹ{�"yS[|���b������x��B���7�K�zZM���:�	2|�$N8���>���֑�y˥ȏ��`���yS�������"������ɑQ%�d��)�� c}%��N�ʗL��l��$���f��p�`�S׈>���0p�
O�ܫ�^�c�>M��{���k�ON�Un��Q�-!���$��W�B�6��&�`�	3U6z�L[ݯ(�F8�������3�*�M���pc��5b�׬y�/:GI�J��+��G�̵v/x}�	�x��4)-�rc�ׅi�˽�U��.�m�z,:�Z�,-�����3p������Rh综�X�i^��1�bϿs��pkg����T��FàQ��@OTR��_�QQx�\h{^l�b��8��Վ�?�h�Q����c�̘jD���ĵGH�>��X,�-�&�d	����8Y��C,��B����� ��L9��bK�}�!�)r�2��k�� =ߞ&u��y�����<�{����8��.+�M��.� ��Ď�D�E�Ɣ"GP�1N���Y���1��:�3oz�����5�ϒ�����y{&�s#�>4���t<�49���<��O1�Pa�"���*�S����Ed��X���٦�bA~���9iz�:�E*��4�<��y�g��Y�O��11�$�[Pz���3/灒�NJ�z`?���i#̣��?Ę�OW9��5{�#��~r�Ibi�Y�8Ƞ ��8�P�c�}��łfX�0��o�5*.ʬ9ıM��g�E>ᬐз��=+�P�|ݳ�Λ0�g
�}�.öڡ����> �ɔ���t�$}V�bg�����j����V�b//QD�Ś���6δ\�c��bᆣv������>`/���1R��T�m�}@�Lw��֠��\Z�����uc%|;�0!�ۑ�01�f�W4C�mM����%�#�ጹ��D����X��b���tN4I��)t'{�>� �)k���A��؍
f�,��2-@�i���:�oFW	���1�� .vjQ�o�l`:�!�%����J�熢U\f)@B`D�j3,�Y^�v�x�!MGmy\w\Nح`FŃ4ҹ�u_Y�J����¡�aI|�M���2��C�I	~2�f9	)@�'
r���}o��RE1Q����L ��d��S�8_��N�	IJ2�3<�XP=_;���Y�e�Ichp���(�LԦZh���]e�xg��#B�4�S��#���KT���V���W��d�Br.a7�Nf�!d��&���U	�:����aBo�� ;�#����7L����#�,��J�-��!��}�je���gOG
T��&�Ot�wI���O���.��󅊏r��j����e�p�~�>��>/���	�fl(�5�qU��8J��N���~gc������2���#Х]Zk��$�mW�&/t��`����-�������<�*[<��v�!SGפ���ZKGF�u��D���@�)��Z��~�T�N{��\��Q�w�y���g�_�9�\��d�j�����Z7z��Y��R�`yk�z�׊�� �RŠ����D�1CI0�{j=���M��N�@�y�ŒJ���Qb�����o�N��ǆ�؈��no�"k��7%�f����K�$����e�z���Ez�}�e�K��@*	�CG/�'X~כ��`d�1�E���^��:�fC�����,�ݞpzQ���ѩf�Ot�T� �OMU�u����]��X�:3D�O��R�!��R
.A� wM�aS�-�bw���5����,�ڙr6���fR��}Du�A��7���É(��>gC����8��0�mԪ���|�צ-������'@XH(K��#k�s�Q&&�s�Y�8��w�����`e�$�� �r����2��۽�Δ��׭2*\`��o�ͫ�,,�z̤�����+�t�t2�-�@6V[qB?p���T-�mgrc�iȼ���B������4;� �D$�^_��C��qbCSf��ƴ�Ĳ��Dp�~V�:�����������&����V�6FIͽ� �SB�n����*�l�^��4��e�tl�9W0T5�	�} ©%º��J�*'jo!rz��I�o��ʺ\�klS�G�����X�Z�L����������s��C㏛^�����k�Z�=���H^�2#"ӅV�b���$�HyL����P;n�O/���I6��'����M!x���R~�W~�W:n��uK�La�9��fT���T������2ߺ�
X��sRVHF���|%�ojS�W��y-�2�x��i�,��� ����rz���TOk�K��).�{����q]�7�6�ޗ��hl��v�FLu�W>��F+iHg�1���qr��r/�����	s������GH4�Ʀ�+��܎�����N%E���.��t�<��h��\)��Tbb���H�w�B�����x'Qq"�d�k�����,��������G��;]�
p�lA�D�0B����('�h��oW{�^�����U�u[���p�b�M?[�E���Ckܦ�6!!F]X0��ұ�}����k7��:t�y�o̒�/�m�`)z d�ѣ��ś��˂��!������^����q��gA�L\ Ep��v�:g�豲��B�=5���ײ�A�j0�	4�)���WR2~q�����q�*��φ��׋�פ<ː,A;V~�D�W�j�8��Q�+��R牔|�	!��=n��hp�E
��6T�?�'��k�\i��xlJ̟CW�In��k��g@|]�N�oߌ��KĪg��׳�bI��\ɕ	q��|�V�������Vvk08�dhi�Hժ+a27��n<mN���xEK��`a���� �_u�y���|m�O?���4��w�>o��	�f��z���d�&ı*UX�*tb�\���#LN���J����'�X(԰�f���Z5�2��;�8˫W�����:�Y�D�,�?��/��2�Q[a	lc���P�6?�Ě�=���?�Q@$9U���Va�L���nN�^��8�m,�W����4c�$�kJ���ˣ�rn�E�ԯ-��T����
����/W� ��2Q�-��lX
_��V�(ÖD�~d�$�e�k�(r�raB��g�ǬY����[�].�$�Y�_/�AX!�ƅ��s~�}�wBk��G��3Z�&����9x:�䒅�Plh}>[i���516P���ﻡ�Q��:ڟ3�|AS4`0Qr�Ռ��f1�����%SӁH��={e����ȜI�>�������M���)�#�c��"V�{`�lH�Ƒk*M!�M}fj;�Ƹ+��(E�H�5����bw��P�P�p��C�5�۪j3�i��O�V��{�����u,���G�����R���ӧ����b=�-�����+���Q)^*�z	�$
Dڪ�Ľ��U�{ãI|�T(sL�7�R�0�T���4�y�u�wrA��f�i�u�O�RI��d-g�đ�Zk���lBOHl�j�(������YA0$�5�hn�5#�������#����r��v|�0_�sCO�̋�N�OUB������H�D(��I�إ��z잎UR��/N#���:��X�:G��y�S[l�~
������2���k��vHT���<S/����n"�������`�z��RxCˠ�l���M�*��M~��pK1�a�˘m�)�e�qX0��f���(x��]'� y�|�&��4b�8F�!�6�:�w#󲩠�����k�����zQ�eH4��7޻��8�́���7��e����/)Na���!��:��Ԁ���W]�ΐ�|��_��/0s�эS0���n��Y�s��)�����B!����`�Eͯ�b8�l �Kj�2������'�[�r�S)/#���1�s��w�I�L�C.���a�h���X�>7cF�U?#�	�A�]�0��3�g��;^��$T�_�9,�3y#��?�鐕NM��!��2)���%�c��-���%���L1��p���n��^�������6{�͓1Z!�Y7"7��oV�g���,�Q&|�[.9�][��A��� ���Z ��ￂ�*J� �?�T:�$"#'����M|�.4l����Pz+#
SuQ���Jz�Y���� �KIP0��aa�%��:㿆-�,G^�K��Z_#�ս߱������s�l2�e��,�C)�>��Od����ѣ)w.$�G�B �+K��OP�G���A&�7g	�l���A�@#��)H��e��Nw;Ç����@�^*��;l0�Vj�X����Lp)p=VF�94�#\���Γ���A$�S�QfI��|�7%��T4��6��x~���H��1|vg��׿T+�Y�}�����֪�ޢ��k�;����i)�p2�*��Ⱦ%2p�|�A��j��g�%p�]��`ڍȗ_��I�o�U˨,~z��?	�(mQ��J�?��$���N&�S�owN;��,]�h�4S���YDS�o��,��G�e�u=���e����(����| w+l��0Z�)4ĝ9�Z�\��l��� �v�u�R-�$ս�I���N�|�{S��pT�ik8�^���Ie 3��&]��GlCB��3yρ�����vn�8�R&��x�័�� ��[�0��� x˄Y�o�"B�̢�&SG��^�
Fâ�8���+Yh0\/3����{(�G������+���0������G}aV�tHp6$�s�5��\�n!�:��p�,�y�U���Ք��<�h�;Պ�^P����|�ݦ��d���t���5Fʛ!�?��M_V�ۀ6����#����Ӓ��-�>���}@CzЅp>#WR���#\���E�е"�%5���&=Ko��
�}�ͣ^9`qJ�,Q57��3󀥎9w2?陠�k�)�dX��A
eV��+zЛr��čwsEB��5O�r�S�l,/ף��t�3(YD��jZ�a���)��>�Ǟ���\�|�'����̡�j�	H����f��&�,��Cq��/�k~�~��`w
�p�hl���H�]Pa�=t
���[��Nt�\��� <O7_^0�������w�n��	�rh���+F9�u+LJ�� ���>~N�M�Zf�
_|.�/���	���{!1�E�%�o3�&�w!~��o��E��x�#�B>��G	\��B-���]SZeخ�ɴIY�/yg8��+bǧ �3:��w�"�R�K�sŌ�c�&*�4�jo�sd�Z��2��}�vR�[F��)��EL�r�/ᮒm�J� �H#���!b̗�&(O��E �"3=4�9�,�DwV�z+g�����f��=Q޺� ]4�s�����΀,�^_�pR���&�K�SHp�;6���E�Y��lĢg���mi�t�"��-��/�
�X0����/�}8�2�9Ԏ�i���y�����x��}���\�ƮϞݙ�o��s��^K��)ƻ�;��&X�3��%2�@�qYI;����|En�.Nb�T%�z����/"�l:�[P��y���v�����j��|���P#�tO�����Y�m�.S���o5���f u���CX�:XDK�	��q�����S��,�̭<v�kUp^�'k���<4D���ծ�)�aM�_
8���#���P{�V
��f�|�)�����	K+Q@,Jý���G�Ax�rOR����Hg���I��b��,�'�kq�3��������/��/�X$�Z��=pZ {R-�ɡ�]`k���\j���P������$D:�vQU=�P�����0�60}���!5d;�ɪ/��o��x�+�>�W�̅��0���+�n��н_�ꃌ�s"J�'�����=�"X�RW*��S�Њ�$�;�J��䟋�7T�ٹ�#����8������EydV�t���Ҽ���P�L9�	ūj���:[��ʈ�>�{��Y���3�MBӌ:�����)䵣���q]��[�@W�{S�fS��������z��j+1�0��ߠp��M��Ė���>d�����d�S���v�>��ni�� 	"���F'���՚�*4�3!W��KL�d\^���g�\�G��G|ڗ͋LY��6�����,'��uP����D>��މ_mHؐ�o_aI��K�ܶ�$��[��q�GY͔�[E�%ǰ_�F�:]�a���V()�4?������)o�2A�;��Y���)`���:T�h�:ȉ#��G���YL�L>�/���w��݅� ���S�K��e+c�A�d&�I$kV'K콩��1�m�^L����P��6h�;:��Qt�UF#f����s�b����+�J�Ϋ��1�|v�W���GM�|��y|�A���,_'��M��3r#�BFs|ț��%L���2ū��<�O�R�/&<�фB���rh�����´6�( �J/�R�k$���;�-
��Z�!ҙބ	3�����g�����I�1DK��p����O�m������ar���<����G�Z���S:�r��e�7'[�:���9`�#�OF�2Lm�I�
oS��GW�(�ὠxY�)~��X�i�
B)�����z�A-����W���������j���.��_p�*��ֻ�k��W�u�]L�O߶
��~����s�V�mnױ��d�G��S�=�w�֏/�$DmM���:�c(�)�D1�vt��$@v�`��6gK$���̴�a�G��݅~�qq� atV��mz��S�|$�,/r��S��*�t�S���F��0<�㩵z�ْ#Cȍr���<_1���Bٟ�:Nb�|�[y�#~���m�^��U����q����+�2�O�v��:z�O�.��?S׻QC���Ѫӽ|E�aE�p�9J=��S�=Ϊ���@A�01Y�\/�a��;)�n�� �Eۋ���y�L5��M������_u�pq�SJ���҅�Q$���i�g�}���l�enřrA1�ZL�"n~b{ňa����@5�xx(ĕמK?RWĬRӰhy��$q�N!�"���xM(x��g��/v�-m>�g��0	�퉛�h;�1�2�'b믪�ҊY�5XH��Q���Z|��#�d��EL'WU��G�2!A����Y�va�;����J�vW8�����pBL�͜ ��8�	�������&���m�=2��Q�)?l&ބ���t��8�����;0�}dxF���ק�mӷ��Dj(w ��b������;�L�8ys��N1ȹ��e��R�e.��f�^[\��=�hJa45�u�0�U�
�kQu�� �,��w�F7�9)I�z�sA�#F��K��IZ�0��e�qaZe3���Z��%��ٸ��kvP]��� ���5�ds
�l`,g>8P(�"o+/��^,���͵� E�'�Y�NA�.edv+�� ����C��&�0���n�<<��[Ь�ڪ��o�j�ݿ�\&����7�y�\2RA���C�}��v�5�v)�9q��C�����-�)lG$��xD����y2����ӒɇV��w���>Z�}i�=`�|�"ۧ�z؁��\ �Fп�{U��<RKm��B�nsq��NF�R�w�b�K�ѫ�~H���W��#UU}N?܄�?VFZ��VBɸ�!�h��}��S�4�h���N�R�����w�U�+4�4Hq�M7�.����K^��r��T7[�����BL���'b�H�xH��h���Цϓ=��n7�e�w���0���w3bPul��%����x�E85?Z���l��`#�E����������*@.���=W�)ma/>���"�1�w�3Ǔ�0unY������{�eu$�5��z ��x���2|�͓Hꄫ���7w��Jv��L�f��n�C /
4ᇗ��~�Q^%����ZQ���;�5�?�Q���V۸A�뫕��5���v���C���ބr�d���B�sgA��e
���"5�jeBK�H��.*���9��d����$Pǿąv�X�o]B]��X,30>U�!��Y��2J�˻�f��1�;�a�]H7ـuj1(�˩ϭ�	�"7��7��@G��e�$M�՘뽹��5���l�S���%�ȴ'P[�H`^H]5��s����>5X7��� p�V�^D�X�1'�nQ��G=�?�Bk0���jۚ��\��͗n�w�{
n�z�=��#��R���F��T�X�p���w�w���$�b���L�yX�H�nq��TI�&saW%&b�kv�.�2H�ׄr�TP�A�@���J�Ae~7�b^1�.f��k�~H�XwU��Hk]���3�1M�t~�E]K�پ��k����h����fnՍ�[�3Pj��TVV��?�L��s'|�}�+;��70[}#�1��!g>�� �~Q�\H?匩�w��ۉ�4�� �5V���$w*�T�n)6b�̱�>̚��V���en�"�4LB�0b���W��%���i�������:����������B�baW_$���15ZEW˅�:�0Н ���Q�4K�[ƛ�	�Y���;���ǡ�8�2�J;���}X�r�h���Tڍ;̻�ٓ�g��u�'�o��T�>+��2�F9��n�T�����P	��-s�a�(5�
�&�i�	�Xer��5����_@�r'���V��K�f�j������
��y�-�~�:I�u��.�4���Lm��S�6x�ykU�x���3���m��w^�mV��F�6D��9r��:P�>@�Qu�-��WS��F�>1���x�s>�A�����ߟlP��n�(��=���g�DY������������R����]Hj�����I�~T���s�)K�l��(Ǚ���������|6���Sb�H��`����)Q��1�X=�ʽO6���=��n����Ͷ�G�����%٪�&=�>�% {v��L�(O))F>��4�Vж>;#�7���
�	1���g������<����PtQ� a�mnzx�6f�V�<�.�8�[�h�Sv֑�D�7�� ��!��Q3�=��D����x��D�V+ ���ܿ�e0��r���1*��|�O�V���Y�������Zg�)L����Y��Ki�6k8��� 6��]̔�'����R9ub�M�M����'��#.Ȳ������[ݲ}*�{�_�X�����ʿu~��P2y[;�ru>Ȼ��+Q"�QD�l(�B׎* �ՌO��X�>��gW�>LVC���|�1��9�ʳ�6���6"H|'��Vr����
�f�L�IY�y �]���%VgF������S�q�X����`����v�x��8��Y�^9�����k��L>q��~E���x#����  �CqO��T^������<::85y�a�����p�_��y�
z
ҕp��5YMa���J��"1W@�"y��O+(���l�*�@>#�	G�\jp�t|�3r�B�Ǉ��b�Hп����ͥ��%���?��y�[��$ǈ�k��d�f��o���^�"xȦE ���}�Pp� ��̠��ӰE�v�vVH�p�	�f�+�����'�8�$��gy���N��:�
�G�+E7�Ԇ��>2(n����q��{���j[��Z�>N[*������X��*�0T���)�c��HS^| �w��qѢ���FS��l��eK���ը�V�Ԉ�U�y�����.Pk^X!���O5��M
 >�	���:�Pd��#�]Y������aZ�����>��X�T��#k/;��C�I���i�,�9_+a��� �x[G������`���\�J�
1�mp(��a�(G_�j��+]�KԦ�x*��A�G{B ��/l������Lc����ݝ���*�N�O	"(�Jj�c�#��~��C�vJk"2�Gu�P�fXA���N&?��G+�M7����~J�>ؔ�\r}#�����w���F }����7��Ķ��e��s�4��]�����&*���w�H��
��/����D.)KkOs6���x�N�0�"w�˱�N��� �5�-K��/%9���cؤ	�]��/���Q�|A�ˁ�%#Pa����͠9E-�j'���k��e.����x�|}i�v��bs��D���(I�m�⑲��ʷ(��u�Q0���������L��rG�~<0R�Mf�����W����ճ\����m�s\wI��XhZ���LH�.%�S�1Д�#�i͏��NяȄ�>�k�bW�[�\�w MԈܦzkT9Y���C�����ӗ׋��9�tOM��)��7%:��&�Ҷ�J?g�ѩ��ۅ\w���muSt�M	�knj�My�	��(M-_n/�oN��Ȭ]�p�,!�@p����t���aэ�@���+��*2�����G�GV>�eY�!$���)�̈́`.�i������V��(N�L���l��x	(���y�ʉ?q�X�Azeɥ�P�Qߏ83�һ
�\Dꜥll9Y_�n��
Nw�G�QYr͆J��lˎp�ĝٳJX��6E�P#������3r��1Ě��u�k(�l���e@�Th1r�@>��1��_j=�&=!;�Qo�=C��D��@F��6��{���@�3g��sW�d�$����m޻Y���꫈�P�-+���8���kWa���cl��@w�a�m�۽��8	�Nڊ0���*�
}�Wv�t`��ZR����hx�����n���[�(/�'2mU�	دa��.�!�V$ui$�`}|�>��ano�h���0?*���oN��UWK��M,����d}HI�^X�Pd�>�;~C:^RJ��nפ?��;��g
Ġ�=�db�v^���Xg��P`�'Bш����2��)hU�0����r�A��L�+'24�����h�s��}��5�iP;P�a���&��n�1�R��lEm#�g�+� �%�M]%��Y#��Y��HȆ*YF:\��C�v�R�c�}���QА��ut�ty����wKy���]$�U��z��P�gdR�9{r��	e�Ԧ�!��D��%I�SŶ���˩x5� �6�z/�G5
��ymEۺ},��u������)�O�YKct�5��<�|0=��-%s�B��
���G�Ȝ�q��d�_�w&T�V��ڛJY���l����6��m�B���+��!"֩�w��d�6��q��O��ޑ�KN򮖀���xkvV���c��C�2*�����Z���	��(�]�Σ*/e�u��y�Z�� 9�`V+9� �����(.En�V�> �� �Q=Ͷڃ��_�D���UB&6�n)��䤪���lY2����B^���}�3D��ZdSs�8U�Ћ������'��L�8�p�f2�R%=�$�	(���C��ܡ*�fƔ���S����z�k�I#�;���IӷBA%�oM����L�1�r3��>E�m�7��G-���.�� ��6Hdx5ke�d��s�b@g���T�n���|]�:�� ����S)�>_2m!`8@Fc*�EAGO9������kBJ�Fk�r�Mt=V�L5�E��.��+�A �A�m��k5�17��!������W��`���l�@𓂺�\�%��j;���w鞺`r�o��ꑤ�Ce(���m%����-��m5���9�c�[H9�&wɵ�4=�wn�d�l�팰��Vq��B�A�v�O�!r4 ��<Y��e5k�K6H���U��'h���@ �6����%�w��cBZ\}���<��(���<�-�Ey_M�
\ق�K��H+�}A@]�U����}��+LsUKf0.	g���)3����q粠�7
��A��og��#�h����{C��Ԭ���|"�h��I"z�v�.���Y� j�����۟3�?R�+� Z�h*��=�B�y�F:��Z����*@�����!~|4+��)�|�2u1i9ݿN1I8���%�}�L��m��S���0F�?:��;%�a!v� Gteʩ����7Tc$����,cR����q�WdI��w�?�{���A����f�8eKP4�����
�b��nA����֑ebp�v��D��9BT��J���e��D&�Ԕ5��{UG-ߙ��>-������G�ѐ�w�
P�w�j��W�V�>�$�� ���L>"Uqb�}qz^�}y3�R�^�੟�L���my�h�e�H����cDk�A���X���N�胜��tv��_ ��kb?�*፞{� f��J7�z��|F�D�b�]I.�����0� A��,$Eh��e�Ә����Խ�!��w2/3(LY#� Г-�@o���N�@UvP�N�M��p��@��>̓�M9[߇�[������7�u'�p4����]�$B�SXb�}�0�v����h��ħ xo���}�$Q�R�%#��m/�L�"G�p\�w��W�s�ʎ�w�U��d�-����|�L��9v��ziA�v���e��Gj}`�AB�S���T��p.���p ��) �.*��mt���� E��cҨr�M;ȴEe�T�n���-����ٛ��gXن#�B�
ǿ�(�q���#�'��RՀ��r����)ݎz<���Fb_�^�t�ٍ?�y��#��^tܷZ԰��[��.I����^mcyu?�Y
�x/�L�!U�﹧�tו.�/�6)8�ϻpŃ\#��D�ް��x�γr�9i�
��07讍蒐tYx��ŔE7dB�V��@�x��5�$0>�9�(�Bi����焉Q�����(���_�,���*�Ů[TA+������kɀ�/x�)
�O}�E6i�U���	��H�쬜Bf���eU�)�����H����� ͤ�=��ix??�Y�_砺��q�������0�1�t��PZ�]��V�x|ʋ�т�!�)h�����\����o�SvgX$���zN��E|����c�.�ݷW�i�2�Aú�}o\�s���1�ꇷ�\i��V�j�70�ɪMY�\��&d��^���eԪ=��b�:��4�-���>�	�aUG^&u�������4}qf�ny����:�C�h����﹠��^�^H�v;G:Ě�IeT�� .'����e���	p[ �ޘ�0?���>`^�0��氡@0'f��C�����9����<�Z5����ƏE�ޟ{l,P�P�<ys_q� &�ץtp�Ц��:����n�i�q�n+�i��}1�7���)ڞ�G�� �"�j�T�4�F�?{���s	��g���PF8$�z����o-O$	}VX�O���v�o�u$J��7�gYi�n��RE��H�3([�Dˆ����A��slDzO�H�^���`���"��|"�п��\ ���D�?�'8���i��f��s�IN���]�>a�;�lkP$�@� �?�]�W�2-;�|�Ƈ����T/��Uq�p�!
�Z�����$��^�cVitW���5Le�4C*h~Uœh�B�YX��ɝzS|GG��u����+s���ͥ1�a��16�s���?�\_��Ҥ*őB���.�&r�Mԃ�[{:���D��iK�RCp/%G�A*د�����qɿ~	:�ﻒ���*{�)V#ͩ�r��=�!_����U�,i�D������^�
�1��%e������I�����tkHTGӵ�غĮ�h�������+2�����:�`Nl�Ǡ���Y/^�f*˴v��f��k�b��t&���g_���,j]�l��$�z	^3Q�w(�V�.��/(�:}C�D���S)Ь����8�uX�Q��a�V/J���|�� �4岦�z��P�Z�%ݕA,�����+V+l��Nو�hg�ǜ u:i�cK��l���0�A��H����Q-�@oR&؏~k��f��������.�FW��҈�X�5���`�qA�h<�B���̕�z�)�T�@v�<����yWj�o�����z滶���0�j�xz&
���Xٍ��P��h�_��qBv�P�KZ��k,MP�֜T����@G�K�_�����3/Z�r	��/��i��P�Z%�W�`�|6�As��@��a���,�O�ŐK\��o�OE�����*�Y�'�imYn��=ʽ�[.��"Ο�`l��G�^��ӿ(��W�>�#ф���si�Z�o���76�;����ŪNZG*�5Y��c+�#��s���Y;c�7'F���"�.;���VO���tN�R7l��k�-�9��A̓g$c�Յ�ɾ~����=A����Us|Y�gѷ��]����(��c 6��~�צ(�r.�Y���$A�N��+�^5�������d��I+��A�����Y.�	��o	�8���;{٥+\���&���G�s��Wa�������gasu��B�?�]����Cɹ������.��P>L oA�	�${���	�
�1���f#&|���&�I��O����پ �#�J(�=+�,a̝o��,B(\�� 2xx�m'�$��3R�Ȏ�z�*iu�������uk�p�W�	��"����3MOJ���p�9��^X�����<���c{��eM���>���g�α���x1�Qy�)��9�U�['RJ���7{r���y�IY۪V������N�`\�}4?�U� &dD� ���š�5�Đ�����[0��^�K��@��� �]�l(�W��cD�	����Mʄ���l���b-dS{f�5��� W��[JE�׭q%R��,�m������[��͏�L�&ޢ��~�:<�I�;h��(�Œ��»���<��l��'�U1�R--p����:'��rJ���Ӫ4Z𱩝��SY�7ͫ�׿�D �н
f�}'\�ĥؽ���I�p�*vL�>
=�L����r���?$�"-GD}
Z$Z�EPoS2ʱ������Ӏ��Պ��){n�zĖ\,w����O�d�U��R/6n�@���+�O^�y:�[�@��i��"0Y�����$W��n6�RR��P��&Cze#��Wk�8�����O��L����kJ	�-�a"���T�B��.�A��Б+<�pJp�8|a�q_t5ƫ	��fF�͏�|��w�ס�Cr��j-j}"i���<g���@�0�ራ�$��t	��;4�{�ph���xo�=�fC(�v+S�M*��0tDdL���T�.���4V\��lF9�m��h�7��$p[�{�z��9'��L�*��1Ujl�CtN5�rt��!�?T-�����_{�x���'Z�wy���i��!�S���V�Q�XU��*�Z��4�n��d�hi�H��0anp�Q@�2t�aq��d� D����8[��� �P"�3q}�~�ދ����H?J�e�	�hp�u}�
�`��{u��Ș$c*Ԕz�����Q�~�qz5�v8�@������R��e;� m����Z�B�P$��sN�"����uq����ϲC���>e�${�:k��ҏ� b3<Y���xq�H�Ƞ���e�Ţ0zəK�i:U~�P�C6��aK�>Pp�H�[̪4A[��aD�+�����J�tE\/y��r=Ko��Mx��,ϵ�e�3'�e�( tSx|n��z�1�>G�j�]�|�Q�+�+\d��j+u�m:�R2���w�rc,�f���6�@�R���.���ބ�ڔ,Z����AC�����k������D�u��C��Y#��lgN��}Q2�� i���<z4�K��˙a����,�ӱ��C�z��������u-4K�r��NXh�w�Z��"�M-q�Y$��m�{ڜ���	T yGǬ4�`��ym���]kEt�D���f��}�v��Zә*25i��T��.{�v� K'TLG�>�/vO�m*��?�ť �"����1�����}���m�K̄&�%�6|��q^
#����4翝�N�>#auJ���c��e6�s<��t�iΤ��e �@�ET)6��`�9�%ׇ��$%��]C�@�X�;���R�wǈ�?΢���Gߔ����/�h\l�/�+XS8r������a��j��<9咨�(!;�H��N7�!j-r��X�K"�� �T�ؠ��3R��f������Id�Ѽ^/b���^I2�u�]#�rs���g^b'�$���>g6��E�,�W��!�S_��h���ND��˵���DY{e�F��	�����_(tP���(i嗪�B-�w�±vM�^S�@|�� k�>�`�:=��c�8x/6ju�x�4���/��VF�A�w���F�L.���uB�C� ��ĥ�_�d~,Գò�������N�,��޸!Y�X,�u~��TX�D�4��t��Xp��	������;����p��9�["�B�<9󂤺z�3	c�Jr-U���t�����g�E:
�h�\����O�S�e��;>'�Q�_�5�J���"��.� �m���U�u��y����ٖ�N<��f[f4�H��,��4ئ�}��4iҰEikP����g�['������Z�Rp��"�{�K`�c�'h�s��n�u�F��L
�,V��M�m�}�L�o����:�|W_�_�j/�V��g�u�|��L�'��&������p��ŧ�P�샹�t��e�v�ݞ&����{���o��'� T�W4>F��3��W�x�I�å�"V���TE�U2f� sj�L���k���:d~�3v3T�oB� ��-ݑ	�m.>�� ����]�IK,_���U=���P�VEC�X����
xbՇ���? �V�m��|P�h���jh�4��V\.;$ Se.I�Q��i5Tz�m��[m���򸫗�;ب�x6Ŧ���+��8�bx�h�I�95W�&����&(@�a3ojf��G��L�TPK��jI����_�d��o=#��"oR�Q��,�C��Z�Bt(և��6T"���|Tv�,�F�h�7� I�G��c\��AΏf�����82$U�|j@:���B�x�[��DN��ӴO�m�0		�!�	lە�=���׽T:\�u�Ü��|d�WL�Ƈ���P�z)��ǐ�D��c4�p��w�-�GLw�%�i��k�0R.b�����E���~ۚ��m��feds��P�o�4foԈ��K3���u�_�@Vɾ���x�����t2�FZb�����5m.���K�m2�xL|-W���� �w�ދ�0e�	�s�I| 	�s[m�}X�&�^�pd}�W��������0�Ӈ������9��a訽�[&����0�=V��ι��V	ܴ	��$��:?'��с���_ǯ�Ѡ�=��f�+��R�.���@&`D;�����d�ԟ]L[.� �I���j��.����>p�$�u7E�$�Ƚ��U�D���<!���tVl�����]o�j�����o尛'�U%ğ1@X�66p�����2�e2*�7WDm+4���<�@�j;e�H�#�D��6HUן.b�[�lPH#>>qK�杨]D�Z;~����-(�]�O��;��S%�i�S��'U���=W�	�o�q��uU��`�p����g3:��'Q���z��W]�6�D����xjt��y�;�F���V���`n��
�5�y�|f����л5ކ��G��h���f*�R��廻�Zw���d,g���NAH����^�[*�n��ա2��''�>&2�0W�)jw��BV|�4�+�T�����w�0G��.�وF���`v�֛o6�����x� �m�� �>���w�XJ �nq��r�?z��*�<��'+���j50�W�Hg�l�����9Y *�Q���E���Ѹ��C+��T��g]1_u7&�v���7�Ǆ-�с��nfuxmX��c��g$�GA����f��-� 2� ��r;8�Т��	ɗ��n6~g�݌"���5��,��o���� ��������a�Ko�cjԐ����n��(c%�����a����8��ͪ8�&�<��'6Y.þF"�I@�{e�_E?�i���?.��o'a�ŏw�i��}m�P۷ꕛ���H�v�F �9T����E�GU`R�	�+i��A��OC�y��� �
,#Y[��Ic��\��%�L���<: [ ��e'v�����}z���03���T�r�L�R��������'Oi�"W��#5I%�Id�4��$EA�k�~:&�3m���%��)��/yO��KZb���ik�`��X�,���I����F{�篳��;#Q���*�@K3�����Z]H{��UE$�����_��pfGg�<,z0�}x/i0�9̻��I��O�A�c��Q#Xw����<�1�#F"q|i���)�2 W��yŋ�8��ɔ	�NI�`�� �(	���YP�WĲ�d<�c*jg]��`=;U�8�xG7`t�IY�5ǖx\ſ{�����Й�d����}��l�GG"�A7W�d�.�%��G���p��hiA��ι@��^��>� ��MW�����n�T��'[yۭ>�� �cH2:
���`f:D����woR�!���=�"��)%}�ԭ��*Ю�嶀��gH��a�"�X�<F�x1���/6=_�x16�ʍ�H�+� ��%BL��w�1�C�j�����޸�$��?~C�_�o?�[��S�a�2�&4BG�d����m������`�N�F&��--��<���G{q���Oy�TU�Iy�%kx;m��zbL�'��V2M��� 9�<�������%� '� 2�@ q� �L��R\�$~)�4Q��k������y��0:�CIfE�噋h�T�?� �-tjf��yG����ӝ
U���y�Sc�8qk9�{ĎCv.]��0-��g�Uf��&j`�����H?����:`�����b]�u�b���K	[�P$���?u�,�������YZ	��Ѥק��nG��5C�_��r/l�,ǙPD��$&"j��Jl��~���_�3 Ժ���P}+�#�5�u��eص"3�,(+�頄�-��\�㏷{<�d���Z#�IERۏ��$x~����E���Am�4�:$����`o/ڥ�K���D]ǚ��KܫXþ�e�w�T�*�H���c�/���1�7�;Z�$;����E8-���[��s�4�а#�ep�N�l��^/
�m�[,1Q��r�ZPRH*U�Ξ$�&�J��A ���m]n��y�����>}YC���Qű�����J-1@�~gN�*�N�:O��?:zi����gPp�Hi`�	��bm�M����V� ]��^Q���A��E|z#m�G���B�U���n3\�ʻ��=���T�Y<�9�B�m�H#c؋��$?/�X�n{�p���1���oYn$
����?]�F���}.,'������*x�>^�e�3�UF<tWR%��!�Y�-�L废�0�(�[1ZN�$Y������;>�0���X�n�բ
A�Z\w��&a�S�j%tr�o(*��U���M��t]���)�i�Z�+ԃ <6d5t�	����C@}�Z���Myb�s�b�v�.,�E����=8 ������1[�({��գ�r9o��k��0B�NF/������ߠ��B�m$$�jff��
�f�kChZ��gקfS��n�$�xc����tR.%�z���~��ɒK)s�7QF6t�3K���Z؀w==�9�$������M�،����/"�N���v���s~@�J �<�u����fk[���Z�$=�Hg��5�V:`�!s��ë�P
 ݦ��SJn'��s�p���~�[����{�KqT�7��~K-^�`���S���8b�9�d^�L	yn^�>�f�ʴ��>��@��/vN;87��SE~/���88�Q�Q^�uOD't̴P0&*�{nSZI8�&��|2�(|0A�����
�ܳ�Z��s~��p��E�W9��z�ŉ�OPv�3�*���aqN�Xʏ�RL 6"w���;�8�}<��ΘHc����?�h?B�ht�����}����Z���+��x$�N}Ɯ���1�#���.����"/m������By��Wm}!���\]��1�F6�x��hG)���_���J}6�j�w����Ts�mf^(�ظ���v���o �>�l�wd��{������xh66�_y[�f)��in��X!%�4wE���z��\�1`R'��u$�cY4�Ћ_k�����0�d�����3��K���(Ԫ�m(�z;���8����1c&����~SV.���Fk��O��w��P��amC�f�=I�&Ű���I��l��4�q5j�ݟ@���s�G��ݍ� AG)ll��>1�$4�@?�����oPi��`�X���M�G�d��+/�h�2�����RK0��9������_�Ybf�ŴN�AT�9/�����<�����9��9� Ӕxϙ���}�S�9�N�r<���,����]�W�0k��|��Y�֪!뽑$h �K�CyS~��-�$�w��1�j B����[�'u2g.mZ.g��L�뙢FsA�h��?�t�z�F�D�+J�n��+=�K���C�;�6����!_vGC
u�Z�3�e: n��p�8�G�SJ�o�m�8�l���>�$K��1�I�-������v>@�!��k��DШJ�����D�ɧ6�\'�R���o�!�����T�E�m�ɉ�eU�x��Z|(�xq�-�v=\2�|��:��v �k����t�`��Z-=��Me��b��T�R�{2q��&!�B뼦;,� =��ү�q���=���Gw;���FQ*z�%顾�myƽ ����е�y��>��b�����ɾ5��Ay�0^����#c��?���WK��ڇ��(Nu�r�'�0ES;�$y��z�۞mkL������'��8��}q�����f���:u����-�@z�4ǖ�ۤ�>E��Q�Y�0%����৺'�H���|{��7c�J���,,��%�M?
�8�\��~��l�3{�	}�sx����S�����esH+�ܭ��vL��f�)��^=���u���W`�s#]�7*"ףɀ$y�Ue%<�j3��w��M��,����E��*1qx�%_�9:v2�n�v{\�Ԫg�u8�ug6�Vt��n�͊�h�KC�Wb%�m�ԉꤣ={%����#G+��P��3�o�lI&��ʏ8�z�Q�����@u��
'�ʄ,��6R�:���|4vZ֎���
��s��l�X�]'��"~��N�P���-�#��q�P�;)��|�8�2Da�y_�V/��{Gv�%/qS���$Z�J$a�^�"�:�>� } Ď��hK���_w�D�_���3`q97�+X�j��j�V�hv�d�1�+�ԛ�C �)�E'���C�/�W��а��W�_��ԏу�������a����+��m��g�GDΉ�.O��-���ل?���9��=!Z�����SQ����#�:KЇ���㖨��<�-�k��ŶO$������	m�yuH؞Kʍ���/gI�]���dy�˽>m�ڧ`������t��~�[h����缦�4��HP���h���d{���{�s�c1o>�l7����0%�)U�Y�����`����a�w%\��>�3-c�z� �oJ�����$(��se�S���s�<�ڠ}S�%�l�q�T�C��rU@*5˼Z���
�����QK�7��"M��F�D	U�f��,�i��>HCF?*mKq��!��^6��塱���I-���p��;0�ղ�~ȉ%�'��B�ڽ�]dD4��^P�-ݭ��� ����U���[z���"�-i4��+��l\��0i*�gG2HI�5Z"�7j�����$�c!~8�kzXO�~8��8dU�(�NH���)�z����h�<�z��+D�ҧ����Dڝ�.g��pU,�n�^�l���֪M����b�R�͹5�(�����۲P��	f���7HB�j��3�A�[�1��k�<{��ؘ����	�s�Z����F�M8BO��S#��Oq�nrXd}�G�K�cx~�B	��k��.e�Bl@��y����}kҦk �Si����ƽ����!�Z�B��i���UK�[�`��àq��c\�A��sI�"N��㰣�Ŏ�������]X{�Sk��/paa�{``�FW�0�m��c8��j�	_��R��>+^��j鮅4Gi|@�z�%sQ�`������O�FUf~)�/���ɔ!��d��	8j�=����<��O�mO%'�M��^���G(਍p�Ard,�4��S�����x�C��2�X'�o����3}d���jA�3�4�Z4!`����װaiM�Z˕���-�x� 	�X0��F;B9���G�sY{k�8�<���I-W�r-p�0	��@�wtX��9m�TYb�6ވ���!�x����(I"��Y+{Ui&!�b>�]+3~���օ[p-��&���.���w������o5ifk�c����$;�Et���%���oS�Q��<��DzP���_���U�8�<�W��1��V0k��[��8��WwX�b��՚hG�E@��l�xÌ��RF�� ��u�a�z�oʹ�g���t����{u�2�).�Α�4��>��B&�6��WЖkUT�2�-��fB�l��A���,ۉ`:U��n*��u���� ���ܴ����
�n8�
qY���˝���*���e�Ԭ��3	c�
n���P4�@�9-�m�h#
\9(����L�F��n�n��6��ۖ5�w���-x�tS�(C͌=���+�Q�����w��Z��B&�� �7���� ���f�J�0/��"5'+��y���r� ������v�g��Ǳ9��ҕ�jT!ܵ�&�4�.)�Vk���;{f����څQ���� ��#ɲ�Uo�x@��%��ȣ'��LE�cR�@����N��b��RBЋ;j��Aq��p�ϨW�0K�iñ��Ԕ��pѡ��gQZ��#�ٞ�4Hn�fZ������Ԫ1Wz�{�y Eא���YPzO�NgH�����V~���t�����`�+'�i��\,�}Qߔ{LG���!���`Sd> ���ؼ�	�"��$�а�a}��m�4z����vk��(7�TK�s0���8��w��vR�� <��X�(5�Q>+�]�
W2>u1�=!���b�j���L$_�~3�m�1���Qa)��Gі[��S^*��=�5��8$�T6z�q���#�dG�d�jnr�Z%��bblvg��c�M�ay��{r�1��jO��a��kd�,@ņ��IS������V���ӹ� �
wQ������D�M�U�"$���bEX�f��?���-G�\�\P�����c?�Z�I�%���m�N՟��|� �H�Զt{�4ME)s#K��. �b��Gb�y �ߖ�Wv^�Y1�Q�<Wp�^���C�t�uxX��3��U7>yA�6�����W����y�y���!I�Q%K�ە��=r���!ٗ�Qb���{�o�C�]�[wz[tp �]�_��7I���yʫ��d�D�"m�m��)yqxk�k��6�� ���8&�!��'N�G(R�({O�Q�_�>Oɨ]��Ju�X/�̂�Ұ�'���	פ�mp�3.��z��R1��f"hWtC�W��Jg�en
�=���E�j?��٘��S�pp���9�Bi��0���>G�Y�
x��˄䫕I[e��������T���b��A���-�x�����8��nD�>�� U�O�UEejq�G�Vbv�v�	��v�R�X��� �`g6B�S>�"c��v��BދuVF��f��R��%����H����T?�^��L�BU<�/��������R�p�Z����-���ha�ǖ 9��:�p�Nw}�dk��aݥA&���`��(�����g�*��ë̂�I��j���(����_.Q� �9���E�u�F񎥼l���<`��cZD�\��m��O��.5+GӼ���)E�:;3��b%�O�Lo�d���i{��bn��C#P��V�Na��R'����7�q��1p�3їq/w��������L�-��a�J��m���c*��Ӯ�9�X�C�C�P��_�`Y�����	K���ȱ�Nӕ����=��+S��G�a��=Ǘ�(�o~�y�ey����~������E��>���"�eU�"����v�I�%&�erH�D� ��^�AB4�W�u�G�~M�G���g<��ēY�LQ��`��f�,Ƃ�T��/�U��Du3Xo� +,g��Y��sY)lLN'�r�3u�y���z&܆Όyր�Įu�[h�%[S�՝z�����EƏ��� ���0�u`�)V��ᙵ�r�GS�cm5W��̂��Aԧ�����(��`�Kg��/�v+E�"Q���4A�x������V�d�I�!i!l�1&�`�@��Y��B�ʐc�p�TE�P[������l�s�F⚸bq��&cd|��|�?���%����`����:"bnU
�������˸7Ë��b�_��+��|��H��osso�"�:[���j\�ճp�qv��gA��n6]AЫ�£�D\��jE��f��g�b~o+�B��2f�>�1%6f�|�QW~�p8ٕ�$�o
|>9�M�@&p#$=��ܬ����{��˚XE��� Ƕ@	+�v��l$�����/��������x�2�Ɇ�����C�-ʜw�׆�\�n�-�-w��j��eɨ|�Տ��Om��K�<%<c����������*hۣ_ݽ�1�j 8�%^"H�N"D�ih{<�A���lj/�[���=v>��Ğ={����%ӊ�V���Q���fX��9�k��/S�b�9����{9�fdc��e���
\zaȨ4M��?+�5Z�V�(r��T$~I'�� Ŧ.�_k)��B��Go�r��m�*�#Ab|�o�6��|�sq�^<2&�RY�_K8���r�^�s��	Z[�K9nǦQ���$c�iE�z[����44θJͭ�ОrwYuh|���z�g-Z챜�hZz�ӵ���6Tdw4��r�Q�X�	j��F^�p�GTZݡZ���ȆT[N/�?DeFɿ��I����#Ǟ��"D��n� ��[�����1Q�eudJ >���06�1��M�덢8�fFF�{��XaeyW�8f7O�W�M�鳘�B�@xφ��>T^ ?W�чŦ��;�L��&]�7�5�������l
[;���X���]z�*�>��3P5p����F��O�:�eS
5������p�U:y��¡@+�U���Qz&�,-��}��[�e[-��ϊ��4ў�`�|:|O�m�6~1{�۳���mԴ�@6ozvp;��[�}�Bi>�3od{�[t�"�K��e�6ֶ�����"u3<�R,7��oe���7�R_l�E����!���A����v��!�ޙ����}��`R�r�=2��-�z��&�S��^����U2r�7��׋�����4�g�H?;۰��W�վޓ�t���mi�C\�x��VG��p9�㮷~;@nDYh_��s80���:��/KX=#-i?�u�Rup�|��D<�T5��8T޹��hѥ��ӦDm57�m{Mn�V��s!&}ĩvT~�a��/P��,qs!=����`�����������׫K�zۮ�U��F|?(=�	�s��#�g/$FA@�ۓ[�\g5��j>�I���ű7yN����򲏂+�P��(l�A#�Sà��������?�X�^n6u����
^���������k�:�D�>��R�Uz*[{�m ���I7��e�rU�QV_����+� B�ϊރ�)�КP�'Jr@�5��^PV�J]22+�;�gS��%�	*��J�(~>�2�kB��'�ῡ��'�����Ѫ]��fY�^@!�b�ǊB����L7�ҿ��ۢ\�������~�X�Iy,�����章FAs�N��E>�W�hN�{ʻ�,}�]I�{��j��)k�]�n�q뇂�0��O?�Ñ��)��A�l��Wr&(֥�� ����q��׿������F��M�AO�	~���f�
�e�2X��~��P\g9lu���hr?�ٰW�D�I�~],(\�`q�µ�S,^�u��y˥�g���i2
��V�$L
\�0�\#�*m�y�^!�:���z�
��yêF��6���@�����jt!G��R:�|�!Ӥ�;�_�n�O=`/0�����({���o��F�Z4��XQ�]��&P�_���d�^��S�s&x�w.Q+W��l�\v����5������q����^�9`�}���+,D-:���
��T��*FKĲ4]VB�^$�tp;�B�N�Y�-˟-=c�Q���G�����AA���`�|A�/�a�B
���}�pG{ӎ�e�!�JQd� FqC�b�Fs���T�x�IT�F��k+֧,��o+`u�CxR�f�@ۛ3o�n!p=�{A9o�!T�����O'N�*��TB>jϣ�r2w���EΚ?J�B\27+9|:k7��q�t8w�i5|&��znn�!�Xˬ�>BA�\�� n(�[���[��{H���5��w~����hI.��Do��R�^�� j`(F�3��H5���Lͺ�#H�A� *��_��c4�N\��a#j�����\�)������ Mmp�����`>�z�Qd�i��w��AG��Y����e=4e�~�O�]�4i�$ň=gc��<�N2��0"F#�7�����:RDͼG����`��ժ�C�H�ҡ,�ڂ�����E�Wά!�YHV��8�����xJ��Ӯ�v�gӣ�-�P��U�p��C�=E�*�ۨ�҇�e�t���fE��+�ʦC`�\e|kJ���r�j�H	aUj*�Ö$�|�f�f+Y�^h\ .��|m�'���}<��]Ud�L"�$2��$�����.﹤��A�x�t,�?k������K.��0�0ޘ�P;lg*�t��4�~uUW���>�%O8?�.)]�w֔{�}9e�Z���}�}�^ĝ���<⢡ܭ���c� 55��=������5u}��ڵ��=i!�G��p�<c�sb�.��fb2��P��0�� �^y���C7�.�/GS3�0�^-_Y�;�2��s�q��1@p�h7@�����|����v��j���n����-�-M�6�H���J@s�Ext�m�s`#]�Wm}��9`b]/�븚��*�6�P�����q�Ga��a5�Ǜ�2�F��R�s�:�9[�!;I#�8���u{R��8;��"!�7��I�7�����Y:�f�I� v�QtV�N��r`�|zs8S>=��Y�UI،����}��� n���~�5�;=W5?�Cr�OY
��>�*OsX��b$�:)�&�p�۴���&�kd�	�����w���'��څ��M��y��\��S U(U̙�X�ৠp�]��><�lʊ�7���r7�E�۹��T#����7�^�\��6�'
JS�QX�Ϫ5�PG�YpAF�G�}��ٕ#�� ���J�AN�Sj��!����d��Y�f��+��[o����
NJj�a�^�I�{��{tF7�@ۯ"�nDLo����Qq4�It�LJ5�r��&��wǚؖv�t�oM�0�i^������C�a1�CS�HM���)�S~w|UJ� T#��B�5�����z+ _�M�Ѐ�4yw���%[�S�*�
��lHߌ�I���=��Q�R�vcކ
mY�GY���l6DQ6�⿠u9���se���&	�U�2�ܼ1,y)�/��V�a�lQ��ݥ��r_�>쵰s:�G�`�(�q�8cFWpp�9��WI�q�� �5��̼�D����ӿR�L��Z7PYd�����|:�������3��P�{�%+d�JQkjI����j;��ܙ�9�(�G�4����@�o�����l,���`�1?��N�kW�ReS���΁$o�`É���O�����X�����/�_��W
���4�^��a[�<���gA|4�;f�%�N�;T/�����#0ힴ�@��J,�oxFO�Qf(�����c���6�8Qs +lW�[�ܙ�~|��kǼ��e��/�q.\Gp8�
��&&3\Ư�� �׉����c?kHN����+yIO=�!��)~���6�K)�ъf��6��/�(�d���ET4��s���UI0���m��p��1�c\����2�\D�r	wg�����U��Q��:}�t�/��p�R�8�0��U����8ܐP]�b�"��� �l�e��W��r�1jyY�*��M�d_'\B�GJ��ٵ�-����Hµ�m�p��3\LɗQ>����E�e/�o�,�m�ܭ �)�u���Ƿ���Е�5�G���ܢ�Pβ�\ts�=3�=e1�#����*�
X`p��kە���Dr*�PSŀJ���Z�����l���wb�/��ma�{Qiͯ���&���ywt��iO��5}&n"�1k�}ڱ]U�m%��X;o�o�x�F.��T�[�Ӹ��j��4Q���{�j����kǘ�����!�ޞ�rãI,�X��J��)����7�.;´�e���܈����D�Y�b]O��	lt�(���B�?�p��Ok
��8�ib���RH���,l�����Y�H�y�m2F������U� F+P�B��_��5��_A((����Z_r�i��C�k�b��.�Gn���������A�+=4�+���¥�A�pXF�'F��Q�cjF(���%�N����f��K����\�5	֧K��|��s'�L,
pA��fF����1
��@�V�)�2*/N��M6������n����c�XΕ!ظ�(����w9CХ�Y.�Џ�3���xm2����s�;�^�����Э��X��ދ����Z���f�=�� d$���P�xDضē`*Ǳ7��l�.�ۤ�bo��9(�̸l钺9��>OB�h̟����e1^O��	�>qiԤ��͉���1�YhUV
�S�j�״Ѕ�s�է�ˬ�O;ֺM�9[6LW*���� v*PRW~� B��L��EJ���P�S,r�l������T����KBUl8��w/�^�����Z�M�8�r��R�
&~c���
����z�aU�8�ҝە��-��E�'����^�&�ye#�xWt��܏�,�U����Oc��� �d����!�J�
(���i�F�0�F3�(��t��i���,��)"��R�D��M�<�����}8��[��:^a���3��gNO��]@ʘ��*-`�2봣{r�yt��49����PX&y%�y����-�ƍ�5�A�J���:��3܉\eD$8 ��[_=��c����I�^h�lds�b��)r� ����4=\+EĎ�,}����1��ź"�B8�UH���/�}�����1�5K��e��-����R{ `�m�P��б�E"��÷x'���)�u���S;W�4���-(�>�aHw��H
H0�C���Q�2M	lݳ!�<�t7��C��2��j6��G��)>�N�킗�;�}�<B;kSׯ\c� $s�#��*
�G"�1�Fj�������r^e��A�C_���%���̓&5��ہCod�OG��>"4^��9�I�)��\t��~d�E���$$xY�X�b�&pC�>��k"����R�L�\S�#�^!�E3W���-��q��F�/<�W���1��/[�6��^:.�O6Ϯ�xP�q�rB�5U|�Yz�S�;�%u��pօB�5�H^�:y�t�a�c��_�R�xN�@����ܬ��}�$��o�p��y��,�:�
�������Ty�@?�|��ܹ�❀'ƅU����<&���lg&5�G�9�F�x��SY�8r�r��hQ)��y�Iݏ7������P��+���e�"�X+>f&[����= nv���ņJ����م���V� �$_j+�n�X>��`.5�@��t�_e��8[ ��j�=�\xb�ޜ#�����.4�U���QV8V��|�o��wڙm�T�h���7�**��E�l�0K����Tz� SVD6�M� cit,u��O:�^�$���1����8�}+I$�z>E3t|j5��D^�ͼ2
���'ݖ��U�M��ۅ�U�W/��!��0�S��>�a�����\@I����my�Ν �O)Z��*�o�x�L�I����6�0�	���KZ���-^qg/�1~��H>;��8��3)8�2Ӳ"����$�<P���DЇ `s���W`�{� �9���$$����n�ޤؒ㌾�f	E�;��Ԕ�e��#�֫.s����;j�GJ�ʿ�`����.�l�6k+��/r�N�����pV��=Hqh�$n���kaI!�����r�а���܇�����s+7��2rj���,�
kx�t��ӭ�+��h#"�_|�iw-X+���V+�3#�ǋ#�7Bm/����^�w�R�Ϫ����S��r�����@���n�����TP4����H-���BoLǙ�˴r���� �b�`M%[�D���d�SkIb �S�؊aU�:<«�����ͨj���4eG[M�h�-��>K�/>�Xi��f�c�� t�)�J�E���T�$2��8��n%�+��Z��I%��Y�j����BZ�7mV���`�h�M�`���ܸ��'���5Y�|kpk�`�V�E�r���ɞ߲>�҂H�w�?轲���� ��@��޳-��S���+!Ϡ��-�Μ��^�b�:j����.��X�Q��(�!�1��tL�RTJ[�9��o��.T��Z��6k"�f��.
4G�}�O���,�;�w���W�m�L�&�H���&{5�M/�4O22G���K��l��ɅHOf�ݍ� ΁�x�>S����>��d2T���� ��)���j/���q+��.���8�"GL��ܑ?Ws�Ѩ�vh!vEr+�YĎ�sMg]���̸|k�X5E�51|���}���E��|���ζ�U��tU���rM�M���/D�#
S�+����X�amE�Fb�x�������O\�	�:5��*7A<�pHy���Yu��XvU���>jq����͖v��q?�6Tᮐi
�N�Wӊ0�\��'Ft|vH��j�]�ţu6� +�66g�mB��6i9%
)�\��ކq!�d�u�Q��f]�E�z��T$�WWj7�5�8������WV���M����GR���v�����/#ӂ�KYA�g�'��O�&ģ�2�q!�����48~����:ki��
�$��\?���g�::$v|3o&�u��-��1�� �����5h�Y��[����^�+��+���^��������r�UM$��I�p5Ʒ�y���`�(9�TT4�G&�Sț���:Q��E+�����?�i ���/�v�.k����d�/�R��9|��u��n����k�&T5�A97�z��6
�DO�2�)֑�Wk':�e�|7�)���is=�g��%�x�".<V���}r:��~��@�P�|�]v��dj�as	L����}=B;A?��b�3��iy��Ó��`�~Z�sY�ow.���6��ch�P��L>T��*��A�����[`!�Y߱�%ü� ��C��*�
�)pJe�U&FZ*��Q5�-��*�xh�{q:Ӂ����I�q����D�
�~>ﮐ@�Ӆ��!%�;�JYn4W{��C�'�O���1O�S�8��)P���S@u\��)Y��~݄��ټ[��_���l @���� ��N�H������O�o�G�E��M��I{��G�َ=04�G�DW�%�(�)@|㭓��t�£f�n�f�����v�"E=�9�Z����b�
y�'�/Co�lN�"#��5���2[����^�·ZtZ�e3)�C�a�p(��Wqϳx�a��c$��h��'A�jHnR���q���ϧ()�N(eV���j��y���2ᴿΓKJ���z��|Wg��_J��ų&rYĨ#����f��Z���P�(.K^P{N�	��U��
tW��(]���9�/�4��C/�ݧ���A�|�l�&�>6�A�y�B���������9O|� <5��.a�[ɰ�8�L��xcR��i:��<�+�vZ�w΁�ٓ����U�4/�KR�[!D�4Hֲg;�~!P��c�:3]�oؔ���F���TC�6�x�5�;T�Q�}UN��[mY��_�O�f�fBU:�^N�c��S���G_�����Ӫ�f����C�:q� ��&n�S�����ӷ@�	�?���}L.��@��!Oh<�- %(j v1�t�b��oX}���]��Stg�b�C�i �z�.��[ zO�E���d��Q̱Gy���-f2�n�eI��m���p��xbPx���2;�^cL�8;�@�ɠ�;���A��Ӭΐ�\��h���~��G05��2ɚ���s�{���7���M����Ai
^Yb���'���t6;(�D��FV�t�R�hZ�<c�{]�ӎq��KaI�M��=��̓��6��	� ��!�_���n0t�]���z�-�'6�8���a6>��,�M�B���l�Tq�ݓm���3F�zq~*�^��Iq�����k��n�1C]��4�Z�)��X�q���.�K���V���"�K��J���/�f��{y"P�F��N�tL�����"�h3�Ğc+�'ɨ�LI���%_���͋eE�3��H��+���q6�`Nƙ�e#	���}M�o"
��b`>J�(���d��H
n����-/"m�}�պ��p����J��v�a�G<�������C�>Llz�w�,G�i${��\�����
�#�dZT��-ǰ�����PY��I�Zu���>��5�ph���+D����nj�0j��T�]�;���6��6��O	s2�#��D���M������\F��Թ��ӾΖ�WJ��Ξ-^���'d�͗����b�o����c��˥�	r�8�o�X>N�������1�p���XΑ`��%�P�^�K��E�}���5�z��/�{ߕˆ�}�,�%H�h� 9!ƈ"��N7�W�L�/�fF.�9UN��'c� b�ʴ�X��g��GQ���FS�x��G��fb~��~S=X��
T�࠶�1iX��+�!�AT�I �X�_�k?��'T�B�4�b�.�iY�2�c�,qKC��چ30�d���>+��+^�����K��E	�!<�a��1GPN���j����Z@���7�5��	ڱ�?��襕8l���-�З4[6��yiz�[}Kc���v��VB�ʸ�ʸw�5O߿ ���{h1}�%lA��.+�e��=I�A����!A��=�%�V��*�˒��VE	�kDX��ˉ7�<Q�V?�`�{�djo:"�"�|��e�)�x��������~f�n,���Q�Bp���V�L��̩�:��{��zR�/ӒP��T�T8���k�	|J�	sh8��JY���8�Q\w��ru�dj� K�w>���>	�|�qg�z�3�a�$�w@j'珘b�)�%�� .�@��0)�sm�g"����$�D�����R<�����j�~m��g!O�kV�ނ,q,V�`}�Dj�j[t�i`�)��yFK��U�L)�E�BsL�׊��x�ٱ����е���B쬈~�\cH͑�4h9����0�%*C�Մ���A�A=6��hj�жl^d�J�q�$%���2�����(6�F�;�P�KѼg����߹KЉ9>��*C�zf�K�H�k�/�l�'����y��Bc��z�z�)`5:z��	�w�<Ik��=��Ka�(�K{���[�_�-0`��Nxu���^�5�ue�$/ԗl��]��Z�GSb3S��ī��z� Xg�/�9'E aO R�K��]o�8Ҋ���]!�?p��3N��M��O�ԕC)�p�5��L�d�5S�Xc��K>�geE*���?aн~��8$��؉
�Ԃ#�Wp���;	j�%�I9~�F�=|�d5���h=�k.�!�Y}���x����L��1�̇x��}�����iL^@8}�ԩ�#��gS^P�)x���羊�^,�{�Ԁ���1� �~>�:mrˢ�A�N:�r@W[-ʭZ(6����%��r�pfd[\�qs %��$�{�ҡ�5�/5�8�뀼{X���M�>��Y��7W�{��?a{U%����s��)RI�~���фE(��#�값8e���Aci>	��D�DTi��LH�ѥ�[����_꽼v��K��a������ж�Y00<���i�z��L�#7-rx�x[U��藝���m2*�������e_9Ixs��2w@�0�W��CSߩ-I�J�i��QJ �C�����?�/�ŷ��
�6��(�kEGf�����^���ˍ�bAH�8
���S:����l�
��_$�7S@����sh�h,k^��f?�f��؄Gu�в$�r�����n/]x�Sj��b�̦ta�����eLꑻ6U]�,yp�����q�����\܃�=�0$�1]Q@3���t$��cNYC�y�z�iX,Lc�]E'{���cAfJ�5��C@�ckf���)U�B@��oH_(
��|���v��g2n�c���xGkd�+A��/�It��G�3%(D�P'���&)oI�i������[ �~��v6��hJIǰN��Bl��.����'�gj�I��V�����;$�8�>!�H��Lp2˾g�����P�0V����r}/s�&��H��)���}��4��p��Ͼ�T��%���=�6U?�7�11��u��6��v�8���Q2�>,�RAT����ں�8��.!��a U��(�����G$uEt2C����u����h��\�ȩCA?TT�ۍ���y��������OO�,!Id!�r�Q�b�#]Z	�2�uH�F�(%Q[T�ipm�]U=�A���]$̈́�es)]|;�al��_��	��r�
�&��
��*K�p�)�����~Le�v�B�b��t�q�t���R��"�e�Z'SjӪ<˾k���mh�VvI`I*�!�oy�������+,}0%rۈB^˵L�[8�h쪑��ؤQ���R��h�0Jġ��ܛEj�V��_s�A'�!9�M������T�SSq���������֍Ma{O�ɒ�t�/��ѩ�>�E��̑�����e��]; �h�c{LK���YF�{.��ե�r��p�b��y���oȌ0^P�ǂC�Ap�������0a����0΀J�t��p�p"�R��O��<���aU���eu`���))��K~4h_��$�u�DRY1��P�lr1�N
4&=h;ד��UB��@�QH*���IϳW��(u$��hL�ϼ�����5t6����mbO>��9�]��]��àt~A�u�h�P�K��};�vdR�O�C���ǿ?u�5�觴�@�����j֯����%��s��~��_aVpqD۫����P�9� ���
\���v"����eV�������%���;�pɖ�`fƤ��B��h�]��F�Xi+��mK��^@� Ph���M�߬G�89�@�7���7����2�:fz�KSz�Y:��<��y�!�`�rȨ
r6������V�8�����3�=ʯ����5JSd
.�S�?G	m��Ї��'FjҜES��^��5�(��Dj>���u�<��S6��fMwR���o�-�J�:й�*��[�K^Ff7h4�C���Jsq�U2Q����@����R��fyZ�g���:<����Q�F$6�L���;���I(m���x )�F�۝�n�`H��O��z�'adSň�/�y$��MP�Ȥ�-������:%O*�@9����NQ�04��l��@_!K��O�T�@(S���F����%e�{����wX��&�^�
Ȩa��7�Eq�����>2��!�i�-B �[A�uB_9ܾV�-1#Jը�0�>A��Y2�ªڧ���cQT��� �_ܬ��������x���4�=^����*��%6����|�|�H|h�����S�uF�3���ɒ2��U(>(�aO^��%_:���ߏ��b%$9�Z �:c�"H�V�3��d��i�_�E7y��?*����L��6��&�}
eb:i4��d�����jj��ҧ�Ȟg��kR(	�Ox�*������>��F�O穘Ѓ���<B��`���u.��"�Xࡵ�g}p�}g��B#�Y	B��hM��t�~\��~�����ɰ��a7��q���w�$���� oD�jի\a�;D p��'�r\��Y�\�ؓ��*s��ג'Z{"��fbJN�6�d:j�5\!08V�J���]Hw�3Q���F$��JmAŝ�}���o,:~�	7w-=3Rj+k�3"|` ��]*uuxew��$>��;�~d���*):�^�I�5N� ���ð�P���F<7wVPQ2EWS	푁ͮA��B�����<v�F�j��Ok����xK�;]^S�&�m� HZ��|���(pv�����j��e�~�hN�\��	��h�����B�s����d�}8zj$i,Fغ㩵F{,�;J2�qLԅ8�x� IK�j�J��'q$kwNv�=�<�.��Q���[��K�ǚ+t	e��Һ9Q�z��d1��d`���QYM��e�
�%UbS~������yy������b �JbT{x�jn�S�W@ux7/�����p��@�����t&.U%�	� +�ׄ	��C�[�G�h�>T�Aq�(U�]��]���'>���h���т{t攠�i�墌՚�����9����;Q�dն�h�T�P�1W9����6R*Ĩx��*�:���O����D�v���I�rt/�X%!��Y�F\�����WIMX���s$%�_VL>"�c#�Z��a%�ۧ<�*L8:x�b�Ńq=�$�v���z(�����RN�Jvi;��Q6�7"t:�> ��֐�:sʾG�^.�z�� �3���%/�Ҹp��QYmT�[��8VEk8L��y�E��m�g����M-ԋ����˕�u�,
��xې�>��a�o�q�~Q0�gc�F�9!��N��(�|��{����KAl��Cd�A6�o���;oI�r�*���h()
k_WqB&~olq^�wS z����~/A�Wf�s��i�=K�;4��`mm+�aYNOw�(��=�_��<2�bn����G _��˸�$��i

)V:����� }��)�Z��6lɹ�L�Do���0���j�m���`�K~ �%��j�*T�r���8��Q�W�EW�~����"{�!��Ӓ��Ht����R}���V�:~�8��؈S���h,��.��!�y����W��;�!�P� �<�T���?0p��44Ke��_�i$@�����~'p�#̚��i
[ʠ�A(��꾠�"Y�R���a�S�VJ�	VZ�ޕJ(Ng�[$צ����-��#JP�&���!=Η�
���UR�N��<寐i����o
���NTف�/��!�g	�;%���ٳ��&����?�Y���?���\A��&ɾ�K��0+'o`´��?L��� �|�4���$,i����st����?���
BQ�7/T��	�dQ�5���z�)IAڀ��O���*�q�@*�\��	��N�����ZE��Uj���6? �f�џ��8��(&[��s��q�čh�h`��`�����l���T����� �WhוZ�m2�˚�)e��Yx�6P�nF��}'�Y��j=L� �W;>HD� �n��"]@7b<Ĵ��	�I��𯁝7qB�L�	X�N���%=��o�毑OV���#�	c:|<[bop��iN)���[W��2Ʃ��y�����@*e�o�G�=���M�]H�y�|hVأ;��)X���F��C��lma9]!ּ}$���z%ځ���qnz(ͽD�98�����M	�=4d5624b����mP#EJئ��:�ɿ9�7�x��"4��pL�]*�X�*����vWH0��O�M|��Ϭ����n����ޛh��1���_MrY�� ��L�5�����߬����D��^��02n�Q'Y9������(�RB?CuO/Ze�ތ_b���$�ה?��!,���� a���#@�Y�Z�����jǠ��-�������d��on�`-�l��xm4a�ЬV�]�]�e��ho�	SG9�D��DN`�s�3����w�38ښ���<��,Ex탛�8�$E���y`�>�!1��c�NJo��W��iKT>�8��'pٌg.hq����G��<�qm}{�uZ�'W�]|��.�S����R	PR�O<[��EV�6&M	[��b`*��{�<\�
sv���������l��-��ǘWzhQOEf��wI���=��o�L\*����p�k9����L/�ī��t����K�UݫL���G=���b�=/���A��մWS����a����#:��v�a�d�c鸶eQ�h�
	Ȕ��{���< ���2������kr(2Ic�i��n�bp��m����0�ڻi�
f�l�@�%�C?�H��e�"@^�~��u�s��e��g�SL#���y6���%���1�H�_R�Q7���߁��!q��	�ޅ?$>������4�*eYE�g.�Δ�H(���]�c�?N���֭o(����sQ��;0�}�J��'��L��PfUq��z0�	�k�3��՛X�r�d�D�/���A�;evs�z�3����_�ˠrAD`���o����C>�5����ߴayn-r-��5�dR�h�Lƫ�MC����
-u�U.G {vؓ�L<��`�PF�v:�L32rG�ۿ����Dj���b�{��0W�������Yr�=gT��AӃQ╵�9���7��p1"�͈���i⼭�_�����­��#F��o[��t[���E�t�&�1�V]d�#~��ʠ��z��sʲ�%�ˬA�F~�a\�s��{����tx�9@ݯ�I�����J��aP�DY�����r�+0�2hW\�^Ȏ!(d��~�7��G\IВ}G�*yזH���(�Qv�r��,�&����!J��
���9'�f%�o��>�K�������E�.�ΓO{��д6F\�d����ia���ɰ-�(�:�\���U�V�}T�o�{]���pr�=�^2󫴴N��^�X�<$�p�������8Gg^lH
Ś5W7=Y1.�2�񄻙�&�s�=�m�t��QX�+�s %}��n ܣ�#��8���B���7 c�z��$��"�M3+��(�ߵ��Nux%���X��vߠWLW��V�L����4Y�LwU �6����=o��E�D��X�E���y�<[ù��Co
�ng~�Έ�:Z)V�,�wj�+��6f��/E.B�G@�΢��R�rhɚl�y��!'[0[�5�+R�)�zP[�7���Y��_�o������ j��)�ܭ��b~�WK;��U�Q�Ӽ�Z�#u��^6"��!.����4%Ip+�2�+����#����\ {Gk�+�u���4&��D�~�0�	t<�tf"k���ȹFCET�|�R�S��0ȳ�+���_W9� �ٚ5��ڎ�g��K(�>G�o�1t5�v�@3�T��!����+Ǯ��>�I̩W�_�¦���<&��շR#��r�jUk�'�f�
����^O�^̒��y����en���U��͒�w1bً�m���ց��0O�Z�P]���L��W�V�n���/i����a�	��PN�=c�b>"���P��+��,Bx9�eź\��	���!�*�B0F��$������W�))����{�r=�9�w�Փ^}D�x�'�w���?u�W��I��Ne�� m����������f[����խ-��
&�- ���������sK�����zE_���g�5,�!ȫ��7�5� �Oպ�g���o�*&|�q��Ffu0��y��Xڦ+�R
��<����r;`��4�WD:����B��Kfj��Df��x�]usT��`3H�/�d�s������k����_
��R���UyĪ�G
U�g�o�+f�(� ��H|(��YI��|(R74�N�(�g�)hqΧ��Ԉ��^]��ٺ�_ 	h�����������B��P-���kGG���v?�7��Ue�U	N��jPT�.ip��񅷷���(~IS(��3~F�o�b @ ����x�*�r-[������.�T����p��j!�'D�Egpн&�^�P)޸�=���fa֪Ɩ}��xaZR�U/3�Sh���z�c���cTٖY']�W�y�Q{�ź�%�g�ϴ�}{t�-֌��1d�`���3�P�A���i�F�n��2���<����/ك�(8��!12��GK$�(o����!�}L�&c���U�W�u�MI��W��J�(h7�~��c �X�Ե�<1KY��u~�����r�8�@�����N�:6��-a�Ru�CG��1kE�"^�u�A浡L�/���?q���L,�5k~�������b�b���?0��W(�� �76oCG|[OfpR�]>��K��_�O)GK�ˣU��4��xEE�&�$K����Z�F N5Ǯ^��,�5T߮����c"S�+IJ�"�\����\�/nE��AKjs;�ρN����Ӭ�Lֳ�����㬲�o�Y�K$�sVq�|L
b"��(}�G��ݦu��92hq��29��9$��#z��la�O�lp�Z��S�Owc4`Vg��~��>5���T���B�����*g�+F���g�'v�р�.���Q���x��G�ߑ��h��MF�XZ?I8�� >�'�2��zVu{���@]#�t��p����g�μ�&|���<���j^��e'�_�������ЄO�V�w� ��e�b ��Yb��,��0�����Fb9��~��U>�>�����~�$�d[�g�!ϗfJ�pv�ϻ�>�Ğ6ހ��һ�24n���}�2I5�3�?ع�w����!���.,��͐L�m��
���Do^��q�#u�~6���R�\Ӿ�5��G����aN?#\��!L�fMu4LU��t�� Qx<�'��xI~���o�!��%�p���u�`Z�y9��M^R�wCZ�S~��	�P��򐠤R�'�IZ���ߤ�VC�`��{�m�c���R3%Q��]

���#7r�&�	I[�Y�%3p��軹�z<Gz��VĴ����c����Q���m��v[�N��ǯ�n��^"�s���I�z����#k������_�,Zmy
gs.nӧ��N�՜�<�K��&���?�}��~^����ޞ�c\Rq�Y�*��rڼ�ڧ�вe���Ͻ����x���7���!�f�G���u)�V�V�M�Kn��u�r�4J\�8��ё�e�[<�%U��>̢���^�U{�;*z�t�Q��PP}�'f�#&!�y������[<G��p�x~7�f�@�?�n���|̇���j��h>ָg�L��pC�i���i�������<��Ml�o�����E���qR)5����(��Y1�K�p��%Ue����)2Q�>�ٯYiL�ɞ�iQ�^�3J0�8P�F�%�7g�:�s�����{��b~-��Lf��1�_�CZh��Sv͂�ʣL\���Bɫ�g�
86X��S�����R~�K�����~xZ�g��<+_Բ_\n�*��4��-D��|G���}$�{�$������?� �Tw%&9���%��i�΁]&�t���D��H� �em���/�
�q�4�V�.���`��~)ۈ߬���6{���~^ZN�9��*����G��}p���(�FG�,�Dg.8��PǫXk]�g�}�K�RQ��hU�MA`���',��m�o����єq�	es��wJ�iɍ�QB]��9�~�O�bq6c�:Q��4F��ȕ؃on�nd��|X��pR�uR�pہ�R����`uZ�T߹07��k�=y|8�y��>:Ϩ�B�-��1Z��b3�,/��y��{���+S��:u��'OV��ZV�}�"�k�?�}e�����-��v].��d�ȡ������Tf��R55������ f������s�&(������wП��#��(��n��|����0�)�ɳ���cr}'.uC�O��D��5IL�L0Vx�L}�H4�.jb���:�7�����ڒ�У��4�	�&�Y$Xf|�����r��x�!�j�Si�Ԙ4�{�≒7slڊ#6���e�sQ.����ى�p*3�$6j� 6i`�Y���*���F4��Ll���PX��G�1�G��p�n�D�#�>K�F}A8�6��~A��#�#��`I�䊚@�*:�����R������W.Y�3����K���#5g��1�l��K�{���dv�vQI�@���:$;ADě�̟�QJJ]�� �M�������z��4��2�\30�6dg��)x�v������;ǤJ>U�����'�m.1�>t�M�l�;�|��-���X�W�L��f�!�H��2�|$��xVϐ�uQq:m]�HLA+j`��F�D�\��Xy(J~�)�{)8�A����� 0�̈́��`eK�i�8m9�xA (�@�d��d�i�o{LĞ�8�By�G�H��:Y'�MjR�$����,F��ߝ��A3^�!Q輖��!s��H�~��-?�Zm��#���L6�6:�����,�f>k��n�s�K�Hl��$S�wt�A� ��)7Gae<�K?�AM���y<���&PFeZ)�� ���|�M�S�+�%��&��D,sPR{߶)r���w���*��cӚX��I�'9�D-��z�t��X_�⤫�)h{Ј�D�KP?53k0*�`/�gZ�r��v���_�1��v���v�2��O�Ĉ���t�c�t�܎��MyZ�{wmB�P���s�+���J:wS���[�8/�G�����׳5-����
T-i�I��R�e�4?�������#[�:��'��򃂬���| �*�k�@�
�h�%F(�r�hD-���#�X��X�n(��P�3���v�E�!����$a�Ԋ����2��Q�Wn�O}��u$Y޻N�u��LRu�+�W]5@V'��ǩ�Nch�j?�$�7T<,��i�4��gUj��;��Nk���[��V���N��x�����;;�3��Vf;a@f�m�J��3��#W5��ۡH0��G>,bm�`,9�F]��ǜ��k���Ej{���©�>�6�7��퐢�/w��v�Y��ɗ<�<�g�&���R^F�<4r�G�S�<�$�Ϙ(��̅%*nz��7�%c=/8A.<�A5��~�m��aAZ�o�k��`�̔jB���|�9 ��<���K���?����#�w���;���C[cC��+�1�?{����L�}�N'�F4^܍�T[/`!�b2��#'�][K.���W"��c�Th��UZ���������� u��S��n�ZpH:ʔe����i����9H�����:�*�_��ȚF�9��!���B�S�,�E"�O�`D(��n��n�.p����N�X��C�%��IΜpϚ&jb�?��	��7�u����,^�Rք�{�k��&��mL������^��0+�{U�t�x���\���& �a�R���v��C�Dk��Cq���Z�^�Mt��\EE	�O`b��~�2�6���7�CNu���$?ve�*S1���%n��h�0̿Lf���D��0�a��Mp�����}��sg��4��^����Y���QTmZ�P�������rL�_C��dc�ݕ��{|O^l]�+��Hd�=�p�� +S!3���M�Ds�桍�g8�2*R�w�D>�s�/���ҹ��=�:���ew���3v���|v�i��$���c��c��9!Lo�	@�w�Ym�}����i}�MFڔzF���$���Ke/�";�5�DR��;��ۄ���h@���O�D�,Rjb�����JA� � ���@Ǒ�4�f��,���s#���Mg����k�-�HX൸NkM@���o�!��@� �ٲwl�UBl��w�#�80���gg�\1�RG;/Yּ�p��]@��;-n�-j�E�FtX:�\q����E���'����p�)�=��hۺ9���z�o��u8$���(����)����FO�2ɒ����U{*U-����Uo�\ǐH/k���$�`�BD����
P�0�	O
P1��\�m�H�u����8ӀJ1O�7L<ߟ��9�G���5�9��9Yw���)�F:ns�nNC�훌�y�!ׁ
T�W��]�#jzf�aE��aДWL�8̏nԝg�^e�x���&(������9��B�b�`���<N.IN�c9L�mƏ�@g�rԲ�:m(��w��6�h`\l��Oc]G�L��w1��$0 �P��2��4nb]k�K�E�H7�z�RS�*}a��spg^�o�S���bŜ�j=���gk��?U��b!@���p�(&��Y�р�1�����RQ�޹�>����1cU[��fYX�F4do����K�2*u���$�ˈ����B�dX���fJۄ�Y&2י�X�?�in(2F����^�2�E4�F SU�����7w�I8�rvcq;�{h}B��'`�1@}_ӥ)���y���G�����"v��i�zb5��!�}r}��k�M8gH�X�ʺpb�<v"�����WH�����A6�p��[�Ļ�u�}Mi[�7��[��!Ȅv�v�;F�ꌙ��Q�g�Ò�2vR��n6g}L��U�j�kP��b���r����<S�Vu��p�;���1�U~������~���Q��A�?&1N��D��f#u�)��q�N���w��HvJ&�v��&���#a~V�ʤz��w2fR�W��[�2{� _҃���-w���ioB!�ꋎ��0��8E�����F��~�k���SЛ�>�JJH5����s�����\Vz���p}�����P�cKw`�Q��b�~��N��X-�T���)R��:�,,,��d�zRָ2Ǳ5}j��u){��Gՠ[�����p9�|�u�!Y`�(����YQ���J��~�]�C2!�+9q�u�w�E�7�t
J��!� ��4zX%��٣�w�y"������	qL�<�Z��:s���y[�t�CFЅ���������8��+�PU����AV�A�~��e���Q���_�����*	w`��I�+l�3�E��8�{���M���PJ@7������:t��#怉�O�I;*j�ބ;}�[�_c�Zp��W���QE(�������Iy�
��"����YL�>��]��R���1]����F�%����I�.
Z<�\@S'Z2�
��ֱl�Ih�w7ܠ��:;���d���XH=/a��n�u?�^Ws�# :AX0";�h�x�W�lhus�H��p�v�YW�Ču�8N$}-�����6�
�ºY1}�^�����S��uT�GS��QX�����.��g�����mK�>f��v�9�!�H�PJ(�5-`��2݂ �7r��vZD����r�$3Z)J�i�wڿ�{�|�����qp�qL�*�������k��6��B���D��屙�0�ʳ�}n�b�)r
n�	0�Mv���9<W�B����[m %&�� /�
ܕ	�w���٨�I�SF
ku)��v�fѐ>�F�4*��XT�tc��D�����t���V��o�XA'\�@����l�h\̅�{y؊���2��-x��lJ�kg���s_cO���f5�1�*�?��#Nh���f�
�0���0���:�����bW3$P���7S��⒫=}$�t��Ov��j�B�VHׁ[hk��aӉf�+v���r� ��Ś�*_�Q����sf�^a���h�bg��'�O�z��_;
A���I�V��d4��e)ny<��3��
�r�WI��q!l�HI{�nA-C;�n�'���%?�mj˨]�s�Ar$���E�����ȩ���23�Aq�	��+X|q�½�)R��T;Y��,�����b#o�Kna����U\���3����ͅ5��Lc�98Θ������	�1��� �VMo)��b� W��xb��ĳ��Y�Z�V5C1��9G��
s�_����)z��0���*l�L�cn}B�x��]@��Ժ3e�-#�0[^�H��9?i�.e�N8 �"mZ�&K+���!�1�����Mv�X����e�%���:σ�R��������>2���~2*0�_��Ro�i�z�f�"�3���I�Q�n5�Qu�@"���CD��\:�x���	�?8@������!�2������V<����a]o��*-�K���f��S	�����+/X�]�8/�9�1JX�O}��3
B�ٮ0X/2���"B�BR����j>��r�B?`�4�Q�������ܶ[��Y���߄�g�"�b:U��d�X�f�w��Ř�5��U�;p0��"z��Q~�ewm#$8����ṿ�`Ҿi�xzڕw�dQ�@{���d�z��_��,%6���g��gIv����;Ò��b���㠼��+&9��\�Q����y����e��ܫ����E��(I���~�"x�x������[b;���������r����
�H/���1�xW��� ��m�9e��/�!6'R�:)>��z�+/�6VL�Y��(���XS}�[�%4�=0�F�2�2R�d��Q�`Iդt���g���~!B�ԇJ�+V�!��H��㳈sه?�.����]7��h ���{�ɉ#J�A��>�Vy��^��т>2����a�j�H�8�ܛin7�ͽo��QJ����p�џ���[�KwQk�E{�޹�@t
���@�Yߓ�L��� ���st0z�A����f7��0]�!)�P¾��ަg3Z���pd�Z�%�W�<�2�ba7����̨rSW���P��!��p��g�&-9�l��d��UV�x�hC4��� ����<�N�T�u2ĺ����|y����7�7Ev`�i�d���o!�A<���4xl�r�ܴQ&�t����X�bҺ�pq�$(��8�
R��ʹR=K0H��S�t��rڤRV�����;k;�q�hv���G͆�H�˶���q��.�T�!���e�L���>}J���1�:���*�y+ 	ƛGհ�DQG�	8��Q����jU��[;�T�=�hw0!N����Y�!ay�iT�N��SǴ�~׃<��ử9��ů�fC����Rwi+、�b�u��2�:�
8��9�KMk���U'd���{4��U��A�s�j��Xi���9Ȓ�.����i�@�2y4`�*팆���,��-��2g�c|���pV�N�.��y:XB��d�(X���\�(�R�%��:63m�u�(��275#�E��z?+�#W�I`	���6�&Y��B+%�$⾯�y($IW���MpQ����8F|zLg�����F,�����͡sx������W~CE��g��pdb��UR[,�J�9�;��׽NC�%GXu>*���Lil��L��u=s�w��Z�9���[�8)�� �Շ)Y0���kMl>v����_���>X���X� �	C���C�������)c�ӽcH��K W'��K�L�"!��۶��}8�B�a)����K����H�5#����|��D�Q���e�I�qo�.�٪��)�"��Q��[��p����E�楴�׳��0����{���;c���X�}G�w��Q��ׇZ����l`�6x�#`��)�9�-rm�"1��k��\6+��p�3%�4�۬���ԣ;䵛�ݺ-_�=3�L �KW���d�x�8z�x�sr�V�`���GǴ�:�b�_�ҋ�����$�ݫ[0��n)AiU���ff.�b�2+ ;�Y��H͠�P!�7��~��	��Y��zw��_�[��u�����=@h�V~��$-�s�}����u<����Yv�D(��J�Z����N��q�P.����\��ߠp(Cv��U2\�#iip|`U2���q����D��#;3�h�+(H@9�?ˏ2/Y�6m�XK�M�S�.Ѻu���!�K��L�F���P���_��!EU��F#��f���7tD�h�@�s����i����9�|����z�d��Gn-%A�=@�����,Ǫ�l��o�dgNܕV
���:���͚�>�Q�'5�@�f�i�N�*�z?��s�!�"̳+J�ϧ���7��D�G�ȓ)b/����T��l�5p�z`j4y��ir#'9x�F�c$'��X*�/U�A@��H�L(�Md�@yM�Lt~K�`�Ҝކ�����Bq�m#%X�m'g�u�"c辄�/0w��U��i
r5���Vp'�`3NP�ci���-�$�G"D)�-��i?,%ռs&��1�r�xf���E�LO/�1{�v�c)AQJP�d:���!��}p�1�~����Bo3�+.��7LX��H}g�j�:N�r�Z�Qm|�t��P�xB�I��;�X��CNV�c0�>���j�u�Vh�m߲!��m7����s�"��Gh=��+
AYAU�A�j
=�*�ϒ[�+SM"o5�)H52P	e��e�޶��|��-�}�y��|m��H�d�/:�c���m˓��Gˬ��T��xa��;���T �V�=����7��'�(tD��F`%��h��B7���N��lTz}-�ެj�`��2r!g"	�d]p~����c�b�aV)#�r�+/ܿʳ���aS��
aԼ�f�ՓN�I�Q���D�<̃���~C�����{#��~��Y��n-�T�|P1�zoo�̚���[,�c�� ��PhxF`֯��H�`�^���Ӧ�:��24�����?p��Z�W?��J��(3QN)8��Xq"c]� ���t�3��%�qy.��XD�n{u������U�H)ّ�s��8f�Tu�\Ϥ
�j<�rx�QM��K}�m�FF,�b�cg�*T#��]+Q.ɧv��'��,!���t��ھ�{E�����*��(ɿ��B:��rЌvF�
4(Qt���Sd��p[�=��WoF}fѪ�4A`vi��@��k@��z��&d	c���)ߎ˿9�|+C)���v�ד�E�0R����"�O�h2���(��&g�H���
�M�)���#��:ߒ��c���Z7����!��>o����۴�6�,�5�P'��l��Hi�?��WgX콅�w(N�٩�ИK�B=��W��?X�.",���n�bS�/+�����!J�ɹ��gJA�̣��6����e �*1 �Ps̤�7�A��B���;>a5����a�.�E>Y���w�&\�IZ�����<��9��*�-1�D��ɔ��e���<�{��x��WP�^WuQ;��d}M��u�٧(�o��׼+g�ZW��9fBu]���b�'�Dm_1N�&�%{D6������H��������rp��!q�I���b��������v)O�8�ρY��K��6�f �a�r;�}��������`H���) ��"e$�_���M��Ȝ�*���p�v���3��Ղ����Gؾ���6˴[/�5��g[{�c�S"�WW{�)�JBz'=��[�@�*�B��r�Q��1(� ۣg\X�&,2:~j���ؤ��;��z������6ƦxY�u�F�p)]E�p9ά�Dx��/��'~�C�[��-)�Y��Ƌ'��kM�jIC�
6d��frBo���ɿt�!R�_�b-9>��iC]�f�B���(7f#�O�
��o�����&�= �ڧp���^v&��oǄ����l]* t�Vt�� ���M��������J�6�j^S�)���l�J.�v��m�,�W�Vl£%yj+�Ҭt���>�.�h�����`:����Y��ͭl����>AT�}o���m�X+�e"���Z�xrNA��gz`���H�&�:7��Gm[�9-0׾�9'j+�~Lc��4�?�?k+��b����D����EqM7s>�I��F?Q�QI[ŷ��}S��6տ4��q_v�U+#����T�^�Oǿ�ïl��b�$B���D,�ք��G��A����z<�����i,b��v Y�a5\�I�I,�#�2�=ZI�rT���%M OA�9};�����yOsqN�3;@���'��̬�(��W�7)������/vD$=��b�2��ó,�Lz�	k��%��B��t��+�l�7O$`Pٴ�^)@=Q�M� z��.�'��7����(:� '�{�1�Xp�1�ed��;-B���y����YF�OE��Q���BW2
�㴐ڈ)bb��w��A��o�ȃ8�������/+�����O��,F����ˈi�X-^&�()��͆=�]C��ޒɜ��o��y@cO���,1�r��? sW��UE�5�'��6�cGV�E��Iv?���'p�	�E*�����fUP�u��J�H��1�u�/-�p��Dy�H020#�t#m�4~t�dt HW��0�Ea�π����d΃���4;��,���ݤ��ۻ���@@�[��q.=��Ehٙ��a����Ń<�0U%�}��ޢ�Gg�ny#�|��9ǀWE b��Ag��Ӻi|ITj���r�6kdǖD��4�W��L�I�~}�#��T���V�7rE�������_�4�����C�(��k@AC+L�@�Ct��ފ^��I�DKW�K����q�oE��p�5^���*77/�3�e��肒���wmIݮ''k��W��H�W�B$m��#�]�wh�� � �5�3m�u�{����1ی���'�� �;���� F1pĊ����s��n�☋	�הFDϺ �j,�ږ�op��ɥ>��@e�>M�Z.�l�O�X4���S%���]�!�M���Dސ'_/�C��f�3�#C��zz�t�f$ט�V��5<t����dOKt(���'���v��%-��r�秾p�"0o���x��%�rz��Ъ�zr���|�J�Πf�0���uM88������ao���#WS{mQ�������<{��{�XBrֲ%�,p�y����,��2�MF1�o4�dZ�-˵��m�;/\������)T����g�w�gd�B����xP����/� ���Y�����o\U0g?2?b��������)�OOK�RN+��;%M$
[��a�jyZ���1��i����!"jc�3������U��8��{S�ޮW��&^a�Q���@G�t�^e�
G��nW���_� �F��I���dy۔�MFf	і����W�헷�x��8�^��B�}I� �3ôd��o������a��85�ux��h�q���\RZ����3���AIʟ�˭�4�a���:��(��~8��z��	�'������CD�j$s����~uB�hoA)YX��F�f��Ǚ��܁�j�OY?A����g�I�N[�B�l~��[�y�G[)˳H}�a
q�!u{��q��`2��>^/�o����$䭯�>��9\��5p7��j��Xվ\ҭ8�
�O	7��:S8�����Z��(t��iQ�����O�42p���RX\�	L��#�±�D���è9���e.��������Ah#�rˢwS�z��шU���%�(�����@�'�J�.�#��P���'��M@g�)}�:�g��g���$cy���+��e>��٪�M��C�B8�O��Fa[#�٤U1�S����Y%q��\��$���q��sP�U�;�ͽކ�� ��IY��m���ĐA��@@{�W1d7�v]0��U���������[d>��lN$���H���}'�e�z�1��W��x9o��r��o�`���Լ�N��{���X�ef]"�T�U�=8�j¼���K_\������Y���!0X*��v���1d�p����i�T�5@#��qx�i�ٚ����R�`(սI�S��p{@v�Z�	����J	`�M���E�d!��M"�:ݯ�9���墤vu�$�4�(}B��W��d [����z���gh̟��is kEL�7|97�\�����6��*��S6]Jt#8�堮�U�g�/��_}b�V�����\S��$��M[��U@W��$�w�D�=b��3���Y�'��ڗ:9�
c{Uӷ~.��G����L���<��>��⾺�Z���=˾"�̧�f�0�?�˵h$
�Y�^RSɠ}���6f�rx�x��-�̹�,Kx���-�	�dPb�V�_*�+�SL�?��C�i��u����{6xi��T�:H��o�[���\�����z�A.�.̷z&
�Ta!�� �5��B�V$+E���x9p�b��ck$�p�]yy,��	�"���h������7d_7���n�^L����B���m4!��w�W�K4�@¬L��Ej����<�K����G���~
>�%4gM��N�%��R�Ze�S�4��k��!��z���ˁ��sN%�hL�[���F����i>ǔ<�g/4DW i}�۩����c�߾�]f��Y����Y�okG13V�C�������N��o�RR��U��ѧjX}��E٠� �����K��� �d�>���4�V��D�T&Yë*ʽ�g��A�/�j-��/
f���+�J���}5O�� hc{�ǯ��|m8a�`�Oj��䂕��_��ʬ�;`�����(�����?#� v�����ך�LsR��a�<-'x�m������.��N]��~�6�m�䆻����Z!��-�dd	Ë撆Lw���)yt�oA-9�#����[�k;�x�q����w7�gE� a���\QڭcHBX�X�S�1S1��߷�DdW����TKp�,,(�D7��N��ռ�K��ke���;��{��� '�\	��#�ø����{���c!;l��ۨ��3;
�!{Y����h[�</!Y,�/7L�gto݌�jj���2B5e�d����,�ߓ|/Bʼg�+g��=&&�C[$����v���$�69�68?�B�\y���"���9�ɴ�zF�"m"�˹�4n�͸���JQE��%��^�2G�t���V۷V2�&����ވn�.+.�z��@��xXı��)�}�<#@y������2��_���	�ZYn�V�6p_sP��dL d�k�ՌJG���,��8<��A��a�c������M�6��PL9C_��h�}a�n3U���V���c�+���ha!��)�q�cvRD�,Z�N�OK�g�'�Ua���U�:T��;�����u������ALNP}ɂ�>���
��c������Q�V�<���D)0��� :'-��}�o��SٸHͰ,./#E��] `��Le��[�j�����'���IP����i�<�!A�g���AԢ=왃�iR�P�-�0I�4�H�~�O��?����E�=��Dl��:�%�������s�b{�^���ɶ�j���>��+-��*~k����7�S�q"t���N>�m�*���w@���!N��x$������e7���l
�0Ųbݪ�-�#9&��_��S��5��fQ�@\�p�����v^6OW��V 5��q�H����5HIR�ǒǳb�=���4�
�kˋ�XƢ�z���bM�ܔ�M?��Q�p�"�*F����g�q�' p[
q��I�؅AG"!����W�fF}PkSߋh�] ���Q�9��b~Q_�o ��I�Bor��[rꢪA��*�IB6�M��D>�S��`Yi�:�h�-���w6�f�hM����0e�6ϤO~���KȘc��=���~��+H�(�≾�eua-��:���ഌ�E���\'�Q���Ωg��pL�Hkxh�Z8�$�M*��A�H]��rUx���$*a����2"�O��UVۄ�LB�w��z/�=h��~r34��|.ᤲ^�Oyt��pΛ3���CCB`Zh�Wr`���?.��d�w�DM�k�e�.x�}��h��%�B(�A�Ǌ��JFYNf
�����B�h���R��Wlx�>�X��"�ϻ�!�=J���Ѕ(�֣j�,�������/���Ԃ�-�k���tr]W�Y�5�8��`
��6茊D0����R�#��n�|�<�u���!h3����4Ws��E��Q�/�	M��#!�2���Ǌ�#
^��j�4�����3���H\�^� ��9����'	�v��5��S�\�g~7ڎK���y�b�4h3#�#<�aG���>�8$�Q��v���d����o	�os���-�bs�R�o�}���/�=�o%A�6�V����
"�YL���7��~�H�؏Wۡ?�z#�q�^�T wAw��ݕ�3D^���Q;��\�����}F�t��*P�y�륡8�����L�4[�����\C�0Xߒ��Y��+�������w�����$�fj��N�Kn�;!���p	>�+6��(c<fx��B�e���[�%�6�i�y�C���A2CSu�eZ+�\�t��֘��9���|ņU�a��Q${�>O���v���`S�H���3C(��f�7�j܁lB
����A[���N���(k�kX��v���P5c��n9�Կ�2'��ZT�������č�p����� a�>c�	"�E�x����iZ�0\l�Av7���D��&AA��Ԝ�
���
����j��t��TOoW�p����+�\ɠ��y�vTR|�&&����<I�M�-̺�j&j��.���հ�BR*�&'G@�^���[���k
�IeRSU,�`� �p���g�H���te�ϻ:>�>�Z��"��C��%`�lDbLt@�u��X���i��m&�Y6Ը뱥2�V���3T-G5�{
�
����K�Zk�U�|��d
Z�� ���,��x�����P(�yOB�}�S��Nuw�ei��&�T7��LfL8�g-w5Ӟ��|�d��e픚Vd�%Bt�0�����s9P[zP;�} �N�h���Z���t�"ޥ���2F�ː s�����7���L&���/��
e��<��z�Q5��oY-,2��+���<�\�qXo�k&a�Q<�g�UrA���/�ȋ�e1�D�%��2�:�1�tY�Du��QH����D4�"��m��b��^
�S��|�w�z��5|V�.�w���yZ���`��uC.�K�7aU^n�P	��)_5��Ru�$R�8����<Y-h���{~��t�O9�qpLhɩ g&ˇ�U��~Df{j�xٰg�������O�%�]@���N)�im�?~ZCذ�����T���lNC�_�>pP��?�̳����lF�`2��h&�qw�:�n)�Z��+�����4��+z�ϔ��f*�KNI�x��j�ss���GĈ�g^���f�*MV��YU�']�e^�PGF��v�=�\@^/�G���~����o'}$��n)�K�<1��t�*9�u�G��ܛ��� �B<�e��с�L�]d�?��"��U%���SN�9�A�A��p<�@5k�]��J����#���Ɖ#$3���H�">�@(e<�ɑ"a	��d���P�z<��]Z_㎢ϱ����X�G�i[le���pUx��X�i`�w�|����B�g�=�/�<ƨ��l�n�OI�E��z�N,p&2��ٟ$���I�2�nɍ#ߨ�sx��&�&V�&|
��ƌ��Cf \P#�R�����_��<��%�]��_y�@��K^�26��lqI_`;�2(��Ϊh�ɮ�8+[ �	>�)�(Np�Z��`l�CSF����vI��yTo��9��.k_�l�4W�����` ?4|$���!'C�؅�1�5�
@WyE���xO� ��U�A�rW��|��~!��E��ͳ�����%D:SZ��˫�mTع|\DXx�V(6��j�t'����RO��Z��0Sѓz�,�ԑ�7�-OpA*źD%��D�S�%�|���΃�d�wKg�����C=�vgS2L�����jӰ9����N��1>�."i����>WȖ������\��Y�~x�Y#b0��Ho�wF�莉&[�!zw\_�ҽ������s��.�v�os�9Ag��=��?�UsE�����Õ�-�(�
8�6ܨd|�ɂj�cϷ/���QKU���7�}�&���x*?�0�i�R��e���yۻ���K��c�8� �!��@:fn�̦q,�9��ۣ���g�W)��k_����&)d�0U������l��7L���',N@�w6 ��'\:uI����'��_b�lt��;|�XP#�Y����$�
��	�x3��kę������E6e}�q��#*$��*��A0�ir�G����RX��87�U�6EQg`efX��KѢK:��#�h�$��W����Ⱦa��]�������z��U::
�C�$
Q�(Z�F��,(�.��N���'�j���9�$�aQ	L$t�_/ 0�%:�w�2�����a C-W!�䲢�ெ'�ǝ���M�)�M�//�h�ͫ�4*a:�{X5?N[}�(�s,���ƻ�@��o�h������o�D%�˫�BSm�ԯ�[�����p�㡠W�G$���W�!�*_����_\b5�S��"ٗ�Qb�Ǳ��,��A═�ؕIS�OH_�˪k�ڎ��@��x� �j���_%�`K�߭��$�����Alv�/q�@��q�~wZ7G
5�}T�� ���[�d(�v�m��:�`�A�_���Ͷ������;N�2�%�A��hp��������xW IZ,���\����r�Zt|��6w�P�ۓ��y�jV�V�g.���p�@�����/Oi�N�[%(Dǫ,E��-��5Һ�S����~��s���1��I�Z�쭝��	7�\7i�cP����T^��0��@��6#_�FP\n�-�^jj�s��8�|Hum�x3uW?�!n\)��,8�a�"�U�f(�|���D"0k�vO޴qA/JEݙ��/c�7��j�]d¢7�2�Jv^n8�	���C�:x�����i�2��vc�����Sy�gM�t]T��k9�(�F�
�k�mu���9Ut�[�*8���x�GۚǤ��%d��V�:{�V�W�!�nW�m���_$؅��Z�TvZ��6x�j����G��.Y�?��)�~r�(Y\���*[i���qI�bF�	F��y
�����ب�t��?������h� e�r��O�:�4���j,�1��<����s`��s/�,�^��*�b��x2 :����j=MԀW&
hӻI'|���7���|��O�	� ��N��/�li�!��d�,qP���;EBj�}�� 9GHq׀�9uj����C�/7 1Me!�쫖��/S�/�N��,(�G`l�^�{�R��� v͕g�ў��yfi����Dh��?Mnc���ʪX���1�,~��d_In��(��|���g�ޞ��U3.�p�V|���WÝ�a����n�����
��i���
���֜JR���g���fq947I�%ǦŤכ��VQ�33� �o���rX�҅����C;rx_��w}	��ΙX�:^�k~���%��֫��M���.m�"ӓ�4�z�'���X�GdE��9����βp��!��.�ޗG��Q��6��-Y6����pa�8��]�1�o�)M���-b5 ,)Y!/�u�As�{L���g�gA*OO\QQ����f�S�h�:��Xn���$	A���[�`�sCGgx^!�����؇eYC��F:���vJ��%[�Lm����}/4�Z�%r������J'Cָ�ũ&�*e}'�_�(��~0$�]K��S��p�2�<AtƔt���5nsBSF��F껭f�Б�w\�M4qH����1�֯��Z���?
�-�ى��d��*����(�a@�%J�++Һ-RB�ψ�v!m�`>����/��pǵD,;.��o�e"����dG��tc��	��=����%��w7v��9�ʓ+��ћ�!���҉�������ya�El�Ƙ��>�~90}f@�������j��>,�����gw���y�>����V����K�A��)oCyhsY�jAu)�k�
ؙ	 S�}���x���[�Lb�Y�n�)��~��P=4̛�e�ҒjՌ7�y����Wz1�*^�� �U d?��ѵz�W�L%8k��L�ы떊 �/��u���I;�ބ�#y��C*�
�B
n�LwKSа(up�p�(��t�p%�$������[~�����S���i��O�򮾟1:mh���4k�n���zDdZ$��|D���N�ݎH�E'�э�O�?'�^ɬ	�"�S�{�$�F)�/o�5g|U�m;�Z����ǿ�;^��������k��d�WR��:����"ݣ���.VK���{��p����RE'a%NA�Lɛ��8�pa������8�(����.�8Wdݜ�Q���.�aG������s�?spa+��A�c�$6�]���wx;j�I��
�bk�3M ��K�b��q�ʧ6�bxJ�J�$�A�mo��=��_�ro���
�;����H��~Yý�v�t��3��;whd�lL���|�W.�lRT��=m��=�qJN������ܵ�_5PdLk�Ϩd�9�ד����x�^�aXguc&�)�D�L����������eS�{����UN~�i�;�p��"�ږGk{B���X�T#����L��&����y?<�]o2k%��*Rꈠ���m��k��Dx±����`����F����G��ѝz�8���IL�4~6�C�'��F�Z2�=�4mwR�R��+z�w=����F@����=C�!R�gbo�m�s��X���' �<ҟ��Iԃ�2���h>>�3�<���cF&��]���#cT�vނ�����z����H^jw��� ҈~5�Ɏ�?34E˞xQF��ĺ}��{Ƶ���ֆ,Aħ.ܶi#�WQ��՚!>gU�CQ��˅*����S��>��j��\�;$a����_�����Y��/�����r�dnpF1�02ə�_3e�6����6�q��ҠkMh�>�&�0K���3�Ҧ]���i�Q�&Ɩ�L��9�qf�g��Ȣ~8|�P�E���_�WF�ӄW�sɐW���\ω:�%z��1ZR�Ҁ��b`0���pvK5cx/FЗ:aY�����t(��a�D&XD�eW{�Lon=�$v`�Qb|ƐG���n�J���J�+�����n΋l\��L�$�m��Yk=�^��s��A���J��y�@͇/��̗^:�Uiٝ���n%?�HR��S)��	+R�|�_<8����L���+�eU0���L]@Mx ���f���gC.�6�[=�_�l79���w@���u��։>���>����*)��e�֦�Y���C2N)����Cl�C���Y��G�����֫��$Zzv?
��N2�ӄ�#b��{�klo��k�fp#���q�ِ��>=��0��V}�&�_���$
`C���Ix(��B@6��E�bd���f��肽GO�e�_� ��;I�=;H4��F5�S��f�ڑ$�!�d��df 9��q��[�&m���"[���@��1��>��9' xeO9��8�CWW�Ku�E�4�7��tx~ўB�ȯ���bu�U��Bwl�C���p�k��S)\N��~�#��!�!sW�(�ｒ�P��m��(>�����]r�8��g�p�L�vy 	���)P厭��s�t�ꔝ�'J=M�arnJ�����^VQ&]^����qO�<�_�$�b���m�WZ���I*�)�s:Y3BzE�] ��0�*w�C��>[�k:á_#�4Q�z���	��3Cy �e�(���-p178~���$�2xHϠ��e��Ĥ1��,o�y�`�l�)ग़gZc�N34�S�������fůoȍ-cQ���zRl�1Z���-��Ei?���?�H@X� ��^�XM�p*�/��2�Mb�{B,5�i�ȋW��L�
9v�Ϊ�J";K�G�f�Or��8R������O��3=���:2���lU���t��{�::D��e�ɱav�eϺJ�6�-9j��������s�;X���0��Ks��%�y/z�mz�\�ս �p-�d�1~ڐ,7�.7۷�1�>�¢��W�]��i�>�������mI���*��y��ڷ.]C�a>,�~��T�.D��4K9��̅�Xn����s�m�LTu�*��8k.��
��)M�|d�K�`�A��ؾ�+�fz �Lq����ǁ@J�y�|ޑA����p�u- �v􆒂Ծ�w-.�^:� �+��i��.8�G�pwU����]�	Q	�J*�|��?6�2�����=�F�2�T_Z�)���<� q�W�Yr0�s�޴+�ᆶ�k�[���[8�v�j����e��SC;�9�V�:W-J_yFV�/0Տ�I�k�G�e�%�b9�z
a4���P����_d�S�V+���U���蛙��Z���l�,i x��H�����:��LjJfeK�_�$�%�}���)�a�6׸�7����?�ؕ�ۨ �I��^�^��@�8��D�z_ϻ:�<���֓���3�I�k��m}��B����_�AY+��������~�S�
�����E;\���)��1��W�������_5�i-R�L�e��W~/ s���?�Dr�{�U��&k�޸����P)���S��H��}���\f`.��l��$���d����"���۳k�I�,IOJ�9�lV��دg��y/�ʒӘǰd�=&nWv�^�Q#+ ��T���ۅ�k\ۖt�[K -.T4F����L��𦡮�,R��T�~�{M��p����W���<�$��ӧP�ݔp�/��F��D�Wk��� L�*a�̑�(��R��lBV֮�[B��*a�1��4x�w��ou�d�G�_�@�@
+ x���nR�`���\8�!��\Cz��§=DR��~\�ehA�[�D����DH�}�K����Oe�1��������ϵ���W�JJ[Ƿso����i��	4!M��N	�a�x�+f�-���1)B���|\?��M<>IH�q>�8���nV.������d��Р%��oSO�K�ژ9;��[0=|��G� ��ѥ�>���t�
��2��`f�qY�z�<�7���l�P�6"��eN�L�K�u]��ZЦB��\{�����1���
C]
���L �08�۫4����nH�G� 8C#��υ�Z���kzs��������(LI#Uݬyo�H�0���qϾ
�L�v���5��F&�c/z������a�h�X����op�I�@����P(���cMx��!��"���Ds�R�N�=/�䂆�n�`�TJ���NP�-��@�M�A7��|��<�SU�9��lTcl�~��`�����%��Ntj�&�jM��d�N>���7�g;=y9/�=աm�ß.�%����퉓�J��u[Ϩq�=Vӭ����Qy	춮���QG�kh�ß�&�b�U�LD%2$�Wk��gV�l�W����}�t�|��+L����\7G�	���\���.�щ���E;\�V�rs�M�iXX��j!}kM�+3\|����ͷʟ�lx�C��ƍ�(>I�8EݳR ���b�����F�^:��hN	��ɏܨ���4֟H4v��2F����/�*�W��]S�A��d6諸T��Toґކժ�|@-
��5k9�����F<r�Ѧ�t6��W��P��i���:�	�ȯM��x�m�'dщ��a��w��a������<Y�>�,A�����(�r��F��G�Y�i�Ģ尐�1��N��Y߽O�PL!��+���mgh�&�.���������*y��dŜ/��ӿ�ĬDGӋӉ0R+����Q���}Au�|�����u��k1��
�����ƞ��� ��=�w���y�պ�^v�,�5�;$.��bf�7I�n�#}�i{mq�vO1`y�B�̊<��s�r/�QHR�������w���@�	�|���r����M���t����]k��[��1��#]9)�Pz�XF#��>�e�H)�5:B�L&sϭBI��"Q�/W�뗂�m��;攀�s�"�+E�JD��!��n � �h�$��e�Uj�{)D��T�u*�u��H=�fK�W�x*C����B�q^DWc�r3g2�]s.�Q���y�O�0�]����dv����&7Ǜ����eue����0"!t>^ܶ�ǩ~�2E�������Q��D�2��b�hN�5\�ͩ��O���G��KitK2�	��䓔��Њ��0��׵�����܁�+&vV�Nj2b�T0\�E2�ڭ0���h���V-F�~���Sj*��{ �B�Ȃuن֠m�;�ܳ�ڼ,&Q���3P�n���\�\3�=��4�/��4

��(�9�5�3�r^���� #���C<�����П��\���5�y��vvKZ��6���I\e``�iU���(��G��|z	1.��E��2@Ⓦ���~YSļ	���/�Z��*öi�P�������U��߶~x��燷��A���Dx:�v�'w��!͎��7f ����rd(�)�3�LeU��ѣG!�#�����P�^��~�G�DSh>m�fl���y��H:�}a���3;C�T�H5�B\)χ���%5�5~1', �SLU#�q�=��{�p�����Em��"��?��4x ����f1;3*+C��:qϝ�Y@��Zr��(c]w��o���(q��2`E����H�Z�|N���5���yye,j +�r�a"�����(���s<	�������!'�P��ҮB��B�L��k�	�%K=\��Lw��Ɗ�(�w�xCF	M"V��<����f!G���u�uz-Y��"!��jD?2�l.)���s>@Qb�OO��NL������c8G�^H��b�	���-ic��(�\k_P�3;D`�Fz��ϙ�r �>>	�v�/�;������qPhj}")V�s������d��Pu���{R	�Gf�-���g��W�s㵦Y*�����%`�'��� X`��>�奁*ge��,T&����h�Y�,��$��$��_�a�~ct���55�~ˉ���34�h3}Օ����0_B8<�1>@��]�m�Ɠ�V�腗!k���V����^NԻ%��YiN����Ia��X=��Bϵtft.����.�C"�Z�gR�{?�E:]��7{
Vz鴅�H�s�m�q��}���(�o;�ˑ�R�a�׫�9����䤴������
s��3�=����.p�3����t��?>�=Y�&A�Rh>%��*���
����r!�^��wi>�<�8�����M"1Aa�5��eQ�5��:����~�I���"���UxK	�'���Q~N#��D
{,c���*�`��#Poh�V��~#���-Y�@��Ǣ3�b ��E���h�@�e�O�i:�� �ۘL��y�2%�Ϯ,���R�T�Γ4�>j�`�.I����B�������ǵS�j�-\�P0W-om��Z`�y�ܕ��N�;˔��7����')*
���Pn�W>��̕����I>����̀��b�伬����DObtD�2 �a'���.��������5uӿ��ظP�	��G����V���R�)��&��s�z	��X�B8N��G�ֶ+C$g��`Z:5W�A�x�*f���\y�T�I�l%���W�w��wi�R.JR2�G�}���u���&�Q�I<1�XЉ
��$��\QWxh	�N�����G|cy�½���ܵ��_t����Y9�ř#Rc1 �(YH��N9�|#�#y�"@} (��1�:n���|p�6�d��_+�L��4���ӳ�3��L�T���*�!lI:�bP������)�ʙ������ 'a%���WEa�?�@����6Բ�c�p���ҵYy%�-D��*�o�_Qx�����#�2\�&��@�.'���@��똗,��P�\`�����\���E�]JT��Ym�ǍzV�ҏ �[<�eΩ˕o��v\*��ų"��f�@PR���A*R�[ѐ���^s��VzVFҚ_��g:� *��*���
�5�T�<X>S��@�).�{=��i������-jPS ���)nL�E?
�8�F�Ƹ��^��;~��a�՝��d�
sA"�.�S$N������h��4λ����\�%�C:��e�D�c�k=��E�Β��F�BN$Pҝ�hiJ��g�`�Ĭ�@ק����@�xW�)����	�f�ݝ��{ϙ��C iT0'_:_�P8��}�~���U� �������
�w7'і�  ���J��7T�ts�ט��ζsX�5��`���Է ެáQg\˽֨ ��o#��"#�H���t��� �����`L[ ��j
kn)�y��>�Ψ�>WC*lL�QdE������<��8��n�m�2Ml�?����Nx�	�>@*�)a�H������K��.���;��<1"�֙��??޾��"h`�F:|{�'�چL���O�-�?O抩�~��`s��ژ�P��mF?ʑ	�E �0'����(�1-�$���
�Ɓ0����@j-���X+݈po�_o\�n��s�"�җ=YQ�籴�v�Ө���k4��10Z���N�D昒�j�}j���;�8��ơ��%e��ί���? ��� �����7��;ܣAU�� �o%���<�_����i�;oc?�j��A%�Cg;�hU�:~$�R��P����9ߧ*�:�-e�]�9�aY��[�<����ώ��F���蝭iL\�-=���>�0e��k+��Zu����?:zQU�yVRq&��c��t]sZa�h,
o����~e��~�q�l|o�7lͺ������n��"�/�=�\�\����8��A��<>9��uh$�P��J��oo�r��H�����~�����;紽�vJ�����_�E}o
 }�t��)�@B��n��H����L��h�X+��wX�ޠ`�NqI�~�LB6hL��ue�w�
����y؛l�b��l�	��ʊ�XI��J1�+����T:��}�A �aw��Z!�tڤ^C w��aJ�P�����SR�
br<yƤ*��t�P��V^-b����i�񗧫?�����@�	+~Nŕ+���)x����R�����.��FwuV\�7�zKB>��+M6-�5j&2�v�8��uǶ�m��x#�������m�z�^E�3���K��U 9+-;���Ma��.p��61�s�1�-�1���"˝�?Z�����`M��.��Er�̦˔�f��K�%���?�O��9�r� ��£��h���Bƍ�߬�D��⒳P�T�U����\�[�Vt�+�nq୊�J}�f�j�#ޚ�� ��i�᪂�����e
����{e(j����1Q��m~!�9g��7��]j`�>a�/����������{��|�Xw:��x��փk+�+l�φ^J��d��mҚ���GZQL g
���Q�������Xk�+��r0(����5�B����B3�s�SEi�f���/���iz'�k�B��)�� 3����_�M�§@�s�V��w����aY�#l&��S��I�\�t���.��5,���gEJ��M��?��g�`\V@0�I�֏B�����J��R�OC�9Q�&���n�ђH�c�ٌie��،����)|��f�䖋�����Q�/J���xh��"�h�a�rgc�5I�l���j��mp1��N/��7u�wc 2ӎ�r@�����"�?�F}Ke��Mf@�5�M�/������D���~uь�se$�Y'��'iF��F<}���=��/��E�u�x+~B0��-�Xz=v��13:�w�B�mO������{=Rը�O1�-v<��>��e�b��*^�>l'-A�P��}ݍU���(����~(,�&<ٟ]+0��b榎�X�sm�<��Dֶ�2Q|�d>�$�������	ͲE��ykP�R~�O�3k9��'��q�hFX��}��#~ �O�> S�Oa�=սU&�O��Uf����*�c*i�D-=�k�3NQ���`.���w����+�'U�"wAR�%2���������Z1��_�"��R��%��s��]Sbڟ;�+>=ͯE��*sz^*����� b��ȅ�C��@���B&�v��c�O�rB�8��E�v�K&7dq�G�r������c��ӯ.��za��?����u/��%��7"g�I�T���n�KB�@/c��+�`�~��_�k�5UFIj��T0��[(F+z��q�S%��Z�b��i3�eR���m��TG��3G��S��-�AK���f��/�[6���E�w�� �S�F�Z��%;D�yuec3�d���pz�~�3�8����c? c���\�x~Hb��̽y��?�����oD��Z����pVC|�ש��of����	5A�x!����+>�u�*���B���2��rJ��qe��n�W�"��'ݺ�҉�Y��G�.���P���ARN��,��Ɠ�J/`u���~�����h�κ�f�[��v�r�e=�v2�F�Z,ޡ��1�cco�m�/�`1�v�A@D�w�\������|���&��`�� C^�B�J�}h};��;�?�#��(�H�v40_5Ppe�cqj�޲o��{bYiN�7�jqNإ�$�$!�	s�T|x ��OCq�#8z��~.����($��G��̼����|-�����#(k��`'D��MK���ι�^Ӵ֣�}(}�*���@W���`��B��|>܉���]�]�IB#�J|�{�)�/$�Kд��oН��Au{���<���]؛��'��dxH����M�4�z^��"/ݍ��ߵ���ȳ4Sb0�P�R��^ퟔ1-ѧ�y�P�,%x��̆Tx�����d���ܣ\���B�ӽ��7ss��,��A��"��l��a[^�0�ZK�kqO}�{���.�$cӼ�E�<[�
�C�@~�����G��<^ ȧ�S\�Z3"���^i;�e�e�2M	�O1�+�������� {̟?
8��יj�#^O��9SN�H��5��_��᰷�1��uk@�Lr�4G'ꌏ��>�t<�e���R�02i񚻦 ��,��Z��W1�@���)�����e�co�f�6��d�QF��z���S��(��"��y/�������(9A	�EmNM��
j�	Җ2�D������yb0_���C���Є:\J�҈\��)���_��+����W����:�\$���o���~�_+�~�l���r[ؖ���K8�AK���G�r1S�ݑ���X,���ͣ�y��uJ����џ�l�Y�a|PL�+��F���أT�[x��aD�ڏ�Eb��b��[9��-��wφ�y�4���\�f*���
���}G<obrt@8�I�X��R��	)��;�D��?�+u����jC�����W<�+�X��vG������ +u:1�a�UI{=&�蝱�T+"1�UgA2,��IG�q��^�5|f����x�q��BxM�tXqPm����#[/����G[(Ez��Q�c#-��	�W[��1@�.���g��of���Xá��R��%����A�8Qv: "<J}��ۼ�.?=�?����ޢ5	O[�2�'�����䅏���VY\��Ż(�,�
:�~�a��c�ӳ����G��8�f{v\&˻�2[R�>hI�r'���J.Q������l�
&*1w�O���5Ք��΅�㕲�~���sh���X�h�Z��y�S�ԧ��L�q%�"۰$�F�q}\������d��E��tS���U�|%�C�f�=$;� ܴJ< Q�;��\���R���2Niturj���}1��F�6��7���X����#o�a�� S�M��Ty@��:'����C�4[�+Qڭ� �2��:f�����'g u<���Sw�c�M�

��^fUw��B�7��(��0M'�rS}� :�JϦ���ug�D���J�8��#����� �8���'�EFr}�=�F,�ed�wS=�@6J�D�z������6�r�նtn�W�
��_��m�M�{�N��@d�CN"��+��N <yE|WC��XE���ׁ9�K+�|l�254dew����~�/N���ɕg��j���W�Ͻ9+�k���?�4�1��o�_���q�M��J�ь�Ό��1�ʏ_I=��(_�V1лh<���X����ۉIE���z�d�c�z��b*�an�x�f����&�8NA0>jÞ7�RIB��J��Hu�B��z�����B�=�ƞ�Ux�����s+�R=U��2�[�Ï��W�Բ�D�{�сĆ��V7}����]��٫$ß],�p�xs�i��/����N����%����cS�����w��שE�� ś5�C�`+�3�6a����m�;�k(	�>u��?�	-��pj9��xJl4�ϣD��fr�#�}	�o��p72��o�Nd��6���:����mij���b���8
�i��E��BwI�>�̋���>�R�S�là��Y���v�L�1���/��Zh�;��f7��оg��W,yT�5�2+�	�GE	k�Y��)�q �U?�zTc��Ue
�����i�]�i'�᥆Tn��=�_L�������Xv��ka
���=b	*%4�т�M��r��>��y7��W��+�e\B��1����!��X�fW?��`�����?(e8ً��0C��1��V�r����yM3ē�娮��`J�(��L�	�� ���:���p���v�g񷋜?�8��ׂ��=�|�VӳxJ�5w�ŷ���Â�m��k�Ͻ_cRo�;��+��x����%C�chA�3Q�*&v2�weN�LoN�}�_����G��>�Y�9km	�2-��,�˦~�����$�{ա�b�孨ؓ�uQ�CQ��h�Q�v�k� ��a��>bq$����\�"V��~����a���q_��|Ƞm�;0�C��dV}���]Ɠ�^X,0v?����[�1�%�9����۩�տ�����}�C�Γ�G�$�����^

#'[d�,x�
��]��%GӲ���Q�ጺq�Rp�d��)�����۳ :�ȼ���$*�jo��X,�^gآ���u�����#�?��X��l���z_��I�mI�\�Д�k͸�ʻ��吪㨑�Z���C�P��q��F�溁G�lXȤLV�
R�\ŕ~�mTdY^���~GX��۰S�!�H �9b�Vإ{0�wT9�nA�SF�p0r�"ϫ�M�-�D�����e�$֌A���pR�L���j,*s(e�e��O�RG%�m��"�~�k�}Go���A������t�EP;�Hg4oH�`�ܦ�ojty.�XQ��*�	T'�ZLl}�E'8d"[R�3N������8p���~�H.;����X�-�Z0jk٬�:����'I��Y�d����u����2����`�s0q�	w�]CK����L�;�$J�mr�� ���,H���L�5�ń��\�/���n_�4s]�H6�Ę��N���,C�o[��`�ۨ���cTKfN��cvu{�ļ��WnH�2�S�ל���檾 PH��6���H%��
*-�ZA5�i!�;s�2�Q�����I���<j7ڦ��������a�jMf�(��jwa��E<ҷŤ;�DEPu�}�L��6O5ՙ�˿să���t�S��E�JQ�Bs)���N���ȩ���r�r�4-���"^�=��� Ƹ,��e6�\�y�\fx6=�a�$İ�d�Z�ǚ�4�!�}1?<�t�*��]ΙW�Dq�으83�f���Z���9ǰ������E��K��j,B�����S����)�6�hB���`T˗�l��-5!|Y�*�"3E�f���k*��+mߒ��Ⱥ�Oɗ��������;���=�u��������Ijex�I�D!�4bK��,���Y�{�|.܆T8��ԁ�g�:j}W���0�x}."��)G) ��C���PY�DI�Q��D�>����}��0	^�4�9���H�6�n�p�n�f�����?�h��),������s��SB���+(��E��%��_<ԁ���������A<����e��]�c�;�jS^�-�3^i��-��)-/�X�H:�K(����72�>I��f_{�ǧ0&L��N��F�%�O�0�{�i�V��i�I�#uf���K��FS����F%�PҎ���c�F�c(��3i0 �ʅ39����-'O��*w��W��/+ E}D��)'�.ϤG*y�Ҹ_�g�|��a�u��b�ӂ�>XlX��O@su���ށ�%�m�~�;ϳ"�\���S���� �.���5F6α�h��e�X;{�]�FY��T�ھ����r��r��s�L�`�=c�0z&�O������n�K�&v�l<𬉑T�$8~�.����	q��ϵ%F�ri��f�zdD(�!�VF��l�%�����I�p��&ݰޖ���(��
��4a���b�`�}d��!͊���L���)��{�7]+�P;��R4�+�bsI~NA�p�dR�V�&W2p�<�A����y�s��{
�S�������0���F�mp[J�����Q��z��%�P��J��a���NtX�����yT��&��-�w�� ���R猪����U�b�}X�$d��C��Ɂ5�|�z=���x����'F��D�[V��S�}C&����~
u�Nki�����\+_�Q�_���_&�'[�o�]� �]��U��P���;*Ƨ6O~w�\�1��1sb�����dR�
ū���q}��M�?���UԽE�PO�r83�D�P]�ye�p$����d��ÿ�pH�/V�[%�U3�����o�*>=%<��jtZ�����I��J8����v�]4<�Qݲ5�+h��&˵`���z��k~����p�0kRù��{��³?���LR�_�՝�v^�����L��AO"X�F&Th*$�Of{��������iK6��}�Ŀީ�/DҚ�g�wŗq�6���(G`��M����;\<�����͘9��/t����>�
�-�[����� Ɠ �����NU�UUL���m���ۃ�ŖCjCM��F.*�?$�3&H̙�iP�|���t�+��y7�h*��H����e���6��rA<a�vgloFZ�:�i=��EZJ ��nr�" ~h��J� z� �s`vó�`���IC/W�B�-_yf�/4le�3���*�`O=Ԛ7�����/i� ���P�jř�\f"Y�**h/H�w���1����J6�0}y Q���0�'��S��o)S����TP��H�v�ߪC��a���� �	0�yݞ�њ"�Z!ᄁl��qy,���{?��þk��5bX�>��w�?鮆�|��0[�����2������y�cͽO�=1t���%���8|)��[�kZ�v������;���h-*Lv?ց��� v�@�1�ї]���ڪx�0�ӹ2|�R*8�Y�Z��s�����N�hX�zʀ��3_z�n���Oi��5�[����U�����j��E4�ł}�Ҏ�:�Y��/?q�|�4;J��W�a+�9�CV�=�
iRF?�C1U�ttp�>��P�s�VA����뚶��B�R�S��?1���ԝ;��d]�r���s�=q�N�9�T�����cÃ{3+��y8pu�жl�NOL���Җ6|M�h3U9j�.n�W�f�� �g3Y�O��拠
�@U��Qx�
(ni5JmZ�oӎm���k�����!�=Ռqb<�� g�c��`��1E9��n3���ؼ�Rq�����AظTPî�#݆���8{��ʼ2�uH�[�;VF��|�0ܔo�)�j��7j���7��-�#��}C�~	�u!�C�������EK3�x���zе�霭"�}�[�7(u7�"�8�3$������	*H%5����*�S"���n��r��U�K=�M[tp�%���?�E��`,'�����MwO��e5w^������g:9��j��nZ�S�f&w��l�q�ahδ�j	�~� �_���o,�깆<K)�O�	?�x~ƣC�m`���^F�@�~�ZB�I�;b%�Ͼ�X�����}-�ϰ@qwU�#��]L	��5��s���+<k�ZR�sJ�'C:�Es���V�X�h�Y�#��=Z��i����矹%껴�f����V�'+�CE�G�:�?�	@j݋�u�?߸�ү�xǏ��dwh�ţ�n"� V��ݷ�-���E����h�����ڈ�;�p3��W�[�L^� .���t��q��W�fG�Ԅ"����U���[��L��$/<d�,DdH��	�cD�*Vz�	b#��j.f�s; zF`W+�n��P��������?o�ʓ��G�EZ���]A�ɖ4|I��Ρ��<����J@��ٔ�kF�z�������{���sk�
=t�iI�*��83�ż>�J�
H*Z��u���2=��cň�	���,�$'�S#3˲ںz��U�O���ZL<I��op̂йL��U�,V�&������l�yv���L$3��d6��`���Ǹ��!��[��X�H�����u�<�� @��>]Q؎3@��|����-����F��H X)̬���ͭ�M.�������q�_�Ȭ�?��c��� �ѹ6CH�lnmaST�=�`\񻹓qƆ`jW��\U�2㸐�ǭA���+�i«�K�n��d	�	�FKt���ƚ���ɛj�돾4"�ǁ�.>>�ו�F��I'��P��r�}�E�Z@�f�Xu�M,H��
C��X��X�*Dۤ��:����E�{7?v��<�B(z
��w�]9g~��
y�8ps�#,Km��RBX��7D�� xDHן�j~�]�uz�!��&�7.�;��Qg�ێD�M8r�/�:��w�?��d8@j�P���6T\gL�V	��c �7��~ο�����}Yb�h���
���C�9�$�ye��q:m/kƩ$5����4�y&�,�@�ڠ3�8�����K�O�&/a=�f�Hs�x6E"����f��u>$���+-�O��l�����3��-���Y�RVt�� �B|�=�7�,B*�Fz3�̰�M�(�0�Du@o*/�~�$="��tH-))B����"��Un��1s�p�(*�:c�ت�|�~��"�a->��6�)k�	yv����i*� �K�ߖ��H5f���no�6���Ax׎��������SL�x�N�Ε�p�ú4���`�a��P߲c6��V�G2��$L�rxb�eF����P�1��D8D��&Y\F𗪦���FȨ�/��v=J��N�����`��[!����z��?}F7�<�{�!걖��[2���,�:WO�,���MM�h���m�l��T�R��r 9�lNtf�[�3�v�8��Kb�Bc~�lի&c1SVI����S�4z�	Bl�����0{�QZ��Z}<e^�[pҐ\șCF|�̃�qL=�ç5wj��I5�o
��_P�[�-|��\r��G@?ͺT�V7,%ݯB�5XL�INS��<�;�;G�QdL>����B�lL��G=�YD��{���C:,�Y�KY��g+�1�@E0oۉV��F������]u�e�}��YA[(rߛ� ���Tl�����ƥ���D�2�:�Z:*6�}�A��]�_�P������,���y��{����\k�Li�bT�>ܥ��?��X2Q�T�IZ��ebJ�';�r"hC�./0MO~04ʡ�FrPT��G1%d�8����!N�6�e��]�]G`�n���Q����6��3juY�SzU���3��xwe�B(k�EFZ�ib"m����0��y_��߼�ܾm%�_������yo�q7�_#���{�hH�&�����$�E�c� ��Y��-��P�á��9ī��a$�2\�#��X�w�?���f�4D3m:�gj/��,� �����FE�h����Ēk�>@0xJ�krH���b��$9��l��-��q�I�ea5f��#Q��o��	<St��}J\�mV7͟�>�k��`D�C���ƺ��>�{�1�/W��4����.u�$��� �r��7�����As��z9H,?�l���#z�
������|6,闈�����Q�6He
��HT�;&�0��K�`�1V!p9��3�3�XW���F����
t�C��5ꟃð���{2:Xڌ#9��!��֡�m�����3����,E�p�<���Ƅ �dr�8"Ysm����]EPm-/�>���zV4�^�j6@AwA2�*�Lz!�G��O�Z[aE,���~��SX�-`,�jֆ^P9J�	�<"2^�E���c��/2m'gK���^���rU��đ9��WF��@�!Ro���܇�a�S��� �2��Α'ԻwwPj�xc��� b�/rĕi�-��F>�����M�Y���L���f�n�x�&m��\p9B�t�E8�h�DRM"ҿ����l�{'5 ;'C���V�c{�-b�R���3wy�LHY6�O3��dR�a廻MC�%����MQ��!�\R�ou�G���e���*��kFpռm�j9[8p�=.��^�eh���z��S�}"
oD�H��
mP����߻Jp�n~\F�slS�4�<P��,�yE���⹛~�#~��`���.a�P����G���S���z��v��Q��5�@ތ�:%5�O��v����������|c�d���K���T�.o��K�i��t67㭭�fɊn�ʌ�o˲��᥎w|z(��K�� k4�}#���J�3jgN ���qƭO���Q7�K��w�����1v6���\��uvC���Mӷ<�_��� D=ťu������f���م5&� �T�<H�Y��Sth-��s��p�Y�����b��Cn�	�a�|dyb��Z�:e�R��0|�3��_A�6
�M_~8ScП9��,+o�l���,ś9ţ).}� -̽�?����8�#{":�ģ�����}r��I�68�s�"�̦�%)���g/u�Q��r�>G��Sz�s�^� �n�����Z���Ͳ�A� �ydіd��JF���[ �d�߉��?���.q���=tm��D~m)l��U��,>����lp*���;-�7�mu�6�
-;T}��ŪCa��$�2��ȯi�;oO��g�Z�C#?���ۦ�ކ�'�����$�� ��G�lR�lZ}�)=���:-�������1�s�:pո�ȅy��28���_[~�ը�xV���܁B�d�ldG.Al���=�C�;]�kJ˪�<B�/�5p��1.͉�j��Aǳ ڊ��V�b�w����{Q�7ն����T<Jk�_}߁@`y���16y�|^l2t�KN �ar�F~AQ�GO���P#V��E��d���QBh)9v��k���Zs��_�iN�z#U��FZ�#��6d��<�~��X�c�^<	m��*_E�{���--�*�5X=8��A��`h�*��D�h��bvb���
���{_ .�}��xx2t��tG�nl*HN���U��?ڑ�5�_�1��u�RN�S. �Y\7}���������v�Z��"�]���צ�N]o��~����"�$\�
1<�� Vt���갢�����pi�7l�̣H?/Ӻ��k6C�
�����iĢ(7z-s%�Խ�E��p-��>�'m@n˦ˬe䍉P��ýGn��{�׼N�hi���@*'q�Lw��ǜ�]���}�M��DKZܗ��GG���<��n�Esj�&C��*B`+�3g�o�γ����KK��TlC�͋��7F_!��d���"1�gr���T��5�̶�d�͟tn����g�5��e������D3��S�Oӡ�d�v�%`ZL�{�ѹx��M��􍉽�g������{�w��O�N�f}�<>�y���S3G̔n���BiL5<���)��3��"�O-<�{@B�C�}��5e��	a��$>ŀI�|�K,!f�쾠6��G��p��I(�ˎ>�Q��kҿr�ߛˌk9�tE!r�Ӵ}��S>��k](��7��gD2נM%�YFS���8�^(�%Tu��1.���n��hJb�X���RY�w��Y��N�~����(���2X�����妚�K��@.R�bBQ^EE}���!��/jh#4A�)<�%�jԕ �m�m��=Z����и����p�f�~�$�ҝ��
�ے��)R;���M�o{vO2M|eC��Ǹ��2mRH{�q�c� �5a���)���`�Ph&ګn�ͨ[��l�����8�WlJ9�V����zت�@>�ȡmQ��-P�$��t���pt��DJ)m�Imbɷ
:\�q��t3΍���fmk�|х�o�1<wp�<�G*��6F9�U-!�����k�z�|�̠�^1�ͪ�c�Yo��v����e���yZ��à��DlF1���������PY�u�ń8�;����D�k�Q�>w"~���r<nv�待Ls���EJ&�WͿ\��⡪���8<{�Y��uك�����)�&B��(ʴ��j��)5�V�nV���+����ϟ���q���6$lqF,a��sd��h��@(���hBx�ҡF���#T�"�Fh<�+n���8�G�[�j����1� j
�L���(�f~6���:$0���<��yB%�� =-l���*n7�ѿ8 ���Dj�F�H����*@�G��`�r�_��C�wn��u�#O�X��rR?��o_��GI�]Vd�I��,Wn�I$��|_(>x����x*��ܝ1a1����S��j!�"��Y,Љr���	L\تY�F𖏒��/���|0b�R�d����B���*Vر������Ok�	�L��%W3���4�K��!}�l����cJ:O��۳��ڝ�yY26�B�rk���%-t�f��F�mf�ë*�#Y�Y�7}�<���u��j��1�]��+���4���y9ʛfүP)�3/�����Y��*e���8�n�=�^�{s*s�2v��0�Ŋ��eHp�N�A3�#U�kû��ad�>KI�7��
�^yR�+թMXBs�b�8�S�Ef�5�216���yX�W�2q�V$��T�M
��N��ًH���c<h�nC�g���
z�
YC�ּH�Mn�G�B�xo����qL�L���Ax�b�+��0���(t�`��[Z~��Q�Xɓ�3��J������m���.W�� ں,e��.���>B�L�X���	�`��P��Ս���냵ԕ�g����H%��[~���@BW�����
�e�����F�L�/��%Enr��F�s����0�p�Pݖe��%[���]M��O��E�K':5=F6��lZ�W��]�}$��O��2Y1�0�J���|;��v�H� L?�}�˭0��v����dJ����3{v�檝-��g��@����hE_�4W\&(h^/�k�̓�Mܡ�a�R����|�� B�l�U`��!��ɀ�7�߅��+:����\}*�� ���Q�N�<V���t�w��,��[⪥K� �\��R^\2{˥�R��&[:����7q�Z�)���!�&��N��_4��UȊ�X�IZgh
�d#�:���@x����	���{�����n�"�eX��G҂�,�,Q��տ�i\��3��*��퇮xG�4UFx�i��k�|
�E�*����v ��q3з�ٯ��a�¹2x�y�0�# ��b}�'�{h���ސ�`g�ч}~^�b��[�[� <8vh=F���/�^=ւ��д�:%hCn�8)%�j��X�y��Պ��|Flv�T6��m;Az1���|�t{���<�%ٵ�j�73�!S�҈$Q������3�b�ߴ���nc����;��W�FA��F�:�-�U�0gF��k)??�k��Q���ЕB��pjqP\���T&
;�)Eǖ�u�ڥ�\Ż�1��_n~[�Qp�f�\<)�;�-vI)ܲ����A��p�+٧,���'�ow'�fr�.Az1���%KT���L=�8�H2_�O[;3=F�E���յe�*P_�sB^��bR���������:KS��t�P��H����`_�sqdR	ٯU4�Q��7�(a�&�8�o|b�s�LZ��2��Gp���Ѩ6e�hj�w�({W�w�P�+��Ȉ���Nh��a~���C�E�Cq���n�
2at�P���E���,���j�9��V�VGKJ9;Z.q�L *��i� \��[@X������ӵy��@�5|��xJ���d�%��T+�d3�ٲA�i�*�nA�^�Z�?1��H`�U�]��RK?#��f+茅��&@��[	ɴ���<��C�]#m���W�B�hm��Q�3N&3T�?��j2aHz�ɇ����K�� ^7 ���G��%��@����_%�u�#u+�8�(���2N��6��q4�W���WlV۵�=���u<��{��1s�>p���k}Ը�K؛ao� b����5ҩ6d撓B���wً8�)\���c��I�!��c/$n{{Pe#3�����}e�_쇑m��h�+�4�ajs��"z�l�[�T���0zp�&L�j �� �mzm�6�(q���O�]�������˙�A�P�Ҧ.����+4���@��0aӈls� ��Y����:eΜ_֬YW)�x����-Q;o2r��O�?b�O�`n#�l0���qQ��D���(���++�n��ó��/��;ƺaO�($�S�g�	�n-���>Ӂ"�(R+�) 7���G��$7_��@�p)Y���k'�Q�y��(̽����<�lg��<�ͽϨYB�.�4)0aݝ;J�V�e����c�zD��-}xJ�p�S17_AkJh�6������ĸ�H����X+/�������9�-y�7��׭;������u����l��v:�	]��$<OE�/�H]�u_*ZR�d��*�)⠓2GZD��kB�m�ǋ��.���L��.���"�P.S��$���{1�yp"�FJ��e�4�Lh�H�5*��i(�禮�~�Y`
��p�{�1��>"�0�Ag�"�Ӡ�i}3�c�z������	m�������j��������"3Q�0pi�1[Xm�!��y��	~�:�zp0��V�A%�XLzW&jK�*��{Z%.I,�7��5��`�1��k��D�#mXç2?ϔV���Ijw�Y'�I]�0Ҕ	A�3*X3�%f��B�+���cM���?��w=SQ�[pb�v	^A�b���R�"H�پ�h�f������8�cN  J,�.�/�X$Ҁ$���a3i��)�]�5ɯ 9���T�|a�baz4�/�x�^V��'r&*[E�>�'��j�C~�������e|���������7�+P�A���� u�Y�:z���tʖ�x'��>o�,�Zt�Y��U�~jJ?A���B#j�u���Q7�+�e �1/�����@���s繉�#M~����@���9'n��@��6�;�bo�v��둝�D����,
 �a`hB	�)V���3��tȀ�m�,��-���(d�&z1SA8@m`[��h�Ƹ��~�~:�3,��{�|��Q�t)ȕ�+���)ت�Q������rx٦�D;�D�R���.g��tV:�I�1YZs1/���oF���;�+c�f����3*�9�#d�0��b�CG��D�l�q'��Xza��c�A45~�ɳ�*�H~T����|�����3�sw?��"�XJ�S����x��^z��b�gj?:cL�#��`�|��������1Bb@�h�6|�D�Uj��{Z��ې��H������tc��u�h�=k$���&��k��jѪ#���֔S�@TU#�V��S�NHr�w0C��d[��+�U�M_�(��(c��{0���d#�l�d�I����@�A�_7��gYY����jP=�{0���d[����p�OF!d�$�*���Pz�2�ꍣ�nT�h� �/Z9���w9�3�u����z?de��C9=�h����NZK��o���9<U�)@�9\���G 9ˉ)&��!%�ax-������v�b;�D���� �'��_��}+�`�LZ�yt�nS竷� �"�^(�N%��o��VD���!\���Ş}/M6 DC���˚^��I�1�a0W�G�x��8���x�^�P<苽����ܱ�_?Hq�s�ԝ)i�cbhO������破����]H2��İ���J�-��l�d�:��}�`FӰ���)\d^��+��(-I�'�z�N�Ԉض)K��ͭ~�i@�}�"�����ǡ$ɞ��4���q�Ř��ըʋ1���B�<�'㑩[e��)y��/]m�N���q:a��M_>o�]�招����6�
ͽ˪7�i}9�gq�D���cY�'��xNNl����������l��4L/���
Ul��V`�����b]9�Rv�A&Q � �pjV�� �j@�O:�Lu�h�Ɇ��Q��X��\5����W}QT���O�\,u��8��!C�-GT`2���}�E��=�/v*J7F�d��:#�B����=�rhV�����N��W�����kM�GH�]9]߿����`���c�xQ�����L��N�s��rZ6%	�r;㥂�����(������C������~���Ͼ�R�~ ��8i᪺x�V�Oߢ��S���٪!��>�5,��|O5���[.�������ݹ��BGqKw*
F�K����]�]^��[�0��+�FO�ңi���Yq�Z!�V� � !��1l�MB
�,�i�Q����W��P�ɷ��f��_��Ӓ��d�w���~��Z��<��ز�'���x�E�$+����k�����~[�df�ʹ�MI�wZ�yy.����'���)�s��֓��]y������ak�9⇗��w8��Dk/Ȅc12ߔ��,�����Q���;m3	�3J:��.�B#��QC\���"U���[3��X�AB7��p����1���r<����V�����7}t���U��-�+���OX�^n'�שi=/��5����L��#��W跌>�a����c�?�����1	]��U���J�>¾��D-�����d�ۗ�� ���� <Y�BK9�}mhvp�����FXJ	��1a�3	h���P��*E=��
��G��2D*z�kX�|�Z/>J.7n^�_���,��i�R��eK��,�?�Z �x�^�M����mV�6]c�_�ۿf��_�xҮ�1]T��_52�1�Vz�΋�h�g&,��%��W������������<l/�>ޟ�B�;� �o����W�vb�u���e�򢎖Է��̲�����{�����m��.���������"Ħ�|8��aQ��͡=��6&��.�3�ӳj����؏�5��������A�:�I�0�bv�{�e'�r�oÐ%h�Zc�{عAj}?��RFa(�h0�oG
�_�͈��!y����v��7+���4�6Y¤���e��y8�%�b����'j�n��3�o�EU�Q@ J-��8���[�����eq+F�.�S
��A.�&;3�h�$4*�I=�OO�`/Ԯ���2X��t)��"m����B8G��+�m���ͅ�R)\�7%�F���\��^��0hg�U=�����Hz��q1Wo���Ù �o�Lt=�w)�>�����v�  d[������
��C�Y|{%�A� 5����䍪����c K�x�;���>}oU-g�ھ�_��e@r��9�-����t܀�S����+Rf�[X��5</��'sy��(t۬�}�~'���X�e�`'d/��X�~��	r�-ݱ���U
�ι$��xG,�:̔dԓ˵ml�9��V�]ߛ]�D�x��.�㱄��φK��� o�G�T@�t�a� �����Vz��]�X��f�$۳sX]� �x���놁���1��jG��(2r�G�]� lc"��;
F#1��Z-��L&�����Bl!~` ���i�ݙ,whrw�|��c�a7	��G���Lg.�)m)���f�N7eن���-P���g5Yo�X��*k6��R���w,m�E-�[�]�p�i*ZH�/%��v�=��5��~�}���5p�E�,�[��ZG��Pe�~�%���_�;�^�}��͚o;�w\$h	�VL벏w��u���S�
�U��T�@NV�>������ѯAZT~m���>u�_E��M��G�t������[��36�p��{�w�I���湝/OE��*�����L��6���ː�
^O��`ȉ�Kˁ���[O�C�w$꿴 oa���-�3��9A�� ���l�Ɗ��QC��x`�ÜB1���p,	=���;��d�Oɔx���1��#�p��I\��[�;���J�("q�/C�/��ȯ �5-��-���~��� ��C���|���,��	�r��=�5�d��µ���]j�/(�u:����s��.ٹ��P�A��8�b�j��aÎ�Rv�� �(���0옱���
p�������c\t��W��l���o�M&Fa+�d��V�37@3��B]����3�E?����4���?ę'�OϾ���#����T���S%kĕ�V7���Q/y��/���O�ĊQ�鞦�*h����E{n�����������su�eӄ��c��mg�B�)>9��" 5�vY|��y]�n�}{,r��Hin=���>"k�{��(��e����A��l��{K���/�P���]R�3��e���}��D��]�6�WФfU��VT���9��؀�)7eT��������T��5�W�wĀR��Ы`�c����Z_mӔ�?X-�$��T2Y��U�Hv�$/3�%�~�����#�4b��Ew�d^��r�3�ʎ6�%��gcd��q��P��9�M$�z���Z��D�"K�u�?�%R]�ch�r-n�f8��K���?��!��nh ��	��WG��@+����D�i��$G�����E
-a�>Lϣ6��-��O1�S����Ĭ�@��;���t���+�/�v%����R@G2�k�Bll~��Y��%��$���n����\ӑIj;��P��ѮI̪�L%��#�F �6hԧf^FI�T��crF:֎�E�@x�JS<�ٿ'�im�{[�q!�}jh�o�=�����CG7���l�ck�]�cDF����P�F�񉍉	�(�Nv8~�<�{Q�dB[��*�b�������>���i'�GJc��սF��l��_��{�w�� �5�� ?T]o3�� �����n�<x=�^����A%�l}'5�d�����1��3�]��f�a <��ٮr(��xެ�'�E� u�~h�hǇL�u��2\#��Ҹ��eJ����N;��7��6V��]_Z�I�݌Ө��}z҄`�Ϙ=Tb;nMV&kc#d2ma�]��V��2�?��o�S�/K2AV�����V���=�]A;��v��e���xO�����o̵ATa��+��Q�P�wK���J-s�,�/�$c�x�P� O��4���6�%���?U�$�V���<�Y҇#�M�ɑ	ou�&k^�xԣ��u�s^{�h������]��ڭ��T��Xb	,�&�#���y��~���y>�����SɪQk����}5�ip�v(BRۇ�F�)bg�7@� NӪϥ�Ik�u��bJ@0?Ssx��$�PY�N�93��&Q�6��.��aH��7���j�u�zm�Ή�&Pbߌف�7ki*�)ō�c>p,/(�J����@����ȼ=P�q���G!�AX|>a�tƗf���1�{�=� .�@�R��Q%HBr�`~+zhMO@Ӏx�R��s���˛M��%ZBzy <@��4uї� %�T�]�=�C��q�8:á\	������2lAy׶��6�����|�ɨe��������Hdtwm�)j�@�9,��\��J=�XY���f1����h�Ŵ�����ʅI����G@�Ka��*�f��Ξ�[7��o;�H��S�M�;熠<X�&��Q�Q�Xv���6��=%���>�G+�H�G���f�t?Fn�����im��4����(1X:��cܱ���jI���]�����+f��b�����/|�F���>.�ۓ%���c�D�%X�^�Q���I��鞑��@�_M�{Z�R54�рK�׀^�Pl�9�������j�P�N�5��A!jo�+�j1�u?�x�H�-$�pޖG���r��"��Э�:d���dF�<��_8��S�3t�R"�`z�:�7T�1��Kَ�n���)����<%��ŘB����5�A�?�J+�#Xs��h&��G{͋��(�0��4w^S~�G�MK􀠽"3	�5��Y�V�bV�!���LX!�>����r��[ǃ{�I�K��h"���*
dy
�����	-�0���%��[`H�"5��*s�S@~��Y�ࣙ	n9���]'��j�|4��VLL4�@}ɳ�!z��WTh��e=:���E:*�7� �k'������C���1�����hG��j�ҕ�,3M��;h��Z��LWV�~B�*�^S��E�@��ڻY�4�$�=�+�ƝQk`m���]�4:�F�u
 �9�V��ӵL�.[��M�<b9����>�)�I1
 �⇧�v�RG��-2�#
�Vt�
ϗ��R�4s��ٝ������rW�PʔP�D�zj��o��X�ښm� �~mq�W_������.*��:���v5��C�虎.�$>�}o�Ҁ�v����o0�l#l��x�Er�Gx��r���� 6���Y��[��c��N�]�JT�e@R{T�~�
m�������C��{����b��x���ob��w��,.]�썒���Y];[�K�N����[���6���Ksԩq��`��ϙ�­d�����Ɩ_�AWP�Bf*u��$iM�Y������@�ϫ�Д\;y��P4؏�P��YL�QV�G�de*���䲀Q�{�;Ǵ�[�lXX@��۴9����g|�H>]�2�a��K�Ҵ�(e~x�Jjpų��e������p���!�4�����f*�<�h>p�s���[ӫ屓W�r6�����]��Z���	@�-�c��r�<�xAȲ�s�b��^�OC�G#���h��U/<�`$ �C�0��N:�r?���u�`��i늻'��rȸ�
ӻ@�x�"F�n�1�s� 7N�7��t��U2ֳ�4D�!�e�~T
�PJ7��"�=������p�#��=�ս^6mC��=�P����y�MV��<w-�f�X��� ���?�6�0����\��h��-��Y"/2`J^�KRc��yc �d�=��T����*D��'�Z�#fU�Q*����[���me>�*L;�SYN]��"�Q�S�nNՁ�^��d�HzlPV��|�������?p?��อ�3D��8jɨ��/��ݡ��`۪�9���3:�:�ϵ��4=�1�Q5xP��Z2o�̒,��?�A������5���~۱:i�A�Xn�`t�پ]:�R���7_65Ӑ#����JAO;�V���JL���<�S�6��%I�W�3a��m�ϖ�*L�.r1INy����G㿵��y��ͻ�����'`V׀
���_���HU{�5Y��o񎁑�H���_e��!Q��C�z�2"I� d��2��
�.��5Ne�.��~����ވynZ��wۤ�Yd�|�>�\�U
~iK���<?��d| �A�`Ě��
��ɽZ��y���y$.�=2E��:ˍ�7N��&_ͬ���C�G�G��a�}���Iu����Y��2[h`]�i���v+����w�
��Mr���;�
;s�cy<?��w���*�H<������m%��f� �/	����aYM���L�ԙ6�f������lq�����K����<��`���Wߗ����Y+���V�?A�V<L�:5'~4е�2<���m�}?Y�I}�p�X�"�dG�f���藛2_J�e�!��Wb�@F�9���U�b�lweOP��|$��Ʒ��@�����)$W�6�����e���̍���-�Fn�Ts�À8*��5"G�9��LľD�-�{�)"��ѭ��ע��l[0��},�=�Vw0}Ne�<&�e��[u�+�%M~q ���7#lϡ��o�U�m:��A��#����$���+�N�P��*h���V`���CM��zS#��Ε��
��\�e��(
Ш����7��7D�]� ��b�:�q�����9/��2���T��t�Ȫ����p+����8�ޏ�O�#����=��n�>P��V�)Uﾈ>��S?Gْ���$�u���D\�7]'v�%���x� ۂ���7%@/z��2Ԓ�=%5c��qP=����G��P�|Fu����|����H�L`��L�f���tv;�b^��߮������� ���6�A�['-���'F�~���G�й7M`Kv�P �E2O0��А��b���#��b��t�SC�r�qB!B&����.��$��1��[Z޼�I����$��%�T�'}��^�Ƹ��<+�99ML�����c\���w?��m��a�JE7�?��ġ�C�v�Q�0�5��D�I��ZMȞQ*�-����z��(�`6Pc?v��	橳���c�.�gI>�7�dעD@��t��u�`�rI,\�$yo(��)/��|��������=!)ǎ±Gj�U�Z�f�A�=�(2a��V���9���1����
6M�b��_��w��6�7ij�n8pSa�'��k�ç��W���)I��rs��A��ȶX*�8g�6��!a�p� ����GU��SM��44{D%U��N�f���VW�}����wkD��F6�:\b+5�~�-?��"��Q=`�-YQ>�T��lӮ-w�\����+��M�%�*�g��e�0����$%L�o�v����ZN�AM�p�4�3�~�}���.0�����M=�٪����|� 7p�Q��� ���R��w�';���,L/�`e�I����cr�U�~6zq��׾��Wp]+����F������ƃ�,(�Eq�ZZ �#��\�L���*�'�z ���*�bzj�.�sO_lAޮc�AV���~L���l�[�z\�	�-xAa�n��b�-6k*V�}�\֓�����΋w�kX�� �O�<p�<�vw����z�fP��]2��EA���ev���њ�JA�����!t�0���E D����lz*�߹D�]�������ZCB��1��?���Mn�� ඁH�p�XN�����I�#h�1�.L��#�������'9�w������:��X�/���4=����ff� |I;"0�v��cؐ|��e�7�P|�W��|�a�a�)Jo�L�^9R���O �S�%�( � ������'�$��8��|#�,e����ou�G0T��?�	����1�&P;���RW�WG&&x�%x8�ui��ɨ$I�;gPA�Ti���M�̫�-�����m_�-�6�/�L�_�wnjDYS���4�{�I+�"+���Ă�gL�B�F�5�e��ٕ?�����:$��q��X��q$yh�b��2&n�ȶ�]朙25+�"��Ձ��M|�M����/���$�z9O^y�n���GH{�d��m(,��6n�ٞL�R1t#����h����_zL��NW~�:'���m�Ir���� �E(D3my֥�j[�g"���$m��7�'P�Q9ǎN��>-��:�ɢp|��:o`�j�L��/Y����,�9e>Su1̇0[�k�6�h�p�:�0��6kl�;f��p���=8�Q��y ���3߯ 'R���������ai0��>�!1i�c�U5�-p�cU�{��ħ="��B��o�@BK�AK0��pj�����ٕ5Ťf��IB�Gw�9���4�9���*���q�\�0|��äj�Yw`�[i�@��i&ҿ"v8 �j������׫Dd���r�NCh��Y�+R\�P�-X��W3V��L	Iܐ-�s*���oy\c%�Ag}��?L����g��zw�����Cr(���˗�|�Q�j���j00a���P������z ͩ�5ժY���\)2Yp�z� ��S�[z7�C7'��.�E�q���M)��:s$��=�Ҽc�'8i��M_1�02	�^q��a��������!aq�by3z��Rq�T�_��o�K��lO�|�@��Y�
�~�"K	mcڊ6���UF����o:��9���Yz��VE�{e��?��^�Sr�+{�	9j!���
c��=:g�aN�q�����.�Z����P7�����$�P�� ���e3G��� �A�G�A���d��^�9��������
0\�^%eG�������l,��l��~��`�V*Q�Fo��TJ5���M�93��W�Am�#	$�U�t��5@�J�o٩�EeM,���,�6� �d(R���+�'%��`����O;qո��v�S*��)�?���S��ܮӤ�%�w��ʂ�i��+~���Zh���Q˭J�?�l|��⎆B\F�������Њ��	hg�P�b	�'Q�lX]�����I��{�w���k�}�_�A+3Q̌?�/����%�	.N��C�746��4��6��h���MNW��O9��R����Aw�W܃��1����D�]�`�*���m�(�D�:h&l�/ڗ��=s�{f�����W�Q�>� <����r�l���/OR��p��E������#��o��(��q�	��[~���/=̓�����R�=C������`w���Ӯ>��?�޺�H�nj�=\81~��wɖ+Lf���+c�)P	|X�e���n�ˆ8�jF��U�I�{?��p���ULHzчeR�Y2���pL.DB&������|x%�jE�|�8��R�m!st.K���?��J$gMD�|�~6�M��+}?[���Id�p��b9%E�p����"���e ���2������P�񘧿W4��u�Z-^?��^�;iq�&��� �79&T���^�k�~�+�e~��g��������{�=뗊#��ҚǶK'���Bv_�t�G�ڇ���L9����_�b����l�$�7��Ճ4"����ŏj�r!&�Ƙ�.)Se�}��v�z��KG����7J}��pԞ�O\>4�9u?�_�h��e:�Z�_%��g��p��3��j82>��^��l�d[>Y?4Qۥ��q�U)��e�Spx��)҆�	��-{d������BS�����a�t���Ȩ������mͷd7���>Q܂�-���Ud��!��}��_w�\Ȧyim2q������c���lYMl��^�)9�]��[��UBt#���F_����϶O�~��8��X2`\f;�<H�F-��N�@���j�eLw�E�,���JG��-�(\�7U\#�5�h�Ű������:�S��/́�h��S�L���Ys�����P�XʭA���w�5(���L��VEX*:i~��HK�#_0@��zf��lB���¹�Y��䅊q���=ֵ���m�у��j��>Jnۅ ����]x��8���k��&0V#�}�6�y��w�]��[��W�����N �L��̯B��.D���tFW�l������"�kN��-��#�����}o�k�D�a(:]�I� �t[M/6}�b��}��� �w�5{�����{يi�>\?m�4Cu�$�}(�	���5�9W�~6f_���&���
�y��#��J��:3\,��bە]�0���7KfCvq��8���9q�U��G0��i�r�Mi�b�d"Th��������hn��&� ��D�v�Oz��3O@�����Mv����p�(����T�f��D���A��k<���3���P�(^*_E�_�ؾb{�g��k��h�����m	8`�"DQ�)闠�̋����U�h��2�<;���L�\��b	�Iq�/$#g��p�l�Y�D�=��k��m=
g�����QO|��o�B��l�K��c�'�V�D!��t&���_�A_�l?`�Kýo俊��i�&4\�吃��ۀ���g�@n3� �Pq2�5fa�/rܪ�g�������7o�d#����%K�SM����&��O���e�;�b�H�
��R��!#rV`��3��ؙ�ⷃ���ʣR?��ޤ7��q����
�ny0�`C1�iZTu#Xh�i.0�ƹd�ýy%�qE��[�k�`<@�o���{ߺ.l�(m.���.�F�s�ۡ�7�垞�	����(��X�#Մ6��b��&ݭ���	������=���'��嘠�!�}�;���9�B����,蟳C;ow��.�g��Mыǆ;P�_s�����Vy�|�z����s	�_�j�?k	���hV���z���O�k/�A܅R���#`�0��
n��*e�� $F��L�#�� �������u6��t"�(�6�G�5("��t�C[��T�����"6�s�g�|��4��(��*�<6ZI�}��$���C� +����lw1�d�BcR������M�P5�.�^�#�>4	�)�2�nF�!_�J��-��j�ܻu��QŴm�����E�g���|���/��s��tW�]tJ�<Q�z6w��9����6υ�*�f_�"�c	��R���8��w����U}���1�[6�g���β3	f���g��N�뽑��I�����.��y��x#u�Z¡{������0]q�_\9��Z����M<�e�e���HG*1�����i����v�l$-��T��7}�P<:����e2B�Bĳ ��y.����ϔ�����,�� ��ϸ�у~Ay�]4kM�3U]��Y����Ϻ8���" �R<Ԩ�~���ڐ�=FA)�u}lVF2Z%�`\����H~�c�fQ�a�����I1�ڽF���c
|�<�9&2��EEܝ�
/]�O�%�(<�����/��j<υ�Z���"�n�<��47���zX�+^ ����̯���c+y��Oوq�Ń���E�m�:���my�˰u��aα�t�H6{�?�ڷ��ΐ�iL&{ƭ�a\Uʃ4������
-��E����pKg�����3���8C[v���\���ԬjB���>۟�S��&Q��ז�V��:EQ���]X&z�`}t���K_/�7�y"����si���0w� /�:G��!����taEݍ�\�~y�Nw<
K	Bbx���M_�- �A��wg���� ·�CWf���A�O�_���� g��b�!��T;�M~�8�d�"E��Xh5��O�6�&�6������hD��px0�'�ٚw(��sZ�TvIoa��J��7���5�}ƤeC��^OZ˧���D�9V&�zd������Nl��6�L�b p��К�(3
�d�,��c��	�q���/^7�̕�9����uB)?R��/�``zo�$��1��'-��{v��p�ר���o����ɯ��{]�˒���U�Γ
\ �̷�A�A'ި��$��<��'�n��0n�������ڲ�;i��,��_����uv#�`�,�H�&�,?ޓ�D��S���lq��gW�����{ݖ�������j��k7���� ��ʙ%��DN�:/_<�N<�U��[�\�c
�j�W�-� ����S��'�$���?�*�B��O�v�&��.;OG_?���Z�6���'��{>7W�
(���b>%�2�����ژp�����J.��f�v�b؇��]K�EV�Y�,�ۭ�-�dlJ�l/�"��ï*F���9Y��:�\��vi�`�ܔ%Hi����7D�J�X��g��I�%�ĭ���A��%t�ǀ�5�<���om(*VDX4�ڟM�ݐp�߂4�ST��)�=�q�̰���� y�Q�[f��@�E�O�^�j;(NO����r�,D��_��m{���FQ���zy"���1ZczH������i��������qB޾x�R]p�DL�
��Q��$�� . ����=�D���Fe�s�G6�An���d3�ж݄���[u�Α�T'��a�Z^��=~b���p���Iވ��5!�0S�c���3� �{�EJ4�m��	&/���X	��h��8��8�l�G���`+�s�2��ݯ*�	��"3��eM�f��?�S�YXmT��k�龼�)�Q��`�>��F�F�
��<w��-<�B�A��7���{ �W�Y��h1�2?�q�5�WK���?�FU����1R�5��?lb�/*ZeT0H�oM�)�~o������<���N�J�Kf�_��𐐸3��}lb�`)��&�7]#�*��fn�o��GJ+�u�	�շ`L�8Yd��,�Z�d}�C,��i�-?hY�DU�� ��������� 5
6�N,��Z�UutpO[d����z��x�.L��V�m1_�o���f�E�T�\�j����j��_9�� �*[��y����Bnm|���"bU�*6���?�Sо"i~Wl��o\Ӌ����LP�¬ڵ�j��6��V��v%�H�8A�����#��^�]��%u9��E"��3��p��̎�-��0�O2������Ϗ�����3���a��o�LJ�օ�������(	�`��,�I�����Lw�IZ�4C�u�u�,H!�ӂ�nBOW�2�Sԓ�zJ�f�)���{Tu�O!b~���v�����ع�)Na��J�)�3��n�]9�L���0R�s=I@:O����%�w��;^�
)�~8-QݿQ�}�?�<��~rBdC�Y�ws(��Sz�
 tT�\ݑߗ�P�3�6B���*�Q�\���܎�NI���ۙC6�q&��P���f��/�m	N(�\"=-���#Fi�V��0��ꦇm�D��:T7��̢{O)�2	W��/�5T��_ͦ�����ԩ�m�M;�c���+��^k	د��r©�eg�2ٌ��y��oa�)�vI��nԋ/8�U6jƩR:�٠�, ��%��ĺ�j�J����Ο%��y5�*c�|$G��{�=�44�]�z���gf���q�N��niEEx�6�+�v�3�/U��ϑpG�L۹Ǜ��[l���J�-�y�����Z���v
6�Vb���kc�!�`q��5��~3#y�&�^��/Y���q�E�9��Z���i�i��c:���:=��2���N�hd�;7�e���L��8����j�u��Ӈ��p4��>^͂�	iо����}�i��7%�}�>	��-�	��kի���KnaDU����E��V�.�۬Ses�V�Vxs�ѡ��j��<E�j|�R�J>�D�*'�[c�7k(3Y95��(>���'�{��KK��~ͩ���:b=�1Yl�c�����nT]�t�w�j�!�P���3ib��--F(�Ķ��z��AE|x�fb�_��-�Bp?2��7CH�� �wڻ��hz9R�% �]��L�� ���-��v�+�OM�(9�[=�]r�����[����XCc��=��Q��2�ꩉ����왫��:��[���I���KI���A�x/C^�
!J�<���;͝q=�{Εּ�jf�E�Ōi�n#T��{�4,���8�5��(�L*XA#�j3��^\�ű�Ǖ&boq�u[l���|���L��z2�]�p��Y�������|zC�ZL����nk��)aZ����0hz)��	J�볟j���IJ=�^(�/.9H�.J&		�	����b�Ct�ܙ`!Ds�1�Z��ٴV�֌4qt ��nڧp����7�C���k|e���ҳ��m�$��>E*���i���j�PY!S�)��І��pf-��1Ă��8_���QXx�fGU, 7HЫ�И�R�`WwK�����@�a�����q�f8�v{�准�5w|�	?[��t�ǵ�)@�u��a�{�lErK�� �l7,��3&gF&���J��HE�B�z���hfo9fZ������uӅ�h,-�@�}�����*\TO̤�M�9��$��vX3m��|�p��x�R-��A�ca@u�z	�$��ƮM�ZBH�i=l�E|�r�o;�}���	�~�(d[:��/}Ooz�:���Z|�g��§j���S�+��������F�km-�rzQ�Pw��C_� ���}�)_���M[�G�O�v���7qq':�����hL���#�:ː:)�=-��(��s?	[l��~.�'^�\�	3�V���D���������s��8E��˘/�)�v#.ׯ�I'i��4l�$oG0o=8��掂3Vgi��D���f��{�b�I*�N�����]�S��"�#�{�}T+��RwHtՏ��V�U֥�1�)I{���<Df�J�-w
|��F�ɓ��c��p4� )�05籌��Ŷ����g�����n���H���^6K20�z�R��z<C��E@���Cbi��ܙmo��~ί!꧔�1yyuhR���K���.q���;�H��pr�����Dn[�:�[U��k��i��L�����ǟ�G�Eϭ���[��l�L��u93I��\?�����g�!m� �`�p�]�W?	v�����J�Pi����,ݫ��>�:����dd�.4;cX�e?`�S-ug�,NaZ�q]*m�Ǿ�(��b`�*Z.�Y0��˂���w`=�Y��Y~����r�;�vI�P��9��XqV-���9.�:��uvX0���K�NL=��]iJ5��y#�}����T85�P��
�2��7���U�m�ߋ��H`ܸ�J�;��2�>0Z��N�K�p��r������g���}��*�	�3	�;�Ae�]�\jN�jY$�ŌUJ7YP�t�������ಮ�R|��a�I�D�%V
tB��w��K�����.��ш����FY�*��5��v�_����d�ް�*�|�b�����	�3;��a��&�I	sR@a]�J��?����W?���}Y��բ����ID��N�s�mzn����$hT�R��p�|�׭'H}�i�0��p�1>��N �Kmڗ�xX�{�N|){�Гh1���>,�6�0�=�|�p�����.�ԗ��T�ĻN��Z4O�V�?-:$͵�Y<kx�����L{wD�����ͺ��) �L}�.
T����`�ne�T�p5��-����V���md�{6M{W5��u��:���ZB��t`�t��J�?� �"cC�"��6���ɹ�R���a�����Vb���X� 5|6��ӑc3�~��s��gr�M�ݳ5��;�3One�\�D����[^�Y��U<?4�����v|�Pla���<��3�h}�}sC}��A@IJ�C��^֑V~h2����Q�V@�	�{�J9��??�d��rJbz$)�)����V�<)ѡ�6o*
�x/�a�x�i�1����U�$�r��ۍk�=,yFV#�\���fτ�F�u��̹P�:������ _LI&5S����?-�T~�[��s#t�C�>�O���ǌ�τ~�t3q����5�%ȁ��ج�2��W�f p���J�R��.lƂл�����S��^��5��#��Pq�
�{�˸]�Fq�����=�:�\e�X7���T%x������>v����"�
8�)�9� �D��~����=M��D�E�C�Y�vQT���fy��-�D����V;mґ���F*[5�&�D#�������@ �#צ0\�����*�u��FEcY��A���.�|�w��9�Q#������V�xnpu}�@Zeqj�]>��e�����)�R覯��ȣ-��{���~c�'�B�rT��SW��H�s:=>��^�I�wbL�R��!NoQ������B�)|�_�jE�ֹm�>qVٜƌY�S��3��3�v+z��5�5?���n�J�n���iO��v����0e!�ە>�7V:[W��|��ń�cs��e��Ci^�Ŷ�
_��j��
nq�%�d�׎�_���[����	�7L���^�j�>']%�<��R~�J��w+�+���״,�
a�To�sb���~�d>Q W6H��j�HJD��2 o�z���"8�a�ri5������!A���mz�9"%�yY��|]�j��ݩ�ޤ��sq���n��K�,9��+*��K�9b��Y�r�	��#R��N![��]@���ˮ�DǶ��! ~pMY���f��p7�to��n���_�B&���73����8�o�4���ޕ��p����P^���Q9�~�����2rL<��.Dߘ/-��)^�a��V�~�@����6�u�t���T-��{�cg]�:�F�U3��n����+�D�<G��D��y��[VS=�m3�"o5{�3�ە� ��)��䄢��΅XC8�T��C�9��%� m$�|�D]�#�!:�")��y��%��y���ފ�k'��?2k���q�'t�e��TX������Ȃ"����f��8%F��٧��"�Q$�V�-_H���1Q�X��ss�ғ-v&�E��$+nt�*�q���A�N�:��V�K�=�Us2:ϕLE�QE�����;�Uϋ���Z��P�h����&���.�P1J� ���*{{*�Kk�e�;b�;*U��Kg䖑Gv	�cLi{����Lwc �6�{D�c%R>r����ޥPP��~?bs�(��<�?���7��-ZcX����5�~��u��k�d�<FfYR��`*#Ө�jW��	�"'@�6 d��i�f��S	MI��΃f%u��b�e5l{@-�x�����i�Z�:�� �2��yA�G�/=�X�kM�B����ODS*w=�<s�?Uءb��)f�>0��K)�!���f&>�!�!�)�/8�5]�����ѵO����bU|;�.3-�.B��Iz��O��ML�O�o-�<��>�S'�#߅�\�9t����z	Q��F >�^h����' |JJ��lw^����kݘ�Y�z��*$*�l�m��������.rN���p�����;�ڭ|�O��~Уr �d����Sn��I}';G~|�[��m�=��ǟ�=tB�N�G���|� ���
 2xzy�D|�3��x��p]�/|���E�'M.�����G���@�^��}�yR(�"��8�ɪ�z�/P��t�s��|��2N�e���łE�PfU��R���t���2���M�&*��gH	n�}"v��+a����=�t��x$��j�$��?�y�K��9E�ٜ�{4�T�FW^Sm|���w��_������	#�b������cN�% �] ����?F� p�C��аb9�/��⼧�rG]W(X�dk����,��f3v݊B�Ef&��Ό��\���<�b�v�f�l�&ua_�w|R��b��f|)��GٺPۄ5G���.�X�{Ic�f�,�C%��f����>�9��#4s⿄��/u��"���w����,	���ik�d���rB_���_�T/3ك��_�׳��?�iN��s}��<��uq+���tB�q R����X�OP_9:7@2����&�+䀀�]�!<��a"�]�T��Ӵ��/Q[���[;��p�Ymz����|s���p������C�0�#U�v�Sɯ��`�p-14��!֓�Gp3b����6��ٞ+�|��J�0����}-`Ë;*b�{�bB��3f��[��]K�(����3����>����h���7(0�����-�kd��~�+��>9�֝����w���G9��'p�_2$�ٓ��^�V�߮FiTD����&��rf6�"y�$1U��u��h���j:�����������
����&�����0*�P+�� K	���S��~n�F�1�C�c��'�llCH�@�h�bބ|�n<:.�@P�)+��	o�n����`x���ޱ�͓����I��Rn�)_9rǨ�����l*d��w�����H��]t�[�#�lP;B %�_�9����#�5�=�5?xF(��4i�a��P7�x��L-�őƙ�zJjM�՗4�=����ũ�a�@�n�*���(+�'k���h�� ��*Xd7�4ʨ;�3�KԳ#���n�
2�D!��<�,h�mP��Q�}K?nCc[n�]�Vrď����������H�}E�<� ����.�EYpe���}����"ɔ:5 v5�\��Bi:T7�=bC��+�悝�4\��!�I��fе� 8v�-Dt���X�9ƥ�ˇ�&z�6*g�W6C#nJ��KW|Y|��,k�,5�f1����Z��oAf��{�1A�j�U"d���{�vU��M���E�M��p���~_�ma	X�bf{\�&��V��yȮ������ #ɝ�-�����3�6�8Z8H��ϲ�6Y�����1��Ec������i��g��|n1�����p	�pES�%�كi����4
�q��}��P�KD�Jg��mN���(˫���4����*�i�ڕ�1̀bm�|ُ��[K>�y�,s��et�;�ܘ��I�)֞:�␋������n�k��VJ�y��O/��kJ4�%�?���Ù��P�4E��p~ �гLED��L|H��7h#�7�?7�M>��q�����Q ��ٕjT��v{�u<�S�y��6�*�^hDT-M��/��⬡��F-7�ƈj�/ÿ�|�=7J/����ͻ}fi(*��c�<,F�i�� �J�l�C.�+a���#B�����#��� i����z��Rʽ7�V"��ݿ��pLD #H�Ri�S`C��U���fUe�6��������:B��k�ǥ
��U�0/*�_~܈~�������DZE�E|~��;VT���L`�����.����6 &�c��S~BE��[5Nc�b�֜+^�s�+��p��]3t���'��D��8G�������h�P��ب��@�x��g����p|E����a�P�\�Ջ�&	�/{� ��N��^���RE�� *>�l�7䢥�Ճ同�Kg7�"n;aDO%��/�I���S�}"q��\f���%��^���Q1���hIF{f�'9�[�6����s�h��iY��s�Se���E�K�Զ���MB����E9)ǋ	3>�N�͊�C;0MU�����VmW�����%7��c�����]p'^��ld�
̘���m!s��c�iт����B�e�*zP��I){g�N$oc�(�pƜc�@�ݩc�;��ZxO�R��b���X��o��C &��Kc	繛��h��V�T (:=4[T�
���'��/Y$2w��b6E��i�bg��9��4���୍s��v��](C;h�U.�v����2ԫ���i����j�1������U�p/��m+n��v^���(�Y�L������cH����L9��+�h�	���$��KG#�����["23F����0�G���b*�I�T�������f�x_X9אtL1��>|�6���#r�`�:�p�1�QK�o5�t�*He�k�s���Ư���]��^��� @��}?	�I���$��Ҧ��4��Dp%u#V��J<�&�{B��>7j�g�7��8J�p�p>{��5>�E��K #͉�;���#�gV���̀d��g�x:vt��͍3�W*�%=:����ȕ_���_ߩ ���b�>�$@f
� ��4~GAi���ݩg<6�b�OA�ߪ��Ɣ����=t�T#�l��X/�5[�Ϳ�vc?͑��q6ďP{B�F}��ӹ�-L�����t9���.o+�U,��X�A>!���"���<���D�g0���q�a�R�:.�S�0�1�]�ί67�}�������L��ޛ"�)�o {�@C.,r)�}͟�@�:���([�:�V��k��O��$P_(��}$���>���7=�ʝmu��/�]76$ ��5�K�ξ�ͅ�(:_fb����,!���f�|uTɿ�I�=�h����k���Q7cJ>P�@���$�$ԟ�]�m�w�\ɓ}F"��L�ԥ�Ȃ�]xxc�s����xפ�R Y�MrݓM{��G���vs�%� �ˣ0"*X���i�~��`©9��J��{jn�g맘�8)���YS̡`�6�[���o������ђ��7^��FM'����M�Ȁ�b<!��@�}G;E�ҜD��!b����~X��Wsg�R����O��7,3m��r|l.mA���K�D�zM�l�DfaC`ހ,� ����o?�aF�F��r���n��7�O8�#�˦��v���j��u@8s"��P�J�!���Z<G���aub4y4&��o���I�1o)%���r���,Ub|h}��V���xᴼ���]9)�H}M�\�=}+����i=�`m��A�m��5Hx�ФC���>��r�
o����������*�`��_�V������7	�Jۇ�ံ|�W1-)oV��(9	�����&!�Ll�p7SkLP�-+�KV��U�	����P/9���<��X�d���;����m��#"�]o�ܡklw����~���z�������(�0[�6n��\hm5n;�"7��ک���!\��`	���t�Q�p�Q�=�����j;(��-�+b��J�\)O��6�>��Gv�X�f6+��"���~"������K�b�L�U�*��q���z�6f-�eb���V�4�Σ��+���ܒ��^��^��*i���P��n����E���Z��c��y�}�v�YZ�5��4����vH��C�.�����)ZH@�{�G��(��ֳ�B���UA��RB�e�ށό��7�s�Zv�l_�?#H����Yp�L��\.EUc�PP�������i3��9�1AW���S?%����h�P���.*��,�~5Xf4�5���D U��D/�>���S
a�>�1x��_��X=��1��������n�|͞7��+����A<��ݤZ�i���_Ӧ�Bt���-���Yal�l��1l7,�i��2f!�i��������z��{Z=:����1�;%|��M;�=�Ӈ��T��8��g�60ZiA8G�|��*�r�4oXX=���g}5M�PT�{��WhEB�4j�o3�SSh����aR~��Q����_c��N�Cmm�-��<�*
��$	_��^N�Be�ˊ	"]m��}/*��%ײ����'M	jA2ggb��4YSԢ�_/�ᶪ�%�ǻ�t���w#�h��� �B~�����u�\��W4Oe?L�� ���\3��#�����j��A �_8n�2f�H��٫xH!g\�g|gX���ܹ}��q���G��=�B���((ˑ|B�՛������`���.��Z��"/�CXe�����dױf�ʔ��d����?�����u6�{�KY�M�&�%��j�I��������:�� ��'1)+������OS�Ʀaf��'��8�%�i�����J|6���k�L�a,~�og�m/��E�_��S���xiV[���f�����%b�^nT��}��l�E�d���5.Gq�h��K8��b����iW��� �G(ʫ�$�4GOM���d���t���L������T����=�2�x�F��v��5���s����*V�o$�?�h�3c� �P�np��y0gBS������W�d��P�b�(��~��I�w
2���$hN���%�|��U�@���MD�Z9��p��s@�nKWO2(}r �ha�"Ku��$�SS�v��(�&z�S*O[ZE��ϧ�t������xxF儣�3�]W�T���K,Z�$]}��!���G�RR�8Z�w]I����m8ҷS�3�	��y���&xb�Us�h�I�le9\���O�,�s�f�y(N���o&G�����B	������Zzd�q�ޱ'�Vc�z�pB��?���C_�;�V�$#f��́Z޳J��)t�\�&�Ø�r����7�b^�:zo�۬� ���M��պE��a�]�>��]P��Kx,��=�v��V�pYN�x{p ��[���(�t�|!��CK^�+��j��Sk0�k��g?�d�F�>������C����-�৊p�ڱ���/�0��J@]R>��rDy�0�Yv�kϩ��jR�,�5��8e�tl&���F���0��J��HCZ������6�ol�J�� ��a���or"���A����e��ݭ�5����/M��ۇ>7�ZW�&`�b,�f�p�������.Cx�׍�:�ސ9�jt��ෝ�~M�>������s�'��pƬ�ں��#4�w�9H�z;W��P��|L'j������v �QN�]��?i���3�[Ŕ���R��L�ڲ��w�{�&D�߅�Y1n�c�Ԯ�HHv��S�W}���%	�8�t�O����ݨ����Ͼ�Wm�?~΁��`T��*�Eՠ,�o�Z���� W?�h�����9���^#k��[�f��{�v'�[�����)+�8�`,�ж3�}��X�8fN� r��2�Y�rK�p;��` wp��P�$�|�E�r�&;ڣUE/tIZ浫��������aKGA|φ jLu��j��H�F�$I�����Mq�w����v�}_�<,�	Ղ!N����N/���IEQ�a[���HiՔ|U8e�Ym�7/���3��Rpԁ����[�*�4�׻�����k����@t����ܱN=}��p&��	�"��?����}D��\�Ɵ���]����_�n�,v߮3T�D6,��:h��������R�2@ʻYv�3 �}���Xm��&�{��xP����3{I{U�z��la��'�G6:��G���O�[R�k�8u�� W��?g��I��]T�t�j.� ��J!"h���*/бB��Mچ6��A��Ӻ >3�Z�.���,��6MaȺ�ܿ∗w~�6��D�%3�=�mk��_����7�F�r����ql����΢���jL���0�$ep�7t�c	H�+cish�(-*��bg^+g��`��Omz459z�X	W1���m32w���&dE�/�+�	Lw���i���w�y��1�͛Kv)��}Y�]�J� (�>�d�y���CϽ �l�"Q���'���@�Bf5|�W��@j)��+��ִz�<���Oɮ��j#�0�<C|c*é��'7j��#�$�c`{��qt��}ElxQ�6��9ρ_Qck��;��7-߀�y�=F����t��:s�|=i��&��]R�6_��%�V�%R�6�jS�� �O��ek�-�R�6�햔L!�Enc�,t�=�G�nSԍ�Ϡb�g���H�p��"���D��v����� J>�8�/��U�T/Mٓ�[GUc*�Y�����D�4~��-L�%l��f���[sd`���H;%���sm���쑽�R��Aڗ�����:$�d��Q�x!���'����e̓V���Z�
��#�6U>�����8�7.�1�"B�n�W8����f(��;�۱hOg����qJ��!N�S4��!2��#[1Jp�Fz�^V,���!����3�mN`"�;�y>��Y����?��[/��qp}�m*�"!�Q&�ՈZ�^zV袜}�·����C�m���MVZ�GIH���}$ܭ���'�9�2�d��H�/�]>��$G�_VPP=q�c9P�z�ƴi�Ψz�7�E"j��'L^��_(��B�����������}.�$���Ĝ���5@O)��_��vޤ�<��4�>�����s�z>@�C���_�a�n0��Rhێq����Cp��9�DBi��Na����DyS �vi]�5�g�n�x�����.��#"���}ߤ�A��.<�w1ř�#��;?w>�y{����_Ð�iNG����¹+�Й�=������;	�.�7�����,]>�D=���=!︝�� ��#L���ήWkťg�yi㽋����=Gv�Q�j�F�:�M�/�(�b�^�S��]��q��FQA}�oyZ�#�ʮ/!��I��tQ�7���>���:��ػ�:��]�4�QL�R�k���qK2��lcg��Ek�C�Ą��t�ԣ��ij�@�!C��6A���������T�)�5a
�B�O����_^��t�8�szÍ2G0=��fѠ�v�;��.Qf3��@���v������8�P���5j-�Iv^�&#�"��_�#�]o�D�Z_��LJ�]K�����Hv��.�s�%��}R8@�vt�g���^?�x�ʌ�k�a{dos3,��(����r�Y�v�;��Y
��3�J����7V	^��Lу��rxL=O[9��^PDc��J@�-
��,y��x��e���YM?���^�^�Dq��)�Ƒc�]k��D��3/�3�poN����>��n�I�%���Z���1��8W\�&�]�*Pm�)9ꊇ�-ɘ�f��[i�z|�r��}�3(�C�[|��h�{�/^��Ռ�֨Z�>J/���i4���eB<'O�>�vJu��œk� �GCEU��ya>�l�u��U��'�JN��(���h^���Eu�W|�7�dᝤY�oxТ�;?X��ke"�B��%Y��rh��CEUl~��1��������؆fy���H��N$��y)��}bcpø-utwj��]��µ �z�<�/^F`r��0+]c�m�n����T07]k�j���Ø���hx��;moR1=���	���kN���s-���5I���R��h*�w�pf/K�*���⯡�Ϟ�!�O�:�3O���?���E��i�r��'m�V�WSSDF�C2��5�좐�y��-��Ci`�~Z�at{(�pX_�̥���d�6�6Ya�ŊT�`�V��G|�旀�J��Lt''I9� ab�16��2�S��wqD 	l`Qo7F%~!Y�3A�atW���p�1�)͹*�՝J��a�"<֒��Qgħ"{_,72� ��<����V1v�\0�Cy�
DPE\�s
K���^)��LÓ��HF5+�I,2-����׿�]耍�d���+�n���>�VN�s"V��Ho������yegb�<A�q�|�h�h�?	��WqY��xI6�'\��o��p�f�+ &��sϒ�����z�Mq3�fz��>$�9��!�z,E�r�o�i�ai�q����E.�tr�A��#�T�d��}T�#�pF��k'S�R`�ʡ��Wa����"�_CU�'�'`�=.��O��I{�@��ꀇ^G�S�Sp�����ƪR�+�}A3�J�,}0�V��gùq�I;�H�m�%�4q�˹Vj�ޒqZ���+I\b*&tfDsqv!�ju�k��e��nՇ �tΖK�EFm�c�0��t)�n�G9ڢY����?�����Řc��'�t���R3+7�۽�4���&�jP杏�˖}�%QWt�|�h�м��PB)�����o�>ƜF �� ��{�ufI��`��*�*)��x#��]V<d��'��툇W���
�;�U"e����*�u$Mx�7���s|�nt���N�`�h��+R&Z%p��}.Lg�^Z�Of2���$��bK�8SHb�bV\���A�Z5]r���v*�6Je��;���Cv`�������������Ҍ�`���*�0|}��?�������(�^��+Y�H�x�/`��r=�؈{�֨�ٷ� ����Q�}+힠�)�=�0	Y���*>A�;am�L;7
��LG@[$��rT� 7��cD���W]�/ۆ�y|
^GUv��J�<J�� ��h��������D,��m�.)��ԇ�򠹠�D��=��^�5�X(%�,ԫC���֏�$���e��N���&&_�9'̳�$��an3��ו� +%`�cj�t׿4q��p�.: ?����<`���D�n���3B�y3�oEmV����3>�x>�G �O
����U-_�õ�j�K��ojI��ٯ0@Ӕ2$u89f?,���r0D�v~����G)�0��^uSA'��ٓ�3�F~�Mr�@� ���ՅOLk~u4~���s�6mXa6k�a��[~P��Ta�i��(�SbPr��
!�ScU|q�����O'�s;�F�A���#�gxl5�Eǣ�D��{��`w�Zl��J��4~l?���0���O���ɏ�hj�7����u��4����9����_,֠����%�-��rW5�>D���0�Q��]�G]]&�/�!�-"ݔd6K���2��ͱ���W�lO�Ls�V7E�f�p�U�\���re�H��8f;�cL��Fi)	����R�kQ�3��=��2��#�S�(�R�_��@��A�^�kv���j���OE�L\���!Oې��.r�v��c;�]�V�j�v��{��Y�x":�ss��+TaA�d�2�$}����.�_��N񿼷F�Z�5�w����b�u��P�8E ��@���JS�øA)�_���{�)��:��	b^7��RHeA��D7f��(+�����W�-ç1I�RC�����
<u�®s�9*؟�y���)����<��w�U�o�@�>�xZ���#��Ѥ�9�� \�@g�|,9b�,�|?��k�*�(ym<g���A�����BS��N�?/b�{
��A<'}��o|�	x�\�h���v�����6��ߒ)"���\�C�s8E�>�	D��If�����ݠ����R7�o�u��՗���x�l��b� ރ
0��B{߾UY˵��"��˝�H���*��{���cJ4��3�h]ӹ�����R����njʵՓk�z3b���I)�F����4B��n�:��ef>'B���!,r�1�.ed`6i%��T��s����`�,HQ�����A(6����K�m:ӂ�����=� ��{�n���W�t�Rf�����jL���@49�^��E�A!���V�P��nE�1�2`o�&������e x�A����y�C|S�KQ����ze�Ă`OEUL&�����:��A�?�JU�|2�V�����K��"p��K��'�$@���Wp�`�M���oLU�fazkd�f8�� O�!������|���<&Y-����������4��=�|��Q]_4����ZSȈm&��o�N�*.B�&�~���f�gi�Ɉ?�OwNs�m}����\hH
.��U2hp)KV<H"^��g,i�����8�D�M�[
EI���fס����[�*��
��Wǧ��6��eI�Ȟ5S�bä�a��.⨎J���L�k_pB6x����Hk$�L�����$G�:��o����.�f#c�?u$�(L�%/���7ٲ���� �~Y�~
y0�a��z�ޏ����k$�RP��B�ݝ�7�*|G�9+���|3�Z�p/04I�iDv�J|r�@@1��-��c3�=9��{��oH�F;�m#�A��g���&��}oR�-��1w�ne�:ϱCp I�H��P��B�VT})�����UAf�5�V̋��0�2��!>0�Z�cG�1��J�֋=
�s�w��;���Yz���
L�4gPR�0k~��f��ğa9��̖RT���*C��Ly֞v������Z�����t���3�דt��#��(RDMU�.y�a}85�۱o��(3i�T������L�`|���:��`�� ���8u�NZ��W�Z:~FD�/2$��J��A�L�E�YzM�Y��6ob�7�#���O��{.�h��
%��ir\�7D�s��-/hX+��A$s�c�o��jN�����X���IE;�(15��C�3G�	�z!�������k�U	�ehK@) ���ܬ��)I�J㽷��MƢ�"���N�3�~�BCN4��V����R{kt�l*����
����}!��xN
١󍾐�S���z����Ÿ�񐃜:zM�`�|��)z�.v+Uo�C$� p�����hқ������05����������n�KzBK�gUF��P&�"�D�)4�B𬁨N	�<�b�J�Mτ�}<���������c郖Q�ǐ�g����/�3�><qu�� ���B�r�Ɯ~�z[�g�����u!��p��>X�ݭ��qVp*K���w!/3�9��YvZ��Ͼ�/<}�m#Rl�1<�%�X��f��j~��	.g1�fJ�}�G�7!\I���X�c�7X(ŏ7d� ��r�Aр�<����>=1�������N�ϻ�d�4'��8��X�Ć�I/�UXD+�I����(��9k�s^X��$��s�AN=�
)�YR^ut[��pW@��Ͱhm�
T65-T��4���kuVӘ���;���;,�9Hc���R�ѾN�w��Q�}۸r�	c.H��j1Ʈ-��)	�k� �d�����D]oB�ʚ`,�^��]�*]���&.�'��w7�,h~�w.�!E��e�����4��T"�<��e�pt_�+w (PW�'_OZ��+�
4C��Lsy�t5~Y�����ʓ���r.�;`�`@� ��b9���=A�S�T���i^��љSP��!��p9De};�^���ϕ!䀶8	uj����xH݊B�`Z9c\ B���z�t[�7�l�i���n9;�e��p,�>o�]�C	�#]��z��b����p- �\�.��8�E�R*7áv��2��m&��L�!����f������Val�d�9�\m
;�k�a�BTNzC+�
 i��v/��oYx�P�}�d��d+C�y��Q`f	�8�;HKugzZ�)��f�����4ԭL%+�UX8�3̢�|T���YZfϒp	��7�Yg����C�.�%������]S�=�Re��Ě(��[e\�=�rM8���2j��[�<����jz��fw`Ԟ1�=$��K�s�6�pܕ销Qb�$��v��!Hg��_F1�2���FoU�RJ^I'IC>g0��k��߫�� n.<\�[88<�ާl���C��x�,�-�W���>�Lv$�I��ɞX����_�$���4D������^���4�x5Ks��"Zޠ�c��!kp���^�T�)�܀{��b }�G��[9����D LU׽�^�VAL�,L�"�sk*�96��G8v��#4G���^>wzzG.�I"�.��0Y�&DO��[?��0MHxNȯ?L�n�WO*���P���)@۠��Ml.�0+�8�=P�=WO��(��@6��3��^DI��߈��e8���hla��N����zZU�o/ǌn�~E����,�8��@kS��U$�����T��V=��@�+Cɢ���{�����=tv
��82q� QnKm��C�9�L]�Q��W~���}иn��4W1G�_ٱE���W^D`��~&E��m�YK��
\
",;9�DE�q��_EW���\__�D3��򁥓}�?�܅an
�F�B����%\��:���8ֺ
�so��󥶉�C���� '�t�ic5���a�����E��NY�	%���p�+�񱽄0��ްH����H����_C"d���!���g>�P�L��A�b<u��ՌN�۵�}�;6�x#z�[/O�Y����n��0��4P�%�3t�k}��m@|t�u��m�_v-�yoJ���*-wTm|�x�;��~���0y'|2h���="�s�/,`r���d��M�ꦕ�fRQ̗��|�o��~ ��t�U ��z�c
��Jd���$�FW�
w���� �G��If�Y6�
$2�F�O3Qv,�d��ڴGbŲ��0�����nD�7�~��}y�@���lV���UU��ça�Rn<ů�1h�����Z;��.�4]�v��CP4�\w�*I�?��Ky���m%��c�0�!����e� ��e�1]o��J&#>	��w,��YiO$���8����U҆r�CkfS�[϶̄.�ywhk��c�m�!%�o�u�fs�C�ޏT3���?YB������.�ҷ�u���/��3ӡ�<vl�Xh�S� ��v�E���!����j��˶w��wB���FJ�3��;���y�ThSTJ��}Q������A8�(��O��o�+(�	߃mS|��m����֜��U���N�\����pT�	ǳ_�}�{:���(��[�Cs8񯯈��,e��-1n�ד �<W@k������ق[�\	�7HAP�����VR��Ӻ�sTKb��/��`C����S"xb?-�[��7Ia�Y�Y�p�������}�ޝOl�WD���)eh`ک���ԉ��f�&'�wL���ݡ��)fga��s�e�y�#���!T�?�I�����k��Z�sl�K�O�B1`�ߠ��!Ⱦ(����~��F�,��G�Ճ\O"\�k���X�����;�ǘ�"�����3����w��Z��e��(]`�6�T�e���y�qe���x/�3v�l��q	9"�7k��� qQ��\mAR�����ںl�����e@+�l�	?����y���~g=l֦5	�	/.��'�D�'a�o��j��F�{^	�����e�tZ0Q!O����L]�F '�W=�
":h�8����c>��&W��\ċX�~a]�|��`�UE[��n�E��r��&��8��^/#u��Wb�ދ�$n�#Z��h�S��5CL�MROx�	L���UL$�c胠�饀�M��d�5��r��=J����c�jϝW�Q�Q\�-ЋYu�;�T�����e�Gk�?�5{?pT�dz(����yE����)�yf���,x_�NA���1됎�j���y��.6�kSHLw_�
��UJZ�V�{�D!�k�"�Ztv\�V)�Jg�ݸ�o��}H��P �q�c��uνc�W���[�h��yQ�Y�/�o��HޡUZ�6nrBP|�f�E����i���������Vü++JH�i��Q]6���_H.�Yi�K���5��&]XH.���&�E[��N��K���0
�e5������ǉ���/�� ���lb�g��-KH��
�b.�F�	|AKc�}4�xE"v0}���,N�<�*�~+�u��S�G��0�/��1�W��M��4��o#<0p"�C((i���P�pi+�y���=�`O`2n�H�.яY%����
>����[t�ZɮS�f;
'�/�m��"QQ
�r�Oy�l4Szw:�r� ����D�aE�޺3AG�TSj���i��ճ��Q&���^?.a��Y�M9�����S8�M�p�|h��<��R�? 0$"�5.������K���D���Ӏ���Cef�7_�P���l*��� �̌��US��/�\�A.ѹ���.�ַ6��{9�6��m����E
I�3L��M:/Ħ?E���P��,�d��_��}�T�d�$�A�������f�KX���Ƶ ����R��]�+�>yd���'�L�딳��.-���
|�t�����h�f�5U�ހ�O<�:!B�s�+�M�7d� �u�
�/ŢwBT����6�w��C�̐JJ�Q���"��Kһ�κo���8z�e�(����q�W(����ܬ�V�X�7#^#��"e�&����~�`��S�!�	z���t>��;���K}Η!��l��ѫ�;�,4@,o��P��RrA'���%� �k#�����:��;i�|�}"�U%�#�г<��js��d�m�i�Bd<�S�̾�!�x��\9ģz��0@���d�H�=��ըF��|.W(u��1xg�󏹨`�c�z���;Wx�͊Z	��Q�"pI8�63}1�.�Hd��}u�Gi�:��+�\���v&�&�3��R���F��V!D�]��S�s�e�_�@�m�Ѩ1�c�X[��6�*1%�Q)$0q�(V����?yi��!YN+�1i��i�]C����r��Jd$�l4}��ގ:�F�P�v^h�s(�>v9����$����£�!��_X�6�+b��ƝT�V�p �!��(���XRJZ�0����F�˚G~�K]�"�0Fۦ��j=�肄{�g�\鐦4���)�o#�32���oE�r4�
��h`��<��y�V8���`���x�*� ��#���gDY�\�$�I�{�h�k`c �^g>�:9�aS9eP�w���=5�]�9	����y��1$D�'`�XkSh�D���&��>���9X�&p�t=-�|�[A�B>lKq$V�B	���Ú�Yz��@V7�Y�_-)�9D.��1�z
���-[�k��iKf��"�|~'!W»QO]�0q�M]D�l��k�^�zS�ʼB�x4����o����~A�O�������S��'�ݘD��J��0����̘��V��^��g��v������I�q��A��:u<�&ϻ��}:^P�<��C$�AHWD8()Q�8�L�ߴ`�,1�W@ǰ,��d�	�$��c��6�_mca{C>���y�w��H�o�<3�b=�-#V���x4���]�͐W#�������s)YAt�eS��ߑD��or� =r��Pa�	�|ñ���*�ZU�	'ߙ*�N��^,fED�(Mu�vݢ6m��9,1`����Vˋ���vyDb��<�+),<#[�o��F~٥��݀syV7O �rw����o�p��Ixi�?l㬔��������L�����c��y�����t�U�S��[UV�"� l�6����,��&� Ī� '��x��l�l�d�|A8�@�ON��eK���Q�i�.>�i^��+"��)B��1ǅ�b>p� ߽qEb����^K�p��VN���޾��4��cL�HhWm��l��;�#9�%�x�y8J�qc�%_��?�� ED:"�{�/��)�!���"8⎹;
Y�ȶ莌p�"'m�4]F��
�^XY%|R��GU��+�.D�������Oo���]׷1c�8C1�V����1	ah�o��mKu�^+n�9�*��:�x{��Ƶ�'2��h�nA��⯯���h��J؞�O.�������2��aw�8-�h�;�����54A��ky���қ�+����!>V�\fz ���*���PL.hr�@ٚ��J7�ִFb9[�R;�����&X�l�+�b�0,G�G�W����W��DH�J���v��q���{�l��4��6�(��E�g3��ܒUZB�󑩋���=��e�U��mf�c��3�!%��Gʍ�H��6 ���D7S����2t^ӦS�* ��5�˵{Ӆ�5H>#���J/��~��k@�h�h����0������W�rU_����ߘ�<�J(J�^<O�~H5��8H��A�F!:�ƌa�3�#��DS{��/���yo�v��7�.�p��ȺK?��-,
�4d��:
�Pb̙���y[�Khȿ+-M��K]���<��0�G���6�!���~���* ��1c�CwZ��L���_�N��w��r�!���Y�ߘr�W6�o'�Y��Jɮ��`n᠔�����&n+����� ���6MUw�� ��N�m��߹���7�U�ӕ%��#�F��G	��Q}���@9d�dӬ�����_Zn��:n�n��
@���w�����"}�S��l�f�\]��B%�9�BY��nX�C��X�U�fz�W����~3�e��!^�2��48=��5����B�@1(��g�������9����nwo;��	�)ۆQ�^�y2�y����`��� vm�T�ax3�wٝ�����9�O=���}�
���2������g���R����sn�$p�1z�
�qN!�ˇ�P���\�<?N.��喚�\ـ���DAO��/���ֽ{���-�Zaݫ�DT����Q��J=���:����	�r֢Y5�Q�u���'�;jjÖcnMn	����=��ą�,���%���
�%�K���GJ�3���y� ���ܹdC��'���թ�۫����k�y�)j1A)9� ��$ �/A_�����t	�����a3ES2�/��͛ߣ+;�+���Lo��n���TC&xi����u(��r�w�����s��`�����P���;��xP�5gǓεʄ����~�ںs�5�� j\d�N��N"�/�7s�����W�L��KA4��&�N���A����!GkP�\�y�>XǷa��:�Ik�j�=˗�Q��&`��{,T�̯D�t����.�堙.ڵ���۶D�7������v�;�^9,����HS��ds��%�T�e���0Y������Q���4��s���3B:��⾓YgN���#��@;��oK^�#'�{4���,}� ���ҋpaTk�q�q-P���	B�'�T�Y��~'�F�
��O��[�淹��]��%Ð�3X�E��E����.�p��w02h)��53�`j�����H}D<�|P���x���ZDD��$�ps�H����u�z�i�5�娏��y��m)������Ĭ�r�ۜ���]�Wg�3K�_��e?��7I�����J����L��w��N�.>��o�>�^tj|h�ҍ�KYJ����f�PN[)�e�z�C�Ac��*�>�HwG��F� �3^-cAg�D���
�7�ì"0�:ڟrM@���I�Q>��pIy^�B��b {�G�>�FC��83��`���P��RWsq�]��������A��Y��'�3z/ΚKͥǨ�rö��ޅ?|���K���r^Qէ�W�#Յ;���C�"�O��!�m/6R��-��=����]��\J������YZF`W��on��,$������.�lUٙaD;����tNKR�q���j�w�͒���8&`����c)�XGN�fI�Zщ�ʻF�9z�������H�����f6�'�!2kQX	�j��z��1T���!��q7��{�����{������[}5�y��ѠQ���[�?A�(�Y5�*��w��x��¿�RSJz~�tq�bɢSC�;��R�����Iɒ��A:�1��E�K�J�P=f�8�.O�B�5���\�K-���|�R8����P�Ucg����-���^F��Z�Tv��l�\8�����p�2H�7vx���%��F���b4,@������{��QS�3��W�KJ�Z���Y��cd���̰�o�5�	nG�Pim�"r�s,UV'�-�m��|T4���K8�|�;C��g�Xؽ�W���@]w�<8rR�95hǶð7+|z
�m��z�(7D�����t	�����[��	;TOgkm��d���|OgMg,�t��p��T�u��� �串���C��� �A�ИӔ7/���i$�&ˠ� #�i����:{����ӫ����:p���>*("=�8������{�~Z\[�Q=܂Y:k��$i&�D�p��z�.��/;��kҔ�?e�����83�׼!�����>��@͞}Q�	y yguߠ��c���zDTRpg@�Q�)�Ғ؂��KT�ŀ,�e�T) î�X��R[���^!��&�8�DI���0�L!G�t3��&��/oS��S6�Oo���Y�ftB�]W�����xGSѭ�.h�v��A�����o�DȖ_sM"S�~J�|�m��(6L�B�8�����5��X��MMc��7����/����k%�q�}��W8���M`�$����(���܁����<�uE�w��8��N�����
�)=I"3��I���ț��٤�<���~e|ЭI	%��U� ,�;������ ��./�h+~|��/�����x�bLI���[�7�%������Mm|�+m"JB�m��ѓ�sgaԊ�P���anoE:C�q��!�G�8�jeu��lfp���2^J��:U>9����ҸjmM�uIe3	 �Uf��x����B�����K �M13�c 61����(%C��E��h@� �V�)b��{��cԽ��p�?ir��} �$p��~>�1��6ݪۙ�9�6$Ӿ��}ֶ@{G��D��]�y�s���fePh@�����kƇ�E�e~�כ�W��Ks,������b�ҷM�)�j�E����#C�������PL�A��"�2$"V�z��.��c�t!�ǚj�b��HN&���
nZ������	�Z�va��.���C��#xB��&���
�� ��م(��B���x�/B���e&zfޮ��F�ʁ�=�L!�/eAuPHZ����@t��{�q� D��!��)�S0�{��m�������Z)݌��Iz��X���(�>���~"��N��>tP�J�W����1/S:���!����j�r�����P��`���<b'+I�����@pAX�L�M,H)6y�z�q��*��-�
鱌Vs��_�h\j��ݓ�^�I$3���]�z�%�8�q�;%�>�%Ϧ��]^z>�J����w��$������k( ��<bW�w-�&u�'!�A�L�M���a#[�ϫR$s_��K���ݣ&.��&/��ku��`Ւ	�4����§���VP��� ���L� �\\;�(*Yw�<*�W0	�K)A�S#�ˍDS{�և*s����t���CLH�o�L� �
&���O�t.sVT,V$ )���往����B�9��D�����9�jW$=�p������gg�@t?��ڕk��pR��Ċ *h�%7�!ՎSVU��<��3:<0Ӆ�!E�긑a�f�j�����N��c�#ǒ.Dt�|�٪����%ֹxwD�R�JO(i2$�>ﯿi�&��?��s����[/����a1�*'�s��]���&����B�$*����EPZw�T1��1�,�BF�yF!���a~K)a��u- :�gb\�e� �4	��I%����	�w����7gq�l{���瑱�r�ruP�,�7�%��"�V`��y���]�F�Ӿ,�}�;��M.g� s��v8���?�����0/I��XT�����0X�7�`x�IS�.��E����D�����Y�k���Ө�L3�A�繐g��O�� M2�q�j���$�]#�����Tj<��o����	Ko"�%�y��<nd��i���Vg��y?��qc����i�y�{���z��?�f헬%��o�[f��}��c����I��k�9��Z��(.�6R���o���jz���5��`�/����Z�*N�6�rz}��\s	6F�"Fw�l��77g2�t�/�&9��f�Qt��O�a{%Eb�O�����Y�ցySU Dǒ�i1jdJ:qz�!����:T��h�cozЉ�x}�%8�8�PTk^���
�)�;���(Sf���f������TsF���AP��=��Q��H�R�i�{�C��o����������z�6�\�b��� ��v�]�7�t�D�w���!ɜ���2�!]�A��-,;7��A?g)��%�9��V%IY��5�Ȯ������p���ҡeg4v�.�79p����)
�)��^�^-��@I���̫�ЅE|8{�-�w�$�sVo�Z�*u���=�3E�\�&d(W�UG��rA�c�-
NKt�Z��C>w�94������΍���
�ր�������Qk2a|SKGe0���"q՛�~� �'�榶��Ml��vi��EWD���{T$�Wx��5�$gU(��ɣ��{���B~�4��s�\,���<�<x��Mu�ҘVd�m���r+���!�$��c�R#pV�����UD�'%>�7��x䦻."�٬7k��g �8�n���p�o�?�kS1c�_�6Y���Z�~N����{�d���^K�.9c_��;�E,�;�2��LM�Mb _��n���X^b@`d.X�W<�87�b�&��1��t�?�����u�=��d�̢0L"1N�A0�"�[�@�x+|y�� \^}x��K6=ߔ�T[^�:T����(tz���Cp-��C��ܛ�P��r4��%%��!�2p	+Bh4>l�+Cvʳ)T�N�7�>]��@�)�x�'����mU5B/���8�G�By(�p�~a��*iP� ���c�Sv޻��e�p��[S�Ep��Hi���[2��Q���HH� ?�2q��
�s�g�7�,��f���(::[�=[~���CoW�,����||�Q� ��G��ҡ��E�I��x��T�ʱ� '�����]���ˇ��E�A���4����`T��7'9�U��^��)�'Hky��鬛��T#��)S��k��k��+�Su 7���u����\���-R�PFL� �b�M��/^�MW.aI�{���t��p���0���=�zA6��p �r�[H���T}[2֌��%��`;�ۍ"�6��	 xt�xy'�j �NKj�����)�g����*>�:�-���T�t�����ڪ\�n���&s�]�E�S����X[3߈p���t�!��WF����?�W���� E��BFQXm�rPG|*M�w�$��w'����8���T�q�R\tt��~�B�D�����|��?���\���	jb��:a���#:�����Vq�����eRӕ�]�T���J2��l�1�Y�C�R�%K1�\�;'��C�FtM����hJ�EyiY��B fpF*��b���r����2Ь��!\d�Ic�y���;��:�Ls���30��'^�.���c��bD��٥��>7�s�q�߆o=-Jn�fT?L�y���}����׎�x)��y	6���x�+�H��Z@k����č�ee�8�S?�"8����?�_�'sm�^���.j2`��$J�	�CO#��#�l��׷7"k���T)�l���z~����X�N �,�Xޤ���E��JwB� �(�e�Md�S���`�ko� d���_n�
0���k�ӣ�۰I��5<u�	+!��v���?�t[?�<xMC��yda(�Ұ�y�?�!Q�����)S�bܝ|��1�� ��fÍڮ3XQe����+�;}y�j"�H�����[������΋���H;;����_�J���p j���?R����ӅQhcpyH"�s�i���ڎ5���[�{�*����_�N����R~�<�h���=��!���.��%L[�2�yJCp�7���)PT�K�X���� k8���n��ʚ={=��K2�ܥX���x��k��(#{�F��qu�~�"?ϔ"(��Xr�m ��@`�O�����Ҿ9�Ss��&ߤk��(���I©�๐a����(��;VƑN霻�nX7��_�ߺckJ.S#i� MPѱ���ǎ��D��|4�����1��L�����r{苵R�J�S�O |�8aSNJ�l���Ve�<}`k�Ǘ�&t�����
��J�Ju3��ǼEN�AYJ���"IؗN��jݣ�/�$s��m�i�7�Iq�J���q
�ɢ �CPG���n.��\%��7h�N�b9s�`���ƪ�j�gs:�:�c"ⷌm��Be�S0�6�#+�h����\����Rhqub�����ն��>��S�Z��������{���^��dW�e��]$�+~�+S5\,P�l#)y�t���쁠��K/*1�~�#�V
ve���'�|g378��(I�|�����Ϻ��v)�݊hv�*8�܅�^�w��w�\,�i�7sJ����u���1����4h�yT1��Wk�PwG0��K2ЗI�������[��p�p%�-�h}B��6$A7�|P�7��(�6���O��'+��̡����?�}�����e&�=�嗽[�l���N�:���t�z�LYQ1�u�	���>��4��p�<G~�(i�>����$A �I�z^ ��wDH���*�r��)TDq�w&�q]�~���A�I�._��t�����e"؀��*� ��B�%�It0/�yo� �
L*�8��2��_t+�=�=��]�'=Y	����2�n��L|���
b��vG����y:���󽮔��Դ��b�[~�{kg�������)�fne�&uz�����íݐF6���>6��F�z!5H+�Bk�R�Z��E�S��oI��"��Qde�3��x��s��I�d�QwRN���lcqMk����-z�N�fn,'�(n����a�n�o�m��]~�<ǆt���yO`\\o�z��-Y�e��`㓘�
ᯱu����U�����;�,��,�m�Ҏ����n	v��|���3ق��������WP�ߐ�n*��a�C;���n
�Ѩm��U�=3%��d?L|+w�V��c����elĚ�t!���u�����3�I,�Ґ�w�h"�4 ��K�$�}c�
� MK�K5i�m�u��d�6f��v59��X/�����SA��&*fy~�4��?�-�%:�֝���k���ث@��DG���EVQ�����>��<�A=�2)״�e�)�s^2�����f�`�k�Hh3�(A�{�ut�&�5+��>Y�j�O�f'Վ�(�O15���{ۙ�/Ʃ:IG�(!��`��Iէ/Z�����T�<:��j�y���m��@U_�`r� 2�����ο�Q�DJ��5МO�T�~�_{Ք{�h�IQ�H��r�~#�����;�C>����$́.�`�q��[����M)�o.��e�!h�h�:����%��u���NtJ��4bS�.�7Y�J�pUS��|�%>B�.OrM��W����FG�$e%e� ��2L��"S�Mn��U�"3�'@#ń�&����3`q U�K�!J��,��\�1�t8-,�;`�O��X�.�:�5��?���e��}~�m�0K���ү��cb��ms���%��� ��BEB> �^X\.�I�|�����ь�f�v��7��*pucq#C�I�Up(y�{�~ion�����)nYc�N�F( �����?Q6�BH��Z���VR�n�� MFD���u��;�^�Z8j���i�|k�{�b$�l���^�i���Y�k\�2�$>Ą�y�{�e�a
}󚿤�JV�5���mY�F�s�K���cѡ[$���@�Z��0���9�vyz-�z�d�Q��b-|�<l��H8����G
YI���w�����_�\�JX��m����z�ՙ���:#X��U	)���_��3�^��ϒ0����__>'XӴx%{)���az`}���R&�'�>�c�q�����ړ2Z�#2 ֕�.��l�������X�E4��/6�gC��E�=^��Cԓ��.�K�����v�2�@�+��%�:>��߷X������_�ӥ�L�+ҴT�)�S��� Zْ�=-���"G���Ֆ�đ�Xz�EC�|��KC@���V�� 1!��Qx>�����v����8@�� �ؔ1�h���i���=<��"�Φ���J�v�\P�g��6�e8�m�2��Ԫ��Xwy��OF$��9).��2��=�������Y�jm�˯�f����@���1P�~�Xӽ��p&)�Ƒ�� �(F�������n;m:����	��m_a�	�ԧ���+}�~�*PL��/q�ѷj��1��y�c����˫<��k�j�b"����%���D�K�L��*�(��H�#���|���3(�ƺA�lPP�T�S[$=��0���3�8�a���l��{�bS�]4^�_���&�=Z�w�oC�)�K�)��:�H�����aXL3l�x��l�"*Oa<�bA���۷����%�X^p�?�yJ�K�gcAU�C���?'�L�9�M��&t@��.c� ���N�c���"	B&j���ƯT��1Y|�u;"� (�̲3�e�'(_�]�@��*�?�p���1d@�n�E��L�S,d"��)���2
��@�¯�E�I��b�f���0X@�9~�����	b��gW��=���t����`�5<��h�U�tuI��/Z�O>l�1�2�D��#?�"w�Jq��ۤ)�ҚS5c�d����ə�f�z�$���\MAը�$"#�y�%Z��'�t�r_��vbߋ�ކ�F�%��[��(�j�Y��Yښ���/^0����:�nN��]�s��j9��GFw�nJ[�IoK)�*'"=\ǧ���0�}L��.CfH�y*�[�]ЗVȗ�DHy����.ۆW'�x)�����1ޝ&�$���C��h;X|[mW�U���S�~#ٔ�+�	Xy�'+�����*��$0���QU(5Ű}
s�a�O�O7j�)x��\{K\��pYIXXyflv�G�Zk��vu]�s����֥5`[s�wK4���^0j�/��{����`i�Ѫ�$�;��E#���L{�2�u����HZ����fwKR�K�rH;�R� �3�2I��\Lr�#��y�{��gw�S��{�+{���
XPO���ZY(�Y�_��;���7� �����-���'T�`\tCy�sr����R�':��1g7�'�� 	|0�t���E�ŗ3��t>leTeEϛ�m,2��َm*!�S�0�PH-�3���1Z"1ٕ0)��ҡ����f�_C�g�i9=4�M㼛�;ï�բ�م�M�^ժ���S���N=���8��v`��]�S��4{B~6�F�\�Vź���ލ�⠳�R�jZ�!�[K!�,��p��'��$y�Z��Cl��`tf�-���?[p�mUIK���p�N�����(䫖�Q�g�/}F��~G/Y�?�9lVJ�D�Y�S��R���z�-��7S?�"��� �R|!���st�:����4�2��7Q�-�m��x�п(��H�m���(�~��)8c5QE�{��!|�»�� }	�ӆ��x+7.����%�5/�Ý#�I����[�8
�A\?��U����?�H�?
�I��ə�֡l�,�q��Fa$��(S�
���td��8�af��:)��c��I"������)�U���ap
ʥ7ARu��E��{�^��D����a=���! ɱ�eց*�d��[�SB�{�3f��G��7��_��@��i�!V4�[p8�R;Ƃi���D`xҊ�0��U�P���ZK'k6����D�-X��}r���ǚ�o�v޳"?1�&��U�B���(��̠+�88�ķ�/��~}8�8:�@�I=cP��)��BA�R�8���H���=�������I����QbD�;��Oty���@iY�̼�FH^���ܺ�.:e�Mg������v(��Z��Wac{ӝ�w�/"�1QHG�PK3lɱ��(W2�;;�x萛] T�5B�u�R��l����ʦ��
������U� �@i���-�+B(}���OmZ��o���>���ȼ&�Q|�p�����،��8�������,�;S�W�#F�R�zԎ��l�Xndk���E�W�O�	7����(��H�� ��Yj ���eP�z���zCd�^�`N:��qR<�A73���h��Lf|�=x&8X~�2��?�sͩ�൉�Qͪ$�E�I����]dM?D��u �ă�Փ��߿��!`ǡ�ߴ�T�(ﹾ���cIlp�ӷ�1���^D(��~�i�|J�RL8�v�p�@��6b��.v?~�b�N�I�R��/$��+p���~��5;��؟�چ?����W�9��o`ze��1�	Bb�{�WФ�:���w!����^�w^�i��l�TQJAF�A��Dٴ�_�[�u}|u����QZ��h�5AW���:Z����Ms�:�^��R�?hda~g�$k�f���_??׽��tS�,���<�RLb%�r:c�,��M7}�܍��F���Xj���
��i-1>�R`��H,������7� �1�Х�4��O�v���k96���z�]B
�#���t'�Bl4�6D��ҋ�ϻ����rqUS;�t�>�3���_�C����S�6�R74H��?��'�s&t\`����V%���[b�ͯ��wA�� ��H�o�bq���'�4_���|��y�`I�cD�l��Y2r���~�=��CMEB_"��O.��848���(郸�ͳ���;��CmOt�	�b����P�����.�cއ�ڮ�v֔A�Y��aɁ7�:=����\�ݗ��Sڌ���C�E����&�����;��%���F1�o��B,=~G�0ݏ��;�Y�4�_`��X��0�R?�uq4��v���t��W���_�$!�kW��Z{���>���$Ul�!M��쿧����j%�ygd�Gu9�JK�xq�%m#k؊���Q[h�1�Ea�\*�	],�՟�^w^�N@�m���p��O�o�"��ج�-V&E����=͜ü��g6�8R��lRF�$�`#��O�e5ƈ��WU���^�����{���J�㾺�{o��l��X�t��%���*6�Շ2;��yЬS��ݢ�,����Ų�մO��佹�Y�޻���2�oSIdƑ�Fu���ϝ~��w���,�����)���QWq�>���M?ߤj��f�*I�kaS�ֿ6��qy�6��j7���uڌF��,�W��&qg��1����l�Ota�M�9dw �5��Q�/�t�T\87 �]�	�FnwP�2=*�*B��L��-<�<&pF�j[���<Vx�)d��s~q�����?�h��"��XD�I�1��*c_��F�<ޕl��V[g @��4T{wUM�1��Th�Zͺ���m	���'`��-�q�=�j����ٕV����L���Djg�-�Q?��)�ߙ��-��<��=�z:���K�dͿal��v�8R��´�!C��	����sIm��6t���7l�z����~�"v��G����~��[�qá�DR(�ڈ��w�z��s��d*|;�+���94����䔣�c� ��X�:���&��R~`��uC������{œ�&��c���W,iP"o|n����]$b�Y��=#�}�B�s����jJ����S�[´e�Gj�I���%`� �k���2�[k�*!č)�%����Y�j��=�~_&ܟ��/)t�	�������R������e�V:bMДl 3�乏O����&�I4�R]O�'��g�`}�x�fs�&re�����m�TgV�m߼�Ӑ k�bFe��zv�Ȇ$��1O�X���_t���h1lm�ZO�z >�evՈ¶ �	@�Tiv�_���.$BF՝�]P�\qc�^~'��Q���0A���>���75$�;��IL���3xdhV���a*,(B��|��o�ۆQ7�y|u(���ف���|}LI����"J���β��`9����N��W���9Zn3���Z�#g�
�Y��b�(���<�3ډ�HӵYY��g�($FOV�I���(
C-�u�YYA��c���(�n-fN%	ቄ�6Kd��|���}X���*N�v�h���(����]2��!	I!�W.�o�#��E�N�&Z��r�4�gf��w)<��b��M�z`��	'c��C�+B�@i�e���`��#�Q�����$+�9�
wQ��C�\1���=� �%ӽ.��-���;~�4�h0|��B���*?���~΅q��A�鳈S�b_mȭ!P���w��>�����^��w�0�QPsBR�g��)ѣ�*�۱}nDc�RGx���L�{i-@T��.�V�`݌z�|^�R=ԯes<=��h74z�_E��b���o���KjO��$@RH�bV�JSzacO4SCJ�:�i&_���:��dV�f,-]��ז������%Ƙ�n����w�!��)W����9�G�*m���\��_���s]�㚚?�!��F���� �N(E}�[�x*�Ȝ܋8-�ނ��v��m�%_�6,/p4����ƶ�&���6:�����i�����������E��ï�g��)�SoF*��� .��;�%��fw%�;�0�mJ��䯍Dj
C9�k	���)���]J�J��6vX�$�WVUz�t��-q��B��P<v6~��H�������b�G�i�^�8,���;���eI�����x���:�HSsyLb�0�:Հ�8s
-M9�]�fc*�;�~���QZ�@��8��7IOg��c�<:�62A��8zh�GK����w�~h�E�w$��(hs��@�e'�Lk��JL�����縻V�	�S,��Ll��D]v�[�),Q06pRH�����Z��[?��wFP���b~��S�)�S�h������iN�	^�N��tS&�X��I�/��E���^���SN5�/�}���]/����hgS-�/���G�?���:�a}?�,IB�Vf�O����B<���[��:�
��/6���b�L2�F�n�"�ذw�X�_�t�,p��Hlti�"��rY�
�⍱V9��,�*b�C+<���Xog�v�3�Kx�@J���5%~����
tv��c�D��ф1).��ũ��O@�Q2����13(�iZ.vS��mQg*IC̬�T�\����g�o����H&��թ��&���S��{<�:��Lu�$K�r�	�(B�vF<���N�9��[�F�?'}�u������YB���XF�G�v��F���L��&,�靎:�s�'��HP��O�iSa]aSц���Ĕ�g=�a�B��~0&!ب�3���JG���*�'g�m(�A@�٦���L���L�<�Ca��0/��uBYb���m��Һ��c� ��E����덅�X�$GK9tOaB��Y:�A)N��u��(m}�Q��\��Pg,+���5m�~�Pbd���+���>��İ�8)���"�ӗ�퉏?�̒9���7e��߅B7+<�?���(ݩ� �$̪�f8����W���^6���yyN�9T���P�3Ȗ/[9m���}1t�Kw|��u��y$�')��r�p�|o��;e�=ș_�t�O���(xs�a�a�l�b�W������>����n��[׆.v��M�;�31h�!1 lײX��rq��G
抈����T��gn�ё �Nѡ'I��T'WǗ-��bv���P���O�����#�C�;��Hw��aҷ��>�_h<w�ǅ=�e'���A��"�������vI/��Vݸ���9ݫe��z����� �Ak�'�T���^��3�y%p�K����ñ�}Кσ	^�:���,,���_@�`p���8��=A ��U���&����t[M{�.����ӳ��?y&�y�so�j�orb�C#'Z+���|Vh�S�-�����Zb��5�9�r~ 2��'ȂA��hrF�NM�j��3����&j���(�E����~��~��z���7*Y��ض�@0/�9��P��22zs�V�^"іfSr\�}�)��Dw�5�\C��4���v,�0~8U�l,s+�2�?�n�L�NO�
���o�x�(���0�[LZ���=#=fz�+��9m'��W����dB�5�~sf$0LSg�ӥboC=GP��0��w��\H�e��]���²\��<������n����/mߡ�#���)�!��w�Y|��(G����^����\4�GӠ���u4��()�0_�d��1��>L��VW���c(�=b*
���P�0�b�5U���,���+�a��-�+���ŗ�3�l�b<_���=Z�OS#����q'C#���at����w�����'Z��+���%fi�א8�����$�:�*\�g��J�]�)�'�Bʚ��X���:�����Д����_��D�<O[ Z�Z�6aܣ�÷jRo���Rt�>��E0)o�й)���ϣ,�QU�|�����!^��
�}-�� rw���)ԩ�M.:�� �SM��&�^����xo��=Gg��&h~����p�=��W؄�"O-3'�W��V�_��9;&_�ЋR7���^+��.85:���=9�
���
=�®���V����_�}E������c����I5H�]�SɎM	h�"��x���G'!�/����+��D�nǕ�	��H�����
L�#C:ߋn��t0᠖�QU0t<�HI����-/3�>[�������*RQ9�`Ŗt�MC��\븞;2N�6���kɻ�@[�v��
_kN/��J!�k����rqu%x�y���,�N��E���A�������,��x���*G.�~$(��9	�!S�A�O�gd�	��k�"��b�[�m�>��-#��#�Ik��A�X�]V��H]S9m�B�G����$��� \�J�Uz��5�1x��qT
���K�AE@������ā5K>F�,^@m��iC�Ӽp�.��^����d=��s�x�8�}���|l�Ϋ��A�R96j������b=˰�)HKH�[<D�-��t��f"��Y�v���`.t G���CI^��;��D�P����
 %g�]�9s4��*��;xON��'��1*��t��@�ZEgY�+��{���Cɾ�x�����d+}њ��h���-�qD�0b���c��#�М�<}��N��؄ZYLXWX����9Qf�G�kjK~�$�p������@�GN�"����|�}G�S�o��G��o!��&�b$4���2t���� V�l��E����0��_�t94���-pN�a����sP�ڈ��Sx8K��^*2h�Dz�H�d��,��[��v����vDj��`n�Ig�te��+��QW��ux��k�"�X���K���������^���O���!����5߾ ���f����2�s�5�(�����
��ڊ�:��d�G2��0<T�	�g �.<x�I �GP1[2'�(ٯY�E)����A����ULf�6;cq���9��'?_	�o�ɂ�!����'����*��&	$�YY�P[�mrp�l���B��rf��ҌN�|c�KeWxۗ����	��]J}9.��f-pP@cw�c�ꄕ���6̵��iC"��U��U���]Ɖ��f�|8�6�FK�㛩�\^��[�� (P1$���6xy�>oLn�q[�!`W�$����T��ã����錿�X��m���Z��� �e�P�9v��E�<#$����e,s�l�2�3��ԝA5
�_�!�:�lG2O,�0��W�"hD�VzD>zy�Z��뤀�ʆh�P֠Q7rW���(��)i	"�mI,L�戨��!U,�c�� ��V(�qꪀf�C��+������.��ߨ�����M{�m�ϛw�ai���y��������܋Y#Z&>����mgm,�wG������k!T"��]@tP"�$�*�y��C�d��z�m&A��j)ƹ鋼��v�V6����yn�+j��֖��3r�M���6����C�?0r��57Z'�N��!��j�Z�X�;��l��Ȗ�D�6�:;��K�A��S�%����9��}Ƙ�N-R�4V]�߻���oW��	�$�-Ț���]�q:�k��1Q�DA�.��7]�}����-��Ub�s���V����ᖩ�n��n�O�ں�a�o;�{8@�l!��S#��Ha���6{ð� i,}$E����@{p��/؉�{'�y�x��P�D�mD�,�~?��#3E�b��s|F]�e���<W��4�������"`S0�<+Ay`-s�Փ��RT��O�7y{�L�?i���������b*,�9j�+F৶����Ѹ��g����K}a7���aܮ2�5��^Kh����o��H���'�6��B5�N	�� ���nƱ�4�h1�9�"��.3]ǱlI��b�@W������&
����ԝ���6��|n�R] �Y���[R���n�`��e3�>=[�kh��R�G�_����Ey��k%OF�����3�VP-O�@N�Z4���hԽ������S�U���('x�k�4Ѣ�+�ͧ�_#r���s��"3�j���m��3N{�$6t�����+F#�Bd*�"Чa��vK�H�$��5\����?���-\~N�`0�ކ�%kx)�e��X!D�pŷo���M9�.q <�;s����Q*��	�"�j��������ڳ�K)��kQ�oSO�o��uKS�f� T�M������ppX�3�V�D�LM�I�h��P�w��"o��G�;y�	��?7)�}�z�\F�D�W�M�K#+k<��4����-��j!-��qq���mi_ĥ·� �-s��M�Y�{U&����:��E\�i6�Y�f�T��W�!�h-�~Vwy��(n�~�F��&ʔ4=���|��{�yX �!���Sφ|�yd
d:5�e���U>� ۆa�6,)֒}i�O?l%��އ^�&j��c=X~?"�i�\_'%g|��	8b]O����dܘ�1M�f�,K5b�E15)�4�Ц�4�cv1b��x�fh���'�\e����c�̲�o�p�i,�tss�i��a���Y��:�Y�D3xGQ��Ӵ�K.�(6~�]�x��f�Kj�7��)����O�����Rc�FQ��ڲ��`Z�&]�o
����G�E��t�P\g��D��E���j��qb}��}�'��)5ٜz6�7/j�&�Mv��>2�K+�Gb�?��|9�����u�7��)�$��=
)��d�0�Z~vۂz�y�X$ek���
'!��fo�^������h,�`,��	���u1��=�va�+��n®Ͻ��ET#��$�?�.hh���RBk�7���֘�E/�G�|��9���P�>Q�����Vi�Ʀ&c��D',V�C���Koc(9�6�DZgF}�s�.@�Eȡ(;�՚ng-D���sٛ�t����z㴵�S�-#I��h-�H��5��[�s��o������C|{@�c��a�/�G/����uD��	����7���Vd�kT�m����V�z0SUvS{a
�j�Y_���=�kӒ�4�*d4=�����:���WΔ�[�2E���	5=�k� ����4���M��2
ͤ�6�Wd[l��9����}ߣ�@y�sm��3N��L(�R���1�~���_�b0��e�e�s�Uw�ObMu�8��_�Eug"�k�~N	�����Y�#�r��h�'8Y��Pz��p2���Y�Ƀ�5#���6������nk���|����2�uӨ|�ُ�1��K��!4:�"׷����R��l�5i��ܶ�D�(�Z޴K(CA,dFqܮB���(�Ӣ����y��,�r�x���-���gMh�Gk���z��xm^�������'�e��K�F��޿�X��B{!	S5T2�ʌ���!kU�yݍ��RQ�P#-wS(z ��JFu&�����n�����:�ү̈��3گZ�M\Ţ�Q�����B�6#o�SH�5x��h�͢�!$h���� �A3��	�:��~�8-Ef�/���!�P��'e.��`eۖX=�s����\]\�f��.-��z�����ċ�H(�nXr]���,�6��qZ?y>D&Kg�j^�&�ތ���N�����aM�mjK��o�ۀ�uN+�q��z��hn��
�X�Tk�zP�	�w-���;�"D~Hc�ə	Y�N�?���7�c�e;����+�HL͂5E}����cY!Q�vZlY��`4��XW�w�ÍPnK�g�JM�|Z���R�;���f��]P�r,���2��{k���9sW}��F\	�`���=J�p`- ���M�q�k+��H�U�4�A�?U�jm�u�Ѭ��vK�!^}R���!h9�m�>t�S����x`>��8���љ��ڔen4L�zգ�{Hbs"Ӏ"�˗��29!�����ߕέ���g���^/�}ML�}S�'�������Ńw2���A�-�K�W V���f��t�a�>��~è��[5�-�PKl�1f�h��(o��$��%��#ׁ�w�M�&�#;(d��0�#@Kݳ�٩}�?�/uA!�!��?8���0T�XL���z#�w;�+�@'y���YQ��	������A۸Scq�A穬eg=��W�$>PZ>�y�~���=Ep9�Q�
+���[����=���;��7"�b��(�-u�~876��_�P{P�!��q���Z��n�,@�D.3�*�t�/�o��!!��g��"�}���<'C+��B���p|i�n��u�Jɰ���,~���KJ8�Hoto���@`�T0��@�5����H7���J�D�4F���aF�=���YJ�/��uqz;�4xPj7���?�Ƞ��>%6s��?���[��4̱�:���ؕ�U�$~p�?�� Y�
���4�>O�/0Z�J0������G���fE��&�����/G;R����Hx���:j�h��3.���a�.;��h�C�U!���3>â�ؾj{���;��[����y�ނ&u
ѐ&�<�^F�ëZ0������|5�]��� b"]���U��҉s�7}�u�� e����@4�nM����,�O�d'�P��,�-_�(�����(��?�{�#V�"@���8�ʹ71�Ϛ
�J�)�w}O��pJp��$i���)��8NY;d2ju`�"��&�/U�=�|4�[L<(��Ӿ\�:��w����M���=��P��ˈw�Z0�U*{8$@�n�Β�z"�){4\h ��9Z]�%u=Ff�z�lL �1$g9�?��H��XQ�� ���fM�2F��{|(�0��#R�6P�g�T��=+V��#Q�;���v� F�eJXLrfl%��C-j~�˕
P�$����O�����1f�Y��%?��ʪ'B|�|��1�֘��18�[�D�R1(��-t���CA�>����_�va ����g" �cMot�љ>����f0���,=c(�00"1��W�J�b���r�ĕ7b��)�%��JE�KM��S�%G)w'�U�FiBV��MULl����Y2mg�*��xWo|<���L�_Rt1A������9�O����Ƴ7�8�O�f��?n��)����Y�.��
NQ%ɑk�� :�����W�K�/��>q��>t@]��I��N���Y�0��a�F\��������[�@H3�y3�qy�4�f�Ͻ���ۈ�b�~�������}��Vl��@��t	��h덏���ͺo��cqFo����GA�%������� +�-���/�w�R���9�Imt\�����[d�a���eRy�H�)/S1i���m^I���:�moN	:�o��Zxʧ����+M���#ǧ#�Cd��)ஞ�����N���Bd΁��q0��6�r^�DV�M�ճ��Q��&�3�� H�@֒|"�����v�(��-�A/#�^���%���x;3'�'�7п����}r��\��ԯDP��ٕH<�g}���/ ;��	T��bҭ%��C����ﯔ��)WD��Z�~��/���>Y��&�g�9����F��Y�L5_?9�Y�9}�Zg03O��{���t��Ĭ�B~O�˺���)Un.���;� ��Ҙ�L�E��n�Ǻ��I��׺h ���;Ǎ�����Vjxy�e���@�*9
6ɷ�{��G��:��ʺh�c���-��7��W��f2������#��$Zy��p��p�D;o���"CG1ZF��oX�/�(I=�rs�?�m9^=�?���f�e\6�%A�۫l�e�^�%:i����n�@���c��[<�b�5�h�o�l���_CAP䗗 ������4ڡ��0�����7���IW�)���r���kl��X���ҧ�YcJ�a��^	^t��;�hr�6�Ձ��[�
��U�;�b%��N7��`��F��ȥ�xT�\`"0�V�
+�UD+'��7��.Z�� }Y_$�r�ْA�D��ʦ��*I�K����o|t�s�:ML�1��D�ϔv6>�� \��i�+�k��q{��sq1+�Vn���hb��S)�kG��3l�w5��qz����ώ������틸$1,�l�1�
�ϰ���zX��'j0��"���]�2�z�M��`Etb��n�8����yoS����C�eX�a�gX 64���n��O� �Rq�z���YC���f�#C���Љ�Z�����O�q0^/Ȳ��(�ˉԠ��5���(=�>���ٴ1�C5ĭ�j���f���;WWwb�}��S%�h��P�m�:���0��s�- !�}�H�JZ�]��|��"�f;�I��m��7`�J��X��+�(���c�k&� vTz����: C�2@�qW|��<o�����74� K ��+կ�c�nCM�^�����9����V.?�>a�)�2N�����5�9��G��ŧD��d9��竻�ߛ��q_�r깹r�m-@�\����y��&E��6������B��߅pM&y����Y�,��Jѧ���QYV�3;��H`�%�B�k2��WȄ���h���	���QqⰣ^��
o��v����M��8	�V6���K�K,�@J"���גTI�9#��7��0s��U����~6�(J ����.�ǭ5�)��X�"h���޶�e��󂎬s4�ۖ1�fe��h.*�!Uh)T`�GD�Y��IQ5E�i1� �r���J��J���"/GT�x���0Ei,۪Y�"�%�m��\,�<%;���&��	�䭈��3}?����@6�x/�`c��$�"�fg��2z�>%�i�a���H���-����c� ��>�u��]��\��&����=E�׹^MN�Y�d���_�-��w-�� x'l�,�lԢ�~>�`,ni�Gx��pVje�U������?�����==񕏊�o���_1�z��b�}�A2�ZS,�6��:��p�&�s�$���`!���1iADP{����S|y��5}�(3�cS&��'�;�;N���}���Pa�]h�ej�ZF:�34�emދ����m�OG4AП"�4�9�����M�[��A� ����te���k�\u̞+�GN���.W�����s���cKF��=�@0���� L��92u��g�Ӄ�r�68|���	T�\�c��l� �L�с�ؙ������_5lB�ڇ��i:mXE��l�P��mpQ%/���p��@Fd񿍄	2v~q�xU�L�;8��+�O!T��'�h.\����X�!ȏ����I�@�H��YD҉�ƺ�!Ey .ݸ��4���r��0����;⌠���UdO�ץy��y4��@��n</Y	��A3�=�L�7u۴���q�Wb�@.�4�>���IX�.o@��Qp\=]�J�y�_5e��}��H&>e��[�,|�N��R��k��Q��n͢Oᗲ��UUI�@�-��*;kn	�X!�O��<�h�օẖ�=�X�ƣ-I'W;K+���j`�!��^�m�A!��ͫ��?�Di�&(7��%��l�����=���3���t�wj��}u�Z�"�W*%KO��,�M��̞者�e` ��i�R�K
�?骢��D�����(Y�� yCX5u�U�¼)<�"���V}���v��R!���Z ���;+
dJ,�����M��zgBb���h-ڮB�"��������;��E�VC�I�7�=ovbm�Pͺ����5�*����+|�d�����ϙ�_^��w�(_d�B��D�C!��q󸘴S�C�)@l/B���H2�L<J�pY�BMiG7�>1�t�~��VΉVduz1����
Y?C��"���vd'3�btS�n�\�P��t���n -�J.�Bd����ŹnBT9����%lp#�מiz�Wu�[��y��Q �"���G V]<�kq���:��s�T$ȉU�@lzȇ�����1��Fz��i����L�;���h�7��B�����+�����w�����{ ��V�B�#�,�0ޝ��Ý��uy�X�64wD!��LY�O�.X1�%���_3��߇V��&��6f���|h|�F�.\'eýI���������.�V�΍��������0+�Q�%Fϕ~C,� 3'��8�"�:V#($ݭ#]����������F��>��H�?~�=�>��J��X���鹽������6\c��H$p�!�0��"��&���EK�c�u����_��i��jS�w���%	?���J�%w��>9�w�s�~M����'�g�� ��D`�	�=�����0���叜"Lv��
&��MC��D�D� N�:}�kW!~@�� ��v����z�x���Qx�&th�6m�N\�ba�yͪ���9�q��]"t�2Q�x���(_N�V��e��{\�ѹ�qM�$a�d.4E3�"R�;�$�̱���i�:�WM�/Tvg�~T"�/�&�{D%ULĹ!�}_Q�	:���U�頼ʹiU	����H��8��
=>&l��0y�C욀#4�f�ΰ��+B���+��q��ҁ��C�}�k��u�����'����2b�0�>�>_B�����kVq�"+T�FZ����t֌��sV)G]�3�A�z��q���9��sBi�A�^���|�Y�-I��$|L�z�P7"�?���̼f��M]u�/�|^>	e�y/x�	5k�-5'�׊��8~����G%�I#��V�*�=�s>���>��&c[(���d�\�L��n�aH�"��:�W��ۮ�h���[�n&0j��'.dF�֠c"�<"%����μ�=���ϕ|;b��sU*s}̺���^��k���x����e[6B��I��0	�m�:ʠ�	� 	l�f_��u��#*�K6��3�Ul�N�l 쎜�y�=']8L ����J	j��A�/⁮��Y�$�&�]��Pg/�g�����F�J���q����M�*���{YPM��ni�#:�Ĳ&��:� L����.n#���W�v�j�A�ꁄZF��`��j�
�`4H�|��"L!�ԗ���]ue�����IW�u[�o
^�=̒�&�h-�떛T�*���F@v�K{ϴ;�Jg}(�s�EE|���}_t��C���I'�DMsHS�!�x�q͋nR��6d�g��ľA�A�W�k@�Y������5�	�b:7 �-I����R8��������r�X��^>��� �j0�i�����2��V�y`���P���PI�}�G�Ѷ*8��\�������c'j͆x#�"[��ſ��P��ɐ+��)�~�$lWg]���1	�1Έd-����ɀr-he7�l�oD�6G	�L��g9E$t��$~��X�պj��s�5(̓��S��k��q�p�f�`�Gf���D��c�`x �J(W*���L${��x:G �HL����J�UwV�"�5������2�N��߭ �I���߫$ /@EBփic��z�r\+�9��#�m0��׿�°��׏���0��L\'�o�1cݸ��tcӧM�5���K.S���jcV���1���u���C�����o|��W�U�޼{��1V8�G\�T�� 3��چ��h:��0I<.�uRh�6!A� �O�e��M��ɝ��V����N�gH��sd���tP���n��=ƚ�a�n��`d.�(�6��:-��W������6o�����l�{3Y�w¸�峚�9w��2!B==�1��g�JŶ1�2���SD�V�&��t��I�ĒB6蜪ޢq0���4���h������}]���$�B8��|Ƈţr+�tKD��Xў���/���x�cr���|z�H\;]8�7ZӧiQ�G�J("F�S+�7S�f*��NL�(�
�����"5�qX�w벭����v����D������G�094Z��ܞ������6-�L�$v<�XDc@�/	k��-�ɼ=��{��I;b'<�Il������������s�9���b��=�.!������Ðf�ꅣ8j� N��w_b�1�Tq>�m�EJm��.z�o�t�hq	������7��A\��������w7%T�+�KD�'��ڇ�q��(�*��J}�R��Wc8�p��9�L���k9��+{���_���@�X�{㠵��1� ��g1g��#f�tu ?�Ї��3a9YL9��d]ۗ���[��:͡���7�m9���s�#I��z�).�Y�Rk�|t�a��f�� ۧ��ЄC�������7H�騲����P��j�lx�:;�ᛊ��6̱&����gN}�ҭQ0�[�h�s2&�����	���Á�S!�91h<�hԿ�3���p�������!�Ҧx�	H�S6*4�5�b�QM?S���3V��_���5�@ ���ǎ
vHϖ�7� z�i4���FF�-�\�C5'd�y=|F��9@�)B?�`f,�gJC�"��ړ��u�=��[�r���/����U[Y��FZ�cXb��T1����n�Ql�=�Im�Z,�-j<�� F�^b`z�c��6�� <ē��T������i�ڕ�}�B7X��X(����Ҧ�ɕ0��Dê���rۚHLa��e�64���
���JE�p�R\�:�����Z���r$^�8���j�8<hQ���f����=�~�J��Iq(�sQ�، e!�f�g��|� ���ˠ|��|��fY$��A�el��e:������������8�sbk��+
Xx�Q~I�e/�z#
!w��`+�hO�s�'�LT�H��>�	r|��܌�����r�Ű. ���̩�%#��R�����[#'1h*R˶o�O��,��+��;��{���!�bؕ�W<�e�īJ�{i8[���vEMj�W�G���kl�D ́��oI��r��O��@�Fmצ���������ͽ<��Ap��%�j-����9a�6��Υ�b���r��ԗX6��=(���D;i@x��ȝO�`�J~�ט�\F�޷���D2\��{ YѢ^{c���4�}T{G����'q��ƺ�,��(��	'��o�Zn���ɮ�Ia{-�؏D�����
�߇����!@}����E)�}y�H�h>䔸f�fN&6��"?�4���x�7�9��w�ߢx�uP˃7w7C�S��$��^duؑT"i�M�ėQQ�z�:Vvɔ�����
Ӯ�)��}�(��nL�h9�a�Uc�Z7�_i�nv={{�n&G*Ӹ	���pW���E��8[S�}X3b�v}�����3��\#~@����&M:pH�8��L$���S�����``�A��;���k<�S<�M!�f;y����(�ͽ:��&_Tj��&�������hX�Kʛ�2H���e(�s��s*�ٺ(����L:H�N�p�1�yA�D<���ԃ�/�R^Z�Q��;1� �U�ߘ��Uk�D%�J�A��ؠ���1�����0�����d7*-�x_���yLi�A��@0I*�B���[�0YM"���J�T�ӳ'v�5�Ma.x��>�dzi�Rԇo�fJ F��z��{�va�A�UL^1!�&x�.�0>��ڭ����#��ū�5��r1���P;o!aY���vH�t�;TN�3�ε;�Nq���~��G#���t*/t��90��S�!�q��5$��ó��Cdk
���C�fӤ��3	����O��XO��������,������&��z�����<4Eb����}Oծ�K����^����х6���9�!��	^3������F�D���z��@̠���ND����v1���{�r�6���.�[W�K�RtfC?��-��Y`����(�wm�O���]C�k��(ζ��n_i�Ձ�����ʀ�^���&��=N���󓏀 �ΈN��F�፷�����锪�(Ƥt}���y({UV��/޺�}"�x��0'+&�j�����B�zs��x7����J�ܖ4@��Y9�P+���a,g3Y�.I][�!&�g�<aT�� �D�f�>$f�]܇ϡY"@�L��pP��*M��?bɛ_�맯U�������.d�Kǝ1R�����͙n��.q%�fi�Qᣖ��z���dp>Y���y�(�Z��05a9��0�r/�{�u�2�@��Ew�&��>�v��3�Ά�����Ke�*e�;?R-����RAl�%���|0�Y"�y��*Я�G���)��6�����t�=i�%iؓ1�Z`�ج(i `:~L4fM�'�S=e������#�*���"as����|���⣧�-��ƲA$��FY�1j�e�Y���0��tS�n�쒪ha�!�
�k�d�uMF{c+֒Ɇff���z �g�ML"yym��6A(�2�5��K�O���ƅK��?��C�=]rLϖ���m]�)؇���� ǉj�(�*������;��<�+e�Y��r6��'N7��I�X���˦�(y�-��tK(��P0�Tw���5�5��σ�
�e�:x�.�Ve9^���ʚ�'�_�P{��¡�7��)����.˔���	�J�0������%!��,����ed5>`���C�1e�ٝh�?<�v���i#��u��=}\,�/\�9��a�#Vx=��&�#$�Py���K\!��K�Dٺ��\*y���>��7��Q�ja�3fP���/�0 QNt�0K����S{yh����:ok�'^�-���ݜC�����Jۢ�?�l]����+z�~�Rʌ/�ro|d�ڈ���;2d��pouX^��U�F�ʝ�
�7�n�B:��s ��.#�Q�7��&:hjx��є��Y�f��B��qfsΎ�J
���rس+��M`�j�-�����,Un[�y���D$���3��;�C+�Q(y���z&���U����?�6��F��H[|��'�/D��qdQ��o�q�{֫P5�{���NKXV��b�Fh�59Tq�y�7 t��|�/bP�JƜ?�h��5Q$I@�?����F����.�Ȼ�rq%¢��tN�b���m�Ȅ�Xڿa�S?�+��?PZ��,����������"��[bP���>�s�ك���h��0��Hz�[�M���I����ƕ c˿{��7N���#��&yo�Փ)
$��B�:�BOǎA�~�d-\��O/f��+�:��e��D�6��O
@[�G`,\_.�v5߹�Ρx|���E�)�(��:pP?�<�5��`(���0�[нg�f�O%�f��~���vl��Wi�u
�8�sdT;ڰ6#�,p���.^I�s�X��w��d:��4���@"�A��F~���(u��Z��2fO�ܝ'�(|�B�~hchM�g�]��6@|�i�WZ\�1�D3B��Da@�F���)0Rt�*fv&h+�Ŀv6);�da������C����NRi�<ϻm��o �f/jt�ے��L����O���q��u����us�"���oS�Gy�J���	8���}�b�(uWO���_>i��&Т��;��IdY����ܥ5�۬*��,�8wz����J��4'Ƨ�9%[�S��I�R�[=Q)�qf��g�Ϭ�d����CO�2650���K�NΧ��,���gx��Hw)�3#��OH	N{X�q���ǒ6�C���K�?lI�z2Üć�I�n����ºM���>�6GD�E�|�4�8�q@�+��g$H=9��<v�e�@��RtJZ�vעp/1��v��KG
M�t�#�a���;q2�3�c���g9���w0ɖj��1d
))к �$�fϔ�YI~_���D�J����Z��6�����}��&�/\#/a6�?f�ؤE����o���w�a
_�Z��"�wm����᪚�
F��L^���*A���2^l�@_VPԏ�8].����*��N���'Rn����P:l��b�p�])��:�J��t�9 iͫ\}�"d�j(jjK�Y���3�w����=�0=��߲�����)x�0�>�*�^��`-�h}�Hܭ!Ju�'��	6��6�(���h�RIu_�}lo6�b���KA��A����l�ڔ�R<��@j���b@2��5Vȑ�:���L4hhD��Ss5��ߵ�M]�T���k��22p���Θ�mo�<�9�SfX��t�܁? ޸�s�U�Z���54-#�f��q�]U9�1�z4��ДI��k�%��^P���^7XQ;�4�~����H���t[�ov,#����-�%�*'�u%�@�`?#[��d�a�M�ԀHyV�����=T�);� �=�i�%٨s3�ו�����;�<l��+�=��?9Lzg�ڒ�⬈�$���&�!x�Aa3偉��ȝ��fP�*S��Nz� ͼ.�X�Xe��<����,�-$D�s����ĩ���ڧb|9t����8�|m��QS������]�.��d�ҠXܚ�� zw%���H�x��2�	4؄� �j��i�w�r��sQX��L�@/<�ا!NF+�ENw4J�~;_UlFizJ���G]�+�!�ߏ�\���6��0�o���U�d7����d&�IC�
�EmiXN eH�"P�ﱩ��f��|���䢯	��3}�CTm�	���e�+L
�V�奇{��8�KQˏk�^�0.ꖏ�S�������Wn�`�)I�s�U�����j��nI�uA�p/Q��MƵ��XI��a#��ER2�x�ЯAS
�*5�@c=$pI�6jE�O{���a�0S���&X����3h�H�-W3��:�ѦZ��k��oUU��Nu��,uԸU�hy?N6`������̂1��
<N�J؛��&��\=�`F������!\��k�|�8�I~���/���'�v��ˌd?.�p|��>c��R!��עK��!?��x��U�#h>t@�����Y8�R֘��Jg��ʨ�����?sx
4��R��*��P@a��M���^�IY�6	��:�Y&^Ӎ[U�'9)cw)��c�(��'�bU}֛�a�lNA�6(06�	�#�!�b��-ո���:%&y�v���M��ˊH��n�qI�F}7�#HMk>(�}�D�=9�u.֡�nipj��3�o��#���g	�v:����v�`�hԟ�,O��ZH�WHM���a����	��z4��kO�W���ʬy+�sr3j�'�(|/���k�M�7��J<zu����sK@�������L��f)m�:P�ƳW�fGļ�v��^�
/���v-�1|k����:o����\�~�/Q�؀	�NIjG.�|��IȥN�B�*�����\����݇# �q��5�۔�p���*��B}�\]�H*�}䚼-T��]++�Lk�3��vȐݏD�?s���W��^�ŠgB�i�k	<���g�/�*1G�d��=sLbu
0Vd/@�sĨ#Q|l$��~��qF'���,����D�c��a�Ij���:�}����\�oVTϙvŏK����vI#E���w�^�WY��C����@�Q���L��MP���vŵ��R/��dN������ ta`)��V>?6M�^�e�m{�g*h��7I�tCx�TE���{�n7���3	��
�6{rs�,�~�|7�(�>��u�����.��޾��/��3��V8��K�P�lŷ$>T�>�u�_���M�Kb���a��索��O1�!�y@�ON?�s"�W�&��? 3p0�{8U�#�I�*�����dZ��]}���E���B\�5e1�Nk��j�i�.o#�X0joB�\�4sō����3����s[;��p �g��\^��c(�ć>�`>?Ya�Ȯ���87SK��ƪ:�9��זW���!e��g?�5�;��sk�Rq��� 7`�1K�[��Aed���!1:��a�%�a�
�H�ۤ���o�����/�������{߱��#���b�]�7�C��m��[�^�i�&�KrZ"gKѨ��Hl�yT,�d`��$Yy�LrL�L��g���S��nm���`O�J!� 5y��U>��F�'链d#+����?ꪷ��6�4��+���gڶhG|c{X�w����l����q����u ��h���<��0�I�ʠ�HX�!�je���߬j^FE���P��������%�*W�s����Q�����BS�9ߍ��5�A��jz����	��,��Xb�YF�$�%�Ngk�e�N���=Wr�^�������{�Y*����5��û0�O*���W��~�;�X�+�03�"�h��d�5'ܼ�{�����`_7d��6�[RXc�a��%}�김a?T3ߢ ���X�\q�A�Q��ׯ���ޖQ��M��Ȉ+����)�|h�<u˴�{��G�پ�­[�_q�~^����NTK7�����9�h@T���nd�b�-6��B�~�I�.�L2�L�U)#`���Ud'�qh1��5��!�v�f�?���ؾ��	�ȇ�М�%�"��b�Ck��s��5�@P����7g�[�LS���&G^׉�i��8T�9A� ;�Ƅ�q�_|#P�{�s+���<��e��L$F�y����I ��@<k	n?��K)��/�y�Ri��n�(��E����d6�J�D��Q� �������zHVג�|���Eb/�, ��S�NC\����(I��H��1�,�s*�DL�0yi��͡h.pr��r�6�q�N��T��N]E��-f����b��Ψ�Ād�`�YZ�%K�I=�z��br7pEv������+l���x����tYēMK�e�����=V�a���M$6.b؄" �������}_�̀Ew6[0tE=@�&�X���r���o��R�����mu��hF����̊q�)�N��{ŭ�&��>�[�ϋ���<��	U����`�	9��s��=�5p�Q[""�fXO$)��|��Mt63�n�����(}-�x�O%un���=���ݷ%jug�V]npM�oĿ�%@H�����[RL+w>U�,�}9�$ۙL�HY�[S``K2�T����n��i�K[&��>�<Ve�V�8�4�&Z��cି�T�]d���L��0�"�c+�:�ٱ�%6#%2Ň)_10}������l����`�N��S�����f�[��9���(%ozP��.���Q�Ȑ$;OA2��e�C:�;�,���
r�~4����d}4QF�~q��ǭ�h�D�H��Y��M@^��E���U�}����ɂ}$К������E`2 �s�'�+j���~.�1Nm_Z��n9)$s��[���������&�b�\c�9V9�Ȑ	D��Yw1�m���w�ڔENU\8��2g󟼄�;cv��E;!��e���D<�}XA�{4�I��~TK"��->�e���}�&�8��q���N���f��_���� %7;fP�Hڃ�RQ�n��c_�Ȅ�|�.Ӆ��qd��(������-�n�?�'H�싲&I��1�Ea�Mښs<�����՞�/����e��^4*r%�wm:���"��h����ՆWAB��I�ch�"�;.Ǉ���T���l�Z+����۝fG�9�1�pVT`���� M��r*P}�:�ʏE��9�%�[A��9���ʗV�G=jS5�a�G�;�^V���x�,�:c���T3"���u��Up���=((? ��!����� �Jٝ�$����p�Ҝ�F��-�f��� ���l������B�f�K*M��tIs$[h�<	�"_�c�JAx�x�=\>ۜ/�JԳ{�g�bJ��Ö������ꜷY��#���^0�@y$�0X6T���p�R��#Zgڶ�'�-�D2V�b��跦\ lj�����_Kް65S#�+��w�Q���� C��0mn"�*�/C�"c���0�"�M������o�hL����3 �E0I�|�P���H�<�h�8Դ�}OR�;��r�|�a�<�č^��Z@��C��	�t����G2��������r7ŊV�&��@	��������#�y���Lq,\�aa
Ļ����z��a���[+{�V�G�w�E���)#h�x~gS1Y���z�,�=��&��m�[�`ۻ�,V/y>�6���7V1���lU3�6�N�\5"ϰ�1�s4�0�dZ��p�8T���ۅ3��a����ME�BZ�W��'dw?>�$>�9z��"�?�=���
� �@�]��\Rav���>������*@O,�Y�ҷv߬����.=��������Qy��&O8{��.����Y�cЍ���G������I^��"1��i�.��{$�Df���rg�#��%&{bu�8Tq�ު�&`�:7���Ҹ�6�4�>E!L�s/����Nk�!�\__p�R���.'�暠�~�%}�7�n�G��d� V�b�Y��#���LR�P��p8h�S�Wz�����)��}���+���X� ���K5&�߆����7����xT�G�Q�[I��b��WF٣h�F�nC����|������jB�x6�PA���J�W=�sj� _��t�g�zm%s^)wK�27���~��>";�R������.���㺰xf�Y	)Q+�=�@1�9?i|1�n.n�]]N�H�y������IM������q��w���l�Kc�c�6/�:T���?���q k��R��X�a�e%�A��6�zC�
��N��%� ���p!5m�& ԰�S���oi�*���aK������bi@ۑ�;�P3��E=3��~�{���1���+xU?��s���5S�>��D����� lV(�N�ﺱyo�U|zd{ʨ��d�ƫ�s]��@��N�:�@A�{)X\Z� DI5��>�]W��U���Gp�J@q�&����;!9�&2�g��P?�4��ء�;���c�{�>b5@�e�D#�!"V K}�R�^�b��m�!!�N�o�����nSLE����d6�2��_U�E7�m��:��X�*��B�. V?l�><�1p�%��W�.K�?dV�;e�r4|�*N�$�Bxga�-f�ҥV�ߛ�Ý�����8�Y�j����u��;��)�ތ��Ț��K(�$K"7�Ȇ|GO�07ƕ�v^��@����mq)�B�-� g�>1�D���Φ�w��M0H�k�a� э	�c!+���;��������p3<�f�����m�%yoD���>##[�^R#xG_w	�>��&�ϋ:�o�Y�Ӂ_Yb�=}�6�;�y��=O1EU�iQC���Y����)�O�V�SڝqӤ�v�" v�6�gAoF�(F\j�����t��(*��������+��+`i<�[�O�6�H��i�·�hR��H{�����H�@Cd�~�>�M��;��ܠ�5��:��`uH주\��Ϋ�#T�9@<7-���+�"+ J����-�FQ9t�q�CL�}|.�V
�aSe)�^�,_����.[2�;�N[	@�ޒO��?��
��P�|�x6?������_�D7��_�1��q.\��f�B&���C�T�Ilռ���2�3���ᅃzv,��l���n��r^�z����h�&�YiC^��4a�J<����)�%�N��G�$%�<�9nϹ�:����59$��;�:�r�w��3u��J��M��SDV�Q�4���.�*y4����^�K��C�����$�3Mc���Cy풓�#��~��/[C�0��X�'i��͑(=i�k'�0d
s�IK���q�*���.�W���&�#O���N������Ջ�ƛ����[xmYd|N|��j)A�k�tՃ\���χ�-&֏�f��}����`�]�į����Y��r���k�����f��&󇭠�/x�L��a�9_�ď:�q�aA���E��}l�7	��}�������[8�:vA`R������U�N��;қ��?0�w ���f���� ӕZ��`�@}bm�c$Լx�4r����R�Bk}��C��Vl�
�ĺaF#��P:�s|����:4�B|i{C	����ݑ6!]�U*��kABJW�Z׽�+�HlƉ�g��Ll��w����@��UE�Qw'�$öU�+3"Q�BY��2��@��B�6(
��>���m�`�=�0j+J��@P"��d�oɿ4�I����R�3�WRbP�h�@�S� |��6��5mV:v�sڰyk��f�b�9A����@��k�ې�٣|Ͻ�z�f~Z����f��Y�Y#��	*1w^.	iL�~�og�Ȉ�k?]u6PD�&/.�ތ��IU`>�~�i��zi�[��:�|{�ҰiOL r'A/`�"�Pè���@��=��ƛ�'��{J��

�a>��c�p���Z�n�	_�ՅX&��j��2�r\�Iu��hd'�w������&�o�jA�}/�SJ4�巀�������]�j=g�(*�D}�+�f#�aݓ�ҋ����S	vu��N1�	Ƥ�oz]���*�:�b�l�[?6"}�lnJPJרD��B� ��}j��{'�0�
İ~��
�Qʧ�����x�]�/��[`9�|�%�Z�����ox�E��A�� ��%��HF���ж�j�8�7^<(���l�0�L��,q����ڮ�
Qu������d8����tF��XA��?�^z��b�N3��)��!�yF�Z#���~u�}^@e��>�ykf_��듷����7S-�欀4�wX�r��B���5؟��Z��X�p��|r_Y��Xv��2k8Uԡv4rI�>L��,�)�B�K1X��|ݗ))ٷ[�V�)/��� �!����,�%����0��mh&Աǯ�@�
@����A�fl����
�B܅�ǃ���&�[�����[�C�)�3�Ps�`w��i�T������T�\�B�_e��Ț�s�6B���!k���>I`����#��O�Np@�H�O	DRbS"�ϡ�1|yɏ"&�#p�N�	(��!t�yQ�u��DD`Q�9!
��X�ΊDh�n��?����{ϳ�p�lX�%煘��R?�׷FHu�8�G=�$/p��}�Ϫ�ZW/�;`o��%��������[� �ɿ����Y��:��Cj�Y�בn-��ҋx!ɠ'3j�R�$���f��AO��#a�B��/Ee��	�(z�y��X���0����*�J��2����.o�y�R	�u��'��3��\έ���	��d�EC�f��Nk3W� >�ha�(i��P������θ��$�siK�/���F���Z��eĴX¥���{�[>��f�GH����&�Cp7�f���DCˠ�^2��������XeS����6QJq�
8�?<����+-έU�Z�4�"�}�1 ���/,	B�����V@�[W���:��t�}�/&�
�4$E������YfA]������V�l<�%NՍ�t�S�*y�,|�p�|�ᐸ-Bj�!#
t0��cb�hs���3H���'"�)qz�0ԙ�z�6+�0c'�P"j��	G�j��7>��o^����!Wl{�/�b�y�i��{H��;T���)�T�$zI���4_���>���)lʄ�H( ��۬�$MS�J�@���W┕����h�
"�Q ����/U�gn�]͈i�~���hrx+��a[�^@��8���[�4���x>�߹��רf������m�o$x.�e�KJ=�O˳,�����z�Y�Mل���4��� ꑊ��� 0��k�gي~U�ۑŖ�%:rQ��Wi�l`IQ�U�*�I���1��Gg��0��N �9�R=00"kz�	I����b���r��M]�ɯ��ܜ��'\��� ��� Ȧ��5�<?n<��cT���r�%}6���N�e�2}�k:,�)$6aryA�����˽�I�\����vp,)�x襕w��/1���%8;F�N��IC�֕D /'���@�M?�I�4�����f놈�D��q�IS�=����w���T��� �����e�S3`��j>�y��O�u� W3H����x�'K���޶�%ixr�S2�ٴ�	:A�=Ǚ��*'F�R�&��vɂ�bA&�"��:9��"�3�7�@8�cB�hc��f<���ޠ��zϨ����Q��h��'�
�e=!����G_G�J9���1AV���p7(@��}��
)(h(�X�ulGZ2�1Q}TvAZ9�#ķ�W0�����|��N�ֱ�e�e{3"� �i;���r��F0H]� G�Y/D�Ǩ$#��e�8���stǛņ2$�� �Yk,k�D(֤Y�FWt�z�椺E��Ň�8�h��]{�.�^�� �d`��^M^�c�é]Wqr����-I*��� ����/7k5<'�#���X%�l|e�e@�ҥT��5�]�8�E��VW�8�;k�_�O��l�	��k��<����-T�Ӱلĉ����Gi���o��Qr(�5� g��=%���U��v� �N��Ϊ��_XC
��C�S7�*��<���&'�|x��7�~�jn��i�.l��m�p�oQ�F	|J��_�ͺ&+{��!��b.1foW�i�������r��	����ؾ3��%��������$�!�Ȃ)=��m9!�ňު�aP�)�������LJI""�E�k�g.��lq#ؼ�K�!����}��q���mgM��o���x#5o��� ��g��ʢ�C)�|��Hb���/�Č���c����WW�p�c�|��wɝ�א�L';�m3v&3�H絻C3!��+��.�X����2ʓ�?5���B��4 ��RO��҉qڷ��i�	͐�cP�a�Y�]R����Y
�O��)��2�(����f�7L���a��Oq�t%|��Y�O���� 0,&���DO��|�f�#������T�,n/sX�Z���={��̽����/��?�<z����Q�j���L=�)�h���ks��_
�fxy:}Ԭ�ac��n�w.�*%�x�8�bK���-�3�ב!��sy�M�uw~b]���i��1�Յ�T�s�����u~�;>c@�� l����7����qy�����v,���|/�����ڋ����T�lo�O�9g��H���r�hD\q�Y�v'�Ԗ�xRq�L/ME��G�Я _	�N�j��g��9���kT)z�	Ԥ��d�4cinb��^�ڹD�!�#���6>��_��#�)� 2h�;AO@n��{�-�JB��?,��r"Пy����[�����ud�vH��QNB�����oV�=5D,2�,�8��efU��-Mi���q���޲I�����ۀx+P� �����p+r� ���Q���c4GA���j��4���e�]_�6F�3eGĀ�w�?;�.:J��Z��
�h�4�&?������}3����� @z�u�D`N��k�F�/�����q>�,�qs�:�h��\%� �fb�O�dr�)L^	y�])�i�������`^	ض��"�F�pҏ�ϭ�6����5��z��+��J978���!�X��ym�������Y[@�����t7_���F��SԜo���%)l��6������+���&� b���#�کAz |Æd�)�̭K�Z]�Y8O��=����ET�G��s�܉�<ggT��8΅����U�X&PZ���g���g�P\��xG3*�#�ϫe]mg�~��"E�g�MRI`��;�)������Ծ�ڏj�9_������8��[z�e�G��,��Q�<T.�1��sG�'��~�o�F�ڋa�0�q�(Rkw��q~��Y�H�}���u$#��%/3�Ž=��}I�D׵f�iox�����}K���D�SHt|:!j:zm+xm��6�M��������=�b�nX���/"X�R�}W��F@��T+"��+�{��JuY�(�3!O
�F
u`���ǆ򠺸ağ�kI݀'|�0*��D*zN�Y�K�����o�ʦf����;{u�֐�N��r����q��&i��) 0����]�nr���}�1�t���~��.@40�X��mA�.�@��X���	�������	(��^�#1,nm�Ř�8�
�bO1*.�����"f��π��~w���Ơ�h}w/=*�a��w|cש!���Ș̥�P��2?���w��d���#��3����V+:ID�$kfׯY����6i�{�AD���t��6�r���TBF����R��D�;r�I�)���V��N��fO�NT�mG,��3XC@o5fD��0Ms�i���MҬ?D-k&��h����*�0�m�");��*�9���jk;���2f�(�Ѱ$�`�ÓK��GH=�z�*V�%	�08�4�� ��`wfj�I^�j0A�Fk�����B���翱F�]��(����)U�o.H�&��B��y��L��[�j��dZ4<3T�>�Vm(y<.uQ��P��M���ٞ��s�GsݥB�4�|��O3y�E}LX��<��J��ҥ��ٿ7h��[��2q /���C��{�-����Y5��HJ��XL���4��
��F�����b��	��y������\��2Z�{Q���H��]��DFXbj?�gA��p� ֍DF�Yi��~��%����~r�D��a��)ю���s������'k�cqr���%��S*�N5�k�h� �u0�l�H8�h�,�l�$]���S��K�oZH�t �R&�������Re�%:�U5�Q=\40����@�gPU�\��P�`�sT����rY�X�G��LOu�oc�.���%|7�������_0�1����e�|�} �gD���zGqE�$��j�U�cT��|E��fS>�U.���*5��9�h]C-�(����	,������ ����<��i���&�G�j��*~�8WM�L��u3&[a�ZS[�2�zj슺Y팜��Vɘ?XJ���H!��FzE���:Rb��+��_� "Z�A�V�"Z� ��#��HaJ^�Nϓ�4Dvn<��w�Ӭj�����G3[�a�Y��E��s����_#�,���"��iX�?%�K�Ԡ3��R6Ae�P}�x� p.��s��j�p�aʣ4�v�֋��MF� �EF�S���w�p
'_}�e�)�
�d	Z�#��y3��3-HB���?��<������1�U`Lgŗt�>����ZȦIM+ڙ�=�M8�o6��cP\�|Kx�[���\z%.@�*k
���|�4�Wʮ�;�&��7+�o�!���ޯ�+����B�4����ݹ;��߂1��V)��JDm��}�ao�ª  ���)y���;�/Fm4�D*�^1�l�,Hq��?�}-P�= Sv�!�1�u�[��A�g�v p��!-Zш�O��@n��{:
��3P��8�nK�Υ�l����ӵ���HU�)��e#���y���������_& ��q6#�M'��3NQ�Jp��� ��E[젪.K�]W;=������@��U:������i����_4;}]^O�����Iu|M�����D�ړK0]��9�(w�C����yUh��6Cw���?����q����	�c}-O~��.nx"�L�W�����/|�%�1�im��K���Đ�k����'�N���n߼W"����+��������d�@���zY]�A5ʦ5��&y��V�ҟ�Ծ����c�KC!�Uv�Kj7urC�����0%C�n�,�@�]�v�Lz%�X��x�IH,����f]���^�	�ŰP��٩A��Q�Oˏ�W��K�3���z�V�tZԃ�úb5 @���bZ��!�2Js�y�;[�Va�7�+�| 4LW�N�~��D#��s�{�V�2�ϱo65��q\P��ψ�^��x-ֻ�M���o�"�zv@�,��n'A�����N��/�EZ1|���f]� ̉=��oa1���ܒ(�T�>B�u�'�ҏ�T���VEN�c�1�Ѧ�u���ʸ���'����y�ў[�'���J97 ���g�c�o#�ڐ��|��jq�{��LGqM\��D~�49A�f��p�L1����p�l+$e���s����ܿ���b��ƅ��$|�����KMVEy����kT�]��n�>[\Fɢ��$!��e��:�K�*��%�_9gI3K�cs�۹F��{���������$Y}~�o��_H3Si���">U,�Y
����e48�Ik�W<�����7��f�1ۏ^Y����ךV�hrH�!W
�I��4dø��x{]�AY`��/ǋ�Ha�f�.��ӗR\��8NY|��L�h�熳���.�ԷL�����#�M@��K�J0mq�¬���/u5�=Wt�{ �� \̈́����N���k`%X�#}�- �=��0������揵R�'����^�@Q�#S��e�/���N�l�cn�Z�D�5�WCW����򸷷�,�2(�r����Or��9�M~~�*?;��O�!1(���I]'.�>�ukR�P� C����v �X�Q��O��%_륣D����=�儜.S�4�^��QeN��X�W�<Ķh�P�����̵�B"�2��Y	�.ER^��HaUgƬW� �o�V���Ǯ4�.0��O�.���>���Y��&�D�E�?D6�2� y����ͼ�ӊŖ�B(jW
���+o������+��z����C-��;}��-�,�<�P���$��PDD�;���=U�//�և��[Ge����h2�OI�2���kR��3|�w��/K~/VZE-�>K��m�EOlc�?/�@M�v7��"e�C�!�4JSu�p������I��[�/��ḇz����J����w�ߙWW,u"~���mh
=l�8H��,4(+�4��o�m���P/F4��i"�n��2$D�ؖj�dQ&U��@�o�*�=ڳCi����D���^��ټ#M�sT>{���Xm��z`�6W;=����3��pç�����	B�7]���`�zȟ�����[�˝xAh]g�	}�SKS��	ͤ�`������|�aFS���9ҐO�@E��t�f6��J4�ga�cC���e�+�U��Q�T��֎��	���V��x��6�[gKI C�c\6�#v���15P^��_��Fc,�p+?�1���S�:�����Jo�ġ������?�p v�wQ��3C�w�7��+m/dtrƕJ��\xȾ8��#et}%���g.�ǨTus-�vФ��"�	Ei��}�q�������>�ҕ f�M8�$�O�^��
1]�T��nD�����
�'�sp527.U�G|����n?�e��Q�rr6k^]�+̠g�gtr���6�����O��A���<%9����ށТU]���3���ۧ���~ ����U�2Kv�zR�����?�H:}J8��銏�����X���b֦0v�I�[�L��X���:���E6�F�����Q�F[~��&�8|z����H���vfk]���z+c�����������?O�"{4��_&RX`��=�4����|�A2h���~5�5��ՂD���Z�GDR��z[	����#W��[�5>����z��/ް�l�� ,2�h�r+p��+�Q��b��h��E�t��?���֊ؐ.�Aus���'��2���Y�/��U�}@J��<��*#�MNC��Z�=8��]�	6Jt[Ǉ�E834��]�������/N����.��
1�_�@��eZr�9V�P��G�x��*T�2u��'�� xa��xՀSv�����kxB%����.�e��_�1�����xL���֌�\H��Ȭ�N�N�d^���'�����q\G�i'�ޤ����ql~���]#��K}�C�vd5�m�m��f�i0_gUu��%?�X��b� �m�$�����̶��~����B*
 ���c���0���s�M��`J�}���5����N�K���Xy�n��w/�-e�ϟA��cv��
����co�z/�9m��v��m���0��;�|ʉ�AFRDu�H�m�����%Rr|�g�b$�95�:Ll~a���p-{+s�v%��=�=��
Ae�5��x�^Ըϔ���T.����H�vg���o���χ��u ���r�!r&Ĕ ��̈��g�7߈-���m����|��L��	�~Pqۙ{d��YcF����Pk�'
*��/�?���e�ρ���AE@�~��{���ZSS,�)��p�.���[� {�斔�3�:�|����MC�W�'Ue��F��S��1} ��P�@�8�<ĩ��:L��Ӎ6��J��ųÑ�T,���w�ה\!B0t�/�?z`���}	����R�����h
)k� W0U��M+�b�$�q�r8�0�7H5����5�u��s��Y�?�B��W#/F��+�eH��ﲷZ�� w�e>�Pu�Ƌ��){Z���3MF�Ju�r4�c�����1��K�7�)�����h-����8�����[��n��5i�;�����n�C�<�N�Wg�A���j�߿��$�b�3S���|�r
g��_�-5Z�/��h+>���<��K�q6��(�w
^�Չ0��pL�<$nYc�9�J*nU��N#�
�@���UD|����vȢW0�n�v��ԇ����n�I��M~�?}>�昩�\Nm"J� �����H�}����A�p�~bv���I�~��^:j:�QL"X����	tt�%���Y Ms�8?��@�{�|��\�c�/X!�5�d[�+3~�b��'��H�q�'����>ҍ:���>����\��j��X\����,+�n�`�R"h��W���3��-A��\%��p��IH�>���6��ā&a��0��nP�gNՃo;��QS2D��c&���Ll��aO�i� w}-ocVZ���f9O�Q]Nq�!�~�@�@�^-�*��$%v��j�0i���'���ꌚt@�i�Eږ�hl7��P/���V���E_��"����7
<TFIܳ	�\M�I�Z��i��.?����t�a�u{��ře8�x��dV@b`�1���4�9,�o�u�#h���,A�b�m������}>橇���jy���"} A�Sȵ/(`}%ׇ��3Jp Ug�}�����M;���B��joݬ�ڣ�Ґ�/r�}m��x�%��6�K�~]YO�pf�x����k��� t��]�BQ�'���A��sB� �/�[�d��q'��D����S�̴���qG>�j C�`��t��ؓ�f��`)̪��Hp��L��+��Ķ�%�������so�5i��߇�S��4��!gM$�m#�x��1�B����Y)S�I��i�+p���]Q��7H���*��]P'��Y�����6W$��[K��Md���;�~�S�w��/�B_���*�@������ؔ�Ǆ��Dά'�j���@���T�[�r������ts��H��u��Ja��?I=M�#�4�we*E�(���~J?�%�-2��-�q�Ǹ��ɾZ+��j��mUv:�Ot�����n�׬��\���Q����a�6��E��<���q���|^�"�̽���I`�a3�Ė)7?2���О��i\FtQZ/	9��r�YCn1���DmJz���*Ilx%�­�􍄅+�F�M淒G�K�O����h촪K��<�ؖWZ��}��f
��[;��{����;0�ßU��n4ι�C�����kT~Q��)�7��n��)qB�c}���0�e�߇5�q^���v���7dbM�`8�Y��a�꫱R�&���i�l96u� �����I���N��aA2��-L+������n�'!�+ٯ�~��"�V	��O�9��s�@\�KǤ�	�+��f��b-8�`��_�p�G��v8���J��q�B��a����N��׼� ���s��x�߹������~�M�-� ��D)R\~���LI/p?�����Eyڊ�7�Odɦ[yP���Z�d~�*���SPB]�S��%�[5����7��p�C_����z�� H����K�����w.]m�Ϲ�8�L��I|���nCdLQ��������胐�x�'����D�d��M}Z��r����z�fP��V@酾mָ����=�_����3�SV��q}�������rY��wgD&{�OL��iĚc�[E+~0�y�r]�7PF���C�����sD��@g0������w^d,��Be�"�����(�H�-J��$}zj�ʣ���Ľu��Y�O�\���ܹe�]�N[�
�C�Gy�I#uV�w��#K����a_V��x8j�_�)��E��﷛�䠸p��2a���Z�XcB�t�/.'�"،&�(V��\6s���2c�x�:�`?�e�*�~��!A�Y�}�%t@�8�����-���uj�1���>e~����� ͇_άi� @�w8�����B�8 UU'*ģ���dXVz�IIg��,�^B�.�SQ|`��al�j?���\��w���!'��T�^e����c���Xx�݇�S�r�ӟ΁cm8?e)�n�\��ܹ��<Ĝ� .H|��X�H�ڒ�f��Q��cD��}0����� ;��^��,�=��y�x1���E�Ŧ�}�]⊽!���8b�'B.<p��ғPl�@�ݾ�2��'�k�Η���Z*��'��v�"��i����2���	�d�$��M2����aL�L�z$1I��/C�c]�-�Ｌ�ߨ*% ]홽.P�A#K N�y��ۮ��R��e�K��`����̼��(�L�H�Ex%�$���)�\�:�vo�z���Jg�GfC�M؎�d��#)����a���%�Ż?��iY��3��8o�%�.��W�OEt5�B�4B���,A�T�z�>7��"?�5�e�l�L�xǤ��2�IJƅ�)w���N�xB�T�b�i�v{���*���AK�}�Pϔ�������vHoPs`�S�-u��*9^d�,d��X����a�xI�]��� ex��-�}��: ��q�ݦ�72�� �n`M��ڿ`}DՀ�~R¥�i������M�C^
eꚻj�'��<��J��Tf�a���CF��I�S2Oɋ���k6�v�S!����}'#Q�w?���z��剄-����7��E&M��`i�D�""���:�U�q�	;�Lm�Xc��"��$�^���C�XKo�:b����Ey| �۝�iW�ob����>1����cK��D�Tf��(�"���� t�em���"���j�{�x)czh\�A-M��Ƿ�:՗=o�b�ms��Z+�=�x3&5�&��ҭ������3�+A�T/_��Gi7 d{
D�"�W����%�XF�qh�w�0��3�X��2Z�u1�M�Y�6F��)%�tE�p*�@�����G%���S�KBW ް�;�[}��,E2�(`�����e�!-� �����ZD�"Q��Mc0�5���j�E���_�u���g xJ��F�_	8�y+�fY��]�ۯ+\������\d��쏥֊Z���3ٞ�T0sb�&���-0eyuПR�j��ݸJ+�ɢ7� ����6��q���v]s�t�Sd��sm�s*��hϣ���T6��(�c�}�y�N*1�ؿ �PbK!\�ߵ�D�t�������5�:[�a~��>Kr��H�4d��(i_K����7���m�W��3�4ٌ��ha�b�^H�`�U~����(�W6%��
��â�	(�~a��b�:Q�f��m4����b���N��NY���󙣇*��H�����Zj�|���ͤ���6/t��ӟ���/��a�l��p��7�����8�v"��t��'k�4.:�����iߛ�5��߭�̱�NT��#>�Ey��M�ֲ��Y��<�:(�3w�:�Y���F�iD	��KnQί���L#x��:����L�+�@qپ��H���6�@[j�g�Ò;�Q�;\˹��oM`�_�,T���B6������X� W2&Z�`��S�)ALxr�	��gG�1�L�zs��h����%^�.�B4��*���5?�f���L;,�k$n��籢L���l�r�����/{�HA��V�E�h��x���y�X��B��Xf���s���%.��ڞ�5C��!�����tu�Ս^k&���������a>"�� Yh��V���<�EW�&�V�'��2(_����^iq�U<�+;�Ty��ɶ�P'=.�k�<�`D�7n�>n��d���{�H��h��E�ͭ
�o����HU�%N{�y�$� � 1ك��-s���QG����~��dB�mc�vr{u�
��)HT�C�j��-ц�n���R�a�c�����p��m�6���Z]?/�"<��qo#��$�f����0�EF���	x~��z��2ua�� �����*Ӻ�M����҅�T��ω�r�1��L�'="���<m&QH��N��v��yt7m;+ �h��?��f|(�� 4��X�o�Y���v�)Ǜ����
��K^D��������Э���V�i��Ӱ/>�ce�����f��z"`��$wd���.�����z҆�w\"�/L�r����k9Z��C,���Leg=��Q�U~I(�n��=��
�K���A�'�Y�4��2�G�I����]P��c"��������.n�����#_I-���2������)�f]��~�{&}�{]���~��A�����{1;$��=B���X���>7pK=�M'�P�Ȓvx�,S"GTV<= g�s���e��JS���������-�V.-	t�M�۫�>5�"�¯�h*�.��	p+˔-�]8֕��i��E���Ws�v1�-�6��j�j����X�o�J�L]m�����/gO�F��0� .p%#���2���[ƉH�7\A*f�'|�Kko<h�Q����^wN�[�H�����|N����vHqw,����\�F�Vs?�.~y)�Vn�a�L�1Zַ��tC�8�Q�L�H>���(����4R�)b_��!�A,D�A}0�{���H�8��@�[=Mr@I��1�J�,��|5�"l��z`�1}���ˌ|Ǜ�u#+�U�]JXР�C7������h.C�^Q�����ιp!?{��쳓 c=@?Al�S�2�-����6o���Vq)(}�^���eB�����r(B9����9A5SP����O �ğ �G�H:.�a���|���8}v�[;c�$)�k����V��@�8��T����ĉ�݅H��BJ���`(m�c�?��{rW�7E#uۭ	������~!��Q�����"a��fh꺜`#"�@l��o٨a�V:�J�r!C�p ���c���X��Qt���\�HG�p���pb1Xk�NU���[��`@��0jy·,�;�멑-�-^�F�r��9���t���֍������5��vz����W_�V��՗d#R�0}���(P^��ݪ���?s(����t+ӵŀ�����9��I>W���M���㋐�+������Ȃ�~����b�={d�o�y�`�6^��ɺ���/�k�S�W����#�7�}t�<�����ҿ�n������Ƀ�;�,p��i���z����(l�)nVe��M]߹������q��BR,��ݣm��n�*�%-��iS��Rm�5���H/6��3���s]��{����^W��a��c.��19�cs�F�y&@����8��y�(#�	�k�Bg�u����h�NH�5Q�6��38���D5���[������o�������U|�L�]�֖{~�2�Y0�9�.�'d'`���j6x��)��-��-rI40�	�������W|�X�?ŵ��x� )~M���g��F�\�S��K%Ѿ
��O@m�b{�Ӂ��$�k��gQ02�uK��ёC�}���y;*|֘���2��$�,gY٬����C�>ި���yp�_&*�v|TK2j���頀�3�V��'A�}@&�p*�V�/Bm��Hc�a`�4�h�����#ˉI� {^�YI��	U�闖~�aU��"�N��*>��62���p���z�F�\U{477_�Rf�S�)��7k�U�,#!��s�d�{a@[��\��1�~�Đ���f�W?���� }�Yg�Bs�s��	Czmx�ޡk��	��P�R!N�����2�3>�D�"֜P�	e���΄�G^���3|`S��x�ԕ�	���^Mq��ƙȤn+�)A���}V��$AA���d @���4|��>us����{�|2&�a�����NAړ�����'S-n��٣��3�E�����aN�%��W��HQڴ�兽��C$�5��u;��1�LR�fuʍ����K�����|�j�ɵ��mS���xV��l��m��G��oK��b�����#���i�"f���u��yCh^�+=Ve����n�M�|g��q"���pX-�������w��Tn�����S3~ ��X7y�_�����`���=�5�oh���6����ʣ�N��fl:�bz��w�g� �	���O���K���aE��#�k��x�
�u��k�͌1��L`�_G��O?�������	��"RO��O������,��Akܿؿ�M��^ѕ�0����}u=D�6w�3W�1�	DK�?W�JJA���6T>S��Ͳm�ꑎ�a���9�K�_3���X�ڴ5;����Y�[����(Uv7���cΔ����ol��e�p6��T2p�ͻ�p��4 &%��{{�ߴ�D�C�e܍�T�ב�uo��+�і\164q<�.���Cj�����D