��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	������&�RS�����c�I�����`�OiM��ި��-���	�6-�l�n8*�l>A�����+`�CاZbC7��ł?h��6�ņ=*�C"���)m/yk�GM$�V�]�Z��qs1Y7�s.5��D�< ���*��ʬ�16�d�F��M<�o�1&���:�vj�m~�w�����n��_Vmm�X �I����Bn>E'��'����0�����bv�blן�]	;}�!�|th�����K`f�uȝ�y�Ivo�@�	���d5ٌh*�l����&1�Lt�aD���O��F����~��������[e\N����Ͻƫc���Ђ���1�7�$���k��?�T@�_�t$�b�DA'�7�~���y���!���a�x�0�+�s�� ��Y�����%�&��`�)�Ôt+B��3̊%ZB���L=��	��GcDI�|e�n�FK�;A���T�����E'@��i�y�=� ��j�*I8��`={/w������g�Ŏ�}MHԩ�4�\l`��#1���^���cT�7�<�ٌ925?����XT��~`H{���&��1��ȶ���_� L�n�,|�rZ^�22�����W�y���2u�	����t�cտ{�/�"�c62�"4��_(j��~|#H�[�x�&�=]n���u5im�UX����ò�{�bI��K�t"��3.�(/@)&�.ЧE���<B|P��4J~��7Ԏ���YRGJ�&��6���x$�31���m�CS���׉����"H��Ds6�p6�^�m�����E��%�}���Le1�$��h�4B��3����㌍�<��z�����
H$��@f��F,�V�C�܈k�u�4�PXc�4ts������D5�I�@�֚���� �f�g� |1�Vu�h9ȸk��A����0�? d�Y����XX�\���:���B��3&�n��<�eD�l�R� �ƵVDЃM�ޚ%0#咐[CiEϟh=^�:�d�詧ꦦx:?IO����pZ�% ]*��b���}&_lb��`��>u�C)e�I?&]��]tM����䣱���v�H
!���
~�(卲�gKiВt!��M��Ā��m�ݼl(�/�]T��mA�#yi�w�����:M.tZu���prϺ��J����bDX8��v��Us>���-��O�G�ȣE~A�8ط�I� �2XhP����.v�a\%�Aބ#�x��U����;�E�Ee2��jp��x�"y�ab�r�� F&4V����j��,�4�=���d֎�0��i��B�=�&aE�,�"����ÔF����n	w��PcޑG[̘vt��խ�nO���GH��l�zz�^�\���������\��͗3͟ F/3ef݊�X������
�pe�ԟ�4�u3�˪5�<�4$=uE��l���/չ�s�Mn��%A��&Hc�c�Ui��q�Y�=J��SC#nX���2��36U�ۖ���<́��u�Q-W�r,Fp�H�b�������.�z�J�����ue��i�QEȗ26��w�gGi�6�nYy��3U�uhm�l��N��e��P�)4h��C�T2�z���d�k�e߉94s�e 
2��S��:M�_Wz C%g�7%U����'�O
6A{}��9%�â=�|t�S��xO�m���W�h/oѷl����1���M6<x6���\��ǁ�[!��#�� �*�`�M8��"�O��#if�K-:��k�>��#w��5s�LX�L!��{$��Aꡏ���.���&�:z�TW��7�{��h�z�O�����aǺ/�V��w�D�33����܋\d����y2�+f�
�7@I47�z��)n��+f�2��o��8����ry�\�W (]����Nm��+^4�Wr�~7�"�t&4��j��;��o�H�S����\Hx��J*�w=�b>�/��2s�ݘ;w.�釈�?�rG��Da��}�Q��������Z��?�����+�d$��	�5�E< 8�dR�%��csٚ�4����&V�S�
Zh����	��:k^A��ŕ-�����݉Zrt/�)A=��9�Q`��5�����$���}( L/�3�"߬�(B����}���]�����/*iI����� n�!E%��7���Հ�W1�\U�Pauv-�u����,.���ʈ�����;������ݙ�w���i/#���9������Ubc��:Z��V�9,z	�&��2A$1� �ηhϦ�E�U� �����WߗQ��Y�%��i��������@�"7R�7Q8��3 �l>w�!�'
|�ՖkQdƏf����f?��znӫ`vS�����?HbkO�l~T��{ɼ��$�xkԹ晴���R@]��:h=�l9�o */�7Y]$PY���WP�����wh�b�����Cr�7*�$IH�2H��~���y��ʽ�v����=e<TDc(%
'����M�n*���h�ݲ����f�"�WJ��4��WPv���Zh�p�ȴ� �u��Y��Q���V!�1�8j����[����-��tL�+%��^��YPs���8�r���K��3���
N���x������}���_ܥh����U����z�����m-DGƅ׼��,��0Ov��=Cz�3/e^<�=�g@�#��|�bO˅�0w��q��*a�t���N�Əj��T�-9cQ��5�i1�m3�Y�j4t�U
H���:����'�LՁ�b<�F�0��)m�|yf0��[�;�|�]9�H3pq���d��b���`
�#����ٮ��Zp�9�QY��G�?'��EA'k{T
� .PD��e�R��9H�2�[]�_	�Y{�w��R�[B;�j�s��K��@���)��O��@Ы~m�F;(ܢ.���Ae���c�3Z��[�6�>�n}�e�ދa)C�
�u����6<�'ŉ��H�rB�MF�%q�S�Q�7Rb8$���,"^IkU��=Q��Ù�;!mv�ݨ�/���P2]�]�i3�x<�E4��h}�[O��Mj �I���ut�"Ne��E*xj,�ZG8��b�o��ݣA�骐�}<w��0#�R2oV�c̽���f��y�`������o��_�8��E���E8F&��9F�μ����BN.��֜�����W�����a��&�"����s )�)1jbR�H����.9*(/�y8��)�)��C�f�E�)"	$�����{5ͅ�	I�jTN�`�E�U��V�Q� �F=z�(���h'!�_G�@���;��\L�Ah�FJ+DA������7/v3uA*�ҧy�#n��V�e��o8��Xp�!}�-�9�@�ӡ�-��;6�Ū�d9n���{�𕤉!��B?�1݇OFAh+�\���)bRL���mB��`Uo�Yhh��H��y�㟙 ��㨡2G"�����rYș3o�>eܪ�����|ob+�ܲה����)���o��������y� K9�>N��g�Ͷ9D���ݖ3Bv"�(�f�\�h���ۯ�2����؈
#�v��ljq����_����QK�%>C��� ��PGT��E�{�Ł~Pw@ �8�5�[,�4鷅S��N���%�&uMO<�,� ���?7ti�gI�K�y6�"��*en��{��Y�&�V�5B�rYΊ���݅{)9��_'��>S��
��&��Wdy���>�1�x��G�]��=��:��O��4�
�_��ͥ���w�6c'���3��3f�����@�Miv���-�̢�ٶ�L�z��e��6�Q���
�B��L��b��Y��h�y��_�h��c�����9�;q>4�+/�Ǉ
Z���"�̀Sk͢��ٖ6�������}���Hb�:��&�9a������٬Ns�/37��@ ���p۸����M@`����u"�:���/��������7%���I���b�U������66H%	Xv��C]�A�/ro����&ɪu���B�E��W�E��=)k���1�pt�W��
i��V�,(��LU�m#AV�;�FDr�����Fw����_1,����z+�2����%4�J�{����۔>�����/iS�!�=���,�$�ޑ�~��U��.*��a/ϾxD6Xה"4hS����]l�0����k$ל"u�o�ύH���C��	x'�iL�P��w�Lz�DHb
��siBwn*3��8�pst@��J��~S�8@����-»�;s�[\G��� H�,b��;I!a�'���?�Xe�CW�c��-\�{��Ȑ���!�z����b]�� V|�R)kL�)��v�q�!�&v<�O>������5y�z4G��>97x��T�ڮ+mb�J��'#���@y�{K�/@X�����ړ��ec��z��7��`�����@�"�Q��<2��9t�����Ē� ?G�pi�&�a�;$v������A��:�㮰MD&1�����kь.��Xu�Im�m=�2|��^��p�Gj���ߔ3�9[������"�_~w
��!"*���h	��_{�ˌAS��GY�!tzʨb����M�-S�r]F�� w`hB��$��Ivc�n�
�r�h��!_�J��6Z�Q{̂��jܝ�sk�&�&:r�4�%�:�~0���]wALȃj�����I#���Z�-w�סM�Z�+��F�l����@Y@P�������bU����K�%�jU��Ra6k�x�jc�*Y�Z�L��{&�fˠ0ָ-�V7M�8�����lz�Eey��ҧ���z�'Kr�;f�aW�!�m��Pu��x�ߑ^��>���q:�o%2�7`Tt����9ɪ6�	���N���l�w~���C���V$���k*D�q��,v���`��
�Ѭ�������$x=�g<ϵ.��#Ԋ����,P�Qҩ�ホ��Mo���.AB�S.�-`��j Z0�օ�݉�- x�`�OO�}A��*��֛��Yz	F��@��"��Z���\����5Ұ��������&d����T����
���[.4Z�S��Gyl�,��e���%E��я�W�*PEԮ`���r��'aϱ�3��
���Ȋ~�	V$8��l��T7�n���^˱Fޙ��\�S+X���B4��)�wH���Μ
���n��\�4>M��6��7�C��Nf8��$g~�2{.k�APĴ��P���^��E1.u��hfĔǲ1N����X{'s�&�8�E���hݤ�w��&��F�ǹ[���,*h�؂=�[L6@PN�[2M��QK�v�
���2u�8L���Q���³H��`�\�o{yb�5 ֎��-��]��I�K"1�WnG�Ze���˔v(y�W	j�3�R׬ ER�`��@{`N<�e��b&G)y��؅�>�z����!���e��9���6CP֛#R1�_��2�䂰����UZ�`C�a��p�YL�}�,�բL{\��l�0aa�L��Xw����K/�������_���07�%��ASĜ�)*S�v?�4�6=�.(����-��[]�)}Uh�U�|9��@�r�܅QV������Ak���:.��̴�~s#����
��BF��/�U/�?朦/ �y0�W�h\�V�� Db�;L�!����r#"w8���;�63�B����C�J]��Ҽ������m��ȍ�:��<��� �2��*��e��<ۄh���Ď���H4����AB_�S�ˑ���8��#?>���`X���XO�҉�"����z�!��^�W�+s�d:�sq�@���M+]���Q�?��!=��H��F��ޗ^8�z�u��30�T�dL*��p���܈�T��#���ȗ����)/�u%ܷ�$��U���e����<�0��we�^�(�v�co�J�	��o0`=�tz�)e,: ��>}3��LV�2*1|-2����ќT{�a��a�����>�[Q	���l	j2~�!d���TN?�[�]��Р��MDSwTI��L�DZ����.,ӍX�����1�Z�m7�2cӏ�R�j���;>��>�0c��,�d�(�珞L��!؝4��e��������N0fK��ъ�8k㡿��u(OB��M��I
��8��ck#�~�5U#�
���>��!y���G�u����|"�����v��)<6����G��]-���)\���̕�d��E�1���Iw�YS�W
ޟ�=�sg�z��@h�Z���i��t)G�hg�nL���E$� �i��z��Z�d��]N�J##4}a^EDa���E����3v�$>E��{����cj������S|Z��˴F�|/�/�b�Vú��0Y��Qe���a%Y�o�֣��N��������&:4Ko�8hd �����k|��'��]�S,��ŭ���dK�����7+;����e�t)8�ˆ��62��G�*�Va�>�aH��w [�㹪�@R_��z����!�����}wU�<1�1wk(,��&;>�P$����0*�g�P}J�����P�����k3/ĹjBs�wMm�Q��{yힶ����U�$��[����V���Y���'��4�T������q�v U�l�Z}N�b�1 v�5�^��͇0��%q��y��%b�k����14��ƨ�j5+�������]y��EWn�!�.F��|(Jb��
��d¨�M~U�2*�ǁ�B�]�{�8�Z�SL�y����+:S����gp b;`p%$���F2p}_��u�TI��ĸ�����y��S;���t{��U6�Q�Ҝk��-(*�1fC���6?���%�:h�%FS�"N���u�-���:�.����);P.�����{�3�q����͘Ǝ������m�x��Į�_iOQ���8y��;6	h�/=�RMh�~=��I�f�.'�*��H/����ޏp{ �,��e��
�}����èip�$�x���=Hk[��Oc�꒜�l���`q���o���(x�VEܖ�a�y��#���#��R=~Be)P�%gyz� *M�s;+�/.�
���NFHkٸB�"B�J�Iǲ��mi��JJS|K��2��בM%�a���m�]���G���^��{�j���:C>s���#y��%���'�6³����rN�Z�R~<N`�)�	c!)���Ί�,���7�D��O��ʄ�ע���2�:�@3�j-qRE�P����'}�6k]��{9!�y�E�&^��7n L{	;2��	��4GW���E�8S2�Z��=>���V�}_|k(��gI}	W�XZ�}��+g����UT|D(�=⭋1��8�M���=���%5��i?��}q��Ipr�����f�BR��?���O@$y���Z"�A�=��,4�� �O~OcXH1Y�!�X������+�Mdis/�g��N;��� }`4�2����
���W���?&��~�7�0�A����i���IS�bC����ߥ;�X����#B�y���vZO1�أ�ۍM�Om��7v�uM��	�6�������g�e��D�(0��C�F��ۮ8�؊q�j����:��0����e�y~��_L' �)Y�+��?"�hbV��eP՜�c�^
��	K`_�E|�|T�7�>C�q�� 1Qh/m[N����&��2��8%!�,(����^1&9�8 �Z�/���!]i�,����r���s8�6�����'>�]&cL1��^�01��1�
\OKR�l��W-+@��+���d�ǋh{+/m<�e�"���Z�H���Ã��YYcwz�4�v�<�|�Ԉ�$��U�!�ʹ����j��"Q
���C�kӓ����3Ah�$��<��;��/���=/�a}�ߌD)�y�~�o�:�^���nr��q�_��1/�"~��!����.� ��Iz������Q��rU�!ɼ�+|亩���iɕ`ue|ES��O��a���:��8����x}�:j��'D��B)��� D�C��xߍ&vc�:A���d��@�1�S�O[a�"�E/G\��R���@�`U�b��<s:/�g����p�Xc>�^tS��'}� WA��mx���\����C�O�'�z v�0Y��#>��P ���*��3���!�8xlW��b�D���7̨�E�$�J�@o��]�sF�f�"��c��Oy5h� ��-,Ez�-�#���Wo�қY2�h�J�^��Ð�b~�Zg���hh�ս I��������,�#�'�o��a4O��j�Rt�U�]vq�1&��:���ݵ��}��x]��L6J�Z�B��4�( ���ѭg��b�&�����/���4���4Bsٞ+6��2����P*vq���nL��1�ɲ[�r�5Vv'��#��+�u�C����J!G�{�Z�Ą����3)�t&+b�s]��h�'�Hq��z
~���T�[z� �VPm�+B��Cw4]��@N�A�G;qe���#{�s���I_��y#���������@4�j���L���Vł}K/ŵ�,AM�C����Zq�9�8��T@�0�����ۜJJ�M$��e��w����
:W�G]����=?���(앒n�h�ĥ2�M��{�^��l/UM���� �ܒ�_蠟�*�ԏ[jTh��)���:���uMsiIg#�h�v���,%hU1c����f�<�Y��A���U�W,=�����Ԟx��yt��Xy������ђ�	�r�b��� ���[�Q��	�FNgր"P �������멱״�A�/N��O��d�e�=K�m���)j��T�RU����6����i(��=82���,�$ln�bx�
��*�#�'�wo�l|O�H�,��������-�X0oۉA0ělY,�9��uT��ǽʭ���0N"�g8��&<��4u����ϼ�@��O{�C
�蓒�\������K�;��C^���+��y����������jZ��?�E���%=Pra�0w���L��L�seke����C[���<���KcL�]�,��B)Fm�5M�	 fX�fh#17JNL��o�5^Ds����7��~�4.���Y�mnN?
P6�D-O��a ž�@�~���>V_�n[�2����J�H�S0�=���t�
M�
�]�@E�ߦ��alߊ��Mȹ��~2�)��n������# ˱��$:�u��7H6Y	�1}:�s��
�o�1����֯EӉL�`oY�b�PkD�/@���/G;V#j^��t�e�L�����<���`��2s�@��Ȅ祴�5�i���r�)���:���5?|\�kb�vl���auA^S�i��`.��d��#�-��_'h��2�l����NI14Pp2�l'�~]V���33���M���I���+$&���m(#����\�wS� j��F�(���s^�V;.��5�I^��&��m�=`;kB%d��2�bI[!�ƕ�'q�N��U���Tw��A� $��և
g7� �,�
����A��M�k݄�����;��eރ�=�!�����n����k��WA��c~ �g��?j�8��$���	��X~�� E�=J-"���Kd�/�� �ǵ������y�ku����?��^�W�W��,!V������<s��J�љ�Ħ*�52���)A���-���I�r�]����N)K�U�"r�3�:(����<�ѐ�SV���C)5���}���5~�N:Ȑ�֫��+c��D�3X�s�FCn�^�m xYpNj]0���Ij��0��GQ��
՗��tM�����Ai�U�����MQO�1$:1^\.~�N]��2���3��6Z���.��-�v��c�h#;w-�l+'Dy�p�/ԥ��n�hi�~u�͘�5� ��2��c���ez���i=�hL��3���:�X��b{�?;,�l2}}'ND�XG%�1���?�<7͈��Op!��V�k_w����p4���j9�a����R�S5zi�=:�7���#���|��	4bB�Ԟ�v�L��ú����d�����u���''aĶ���^���P<n�f�<�./F�o$=e��g|�k� g��(�ݕ�15���-����w_��qZ�3J����l�W��V�C3��>:${����MbȾ�0;{���M�v@�di���hI0�Ỹ��q�J4�c��#��O[u�<Ui� @�]�{&Z=hQ.�$)�o�u=�!-�!�8��\jvT�+��=�ï��(�5�Y䷼��s���f'|\�Z�UbI�X��
Y!�'���z��ף��`�k���9o�%{����_�22�@L��!(c��@w?��k1xX���=ߠh?B�4� �g�K���e�������册�m�Q5�d��Ḵ���.�.��wd>F��$�_���*>�E�����$ar��۾�$MV+M*�|eS��o��y�
GSD�ׅk�c��S�$�9ܱV�SOri�kb���u��1Iww��Hǲ�C�z`�a�m?��F�Hr�r��W�'��r�(W$�-��p-�!��gbCv�
�[/眑��4',��D̷��p~�d���1�-
�p ʅ�D�r��!�s���S���3�:F�NoQ���Q���ʮ��%2^�O��!��}�0��kA�I��)%�AA����Dk��㍀a���*ub��cA-ڟ^t��Tg�k=6��א�R��Ӣ/:Z���nz����W&��	<��_���~	��X��7XmI�����Ŕx�>�h�O�L�Aҳ�vv��	*�N3�톶3��.#�'�/�MPZZw.��e1�.|*\���w�Km<Be���t�q�0 ���+DQQ�����؋CMl�e��F��3�V�эJ�	�]}*�clIxj��d��}d�;�)E�f��@q����X5n"�����&ç��UT�x���+ބ�/�LT�bw|iKU��{��o�;��[�TRn�5د7��/�����~at���?C��%�WV C�V��B?�)���$��H+�P�z�t�0�4�R}NJ|����2�r�iy�q��$ȉD�9Ʉ3"T>4f�	�x02�V�8�2t���z�����a�������5�S��R�_y����6���4��*ȼ��6qH�0E?�92˕�fm���8]���Q����'j+���A?>^{42CP{�*x�'��^z�"�q��w��Zł��'o~J�2��QR�P,�������#�FY~zn�{X�yb�䙳8<��T@V'վʭA����#RC���5�
6���)ϴ�H��j�
�ʚ'���,cK%�=�O���Lu���Z�$XE�v�(͠�V�2���"�rVa���&\h����|�s�ꓪ� ���K�Z�[Sk�D�"W-̌Ē-�Ҏ�j~�T����Ʊ�E�o�1�;6��	�e��qa�w�)WZ���U�v�4^�y`>0j^.�M�80�����f�Ah:�eT���m��f믧��7#���u�/�*��B<cI���C���`$cVv�c=��k�*��%	_�̖W�&�ʀ��oͮ�)r�� b�}���f�g���j�M�C%���ױӄ��z�Ρ�%nV�{A�.��1��Ahs�Ԕ �y�RPT���w�_�${i�J�p�Ԣ��QB]9��3�
Y���K���QL���(����6�C� ���Z���L7�.ֵ3T���D4-�m�d���S�=������]��j7�2�˻\tN?��1,|���C�ί-:$6�"|�eTo���'�|��.��W.�FЯ%hϐJ<��f�"��{8"&�r}�[r�	u���,y�U�Ձ[���Eq�?�h��U��>�� �!/L3J�H��A�~��S��U���.9
	� ����å� �>�xy���x.�2S:�- [xtbP�6��}0���x
l5�ّ�RQ��k�@;���hV�w����%��H���|�,Y�9j,Քh�P��ж�JП�ۍOp5�Yy��uf�^�.4ȏk
��b]�i���D�I�^��ݾ3��\u������^'��Z��	�@�T�-#n+ח��3d�=i5���	S"�[��&��>\n&Ex�B��`��"ѯL��!�y#��L�8ۡ�QA>��f�tj�c�̔�p-m�_/��!�� ��Ж�d�Cx�>ȯԲ�Gze+p�J���YJ�j���Rz��N�@�|{��yhkN�	�.W�U���,L��HjDͥ�"'h���L�ᦿ)�-1d�sk,B�e���K<����^�4 ��]���b(�/��GH�XA�V��ht�����t�]����M��(�����@�sO�T(�0�1������u��%���?vBY-_j�\�cH�mc_�_�Vi�>��W���,9�40���s��<���&kc3@�c�S�/�eB-��e�V�����s��;��l��������1�_�9fhU8T��z�ݶ�՝�V�-�[V|�B.%i�(,L��)�½r���zB+bB�kmV�Fv �RniS�>��B&oW���@Ɲ�����J!g��^RZ��V8��m]��C�T?P���wU]{�_����\���Dgn�鈍�d�{�/�<Ju�mɵ�l�-�b(h]9!2����;|VXR]&׊r�z��U�r�}j�s��c��w�ԥ)��t����Yv�\����I-[:W��{����HG�1����u��R]��S��N��`kA����� HQ|;oG�X�v�@�<�$��!�w�q0���يv��}�u�Ff�����8��YL�~�h_<E��Ћ9~�W\��5{�!�V��!���P�6-��"����/�e���J��<1g��m�{���ˁ�;Cސ����e�����V��������j)������B�;�X���|{",eXMQ�^�7���G��ݺ���1��u$���g��B
��gZ�R
fYy�b�k��|���p��f�/#��W��N��U`N�f�J�����^g��4cf��*�>��S7p姯'�_�������1��W�;��<��̨qeV�K�c	맫0xw��ǈ/5�%�<�����l0|d✗uW��3��J��V��%�)g�]]����3�oR�$q�Kd�tȗ1Ԗei=N^��0WT�5��=���&�J���Qۭ���À�)����y[j�nrq����v���Z`R��>��`L�v�	���M��Ga
3nA����Y�OZ;���pI�<B���=�E�>2o���բ��2�l��'����U�R9čH�;Q��N��� F3���v.��V������M����v�I��
+#I�x��q��$��ܦ������D׈���g�On�[���"�k��C�E�_�N=M�����7&qRt�e(+����sps[3��2�^'8�$cy]�]U���}6�7��7�6Is�[�q��L�8�yq�aN"e�a��'<�M5o��D`�
c���DѪl+% 5�����%d�9mOn���a
H�_t�3s�k0;���1hD�H�@AA�r�75�|�*�|�r�qW�J<�a� >� &)���4sl�stmnS���E��
���Yquǩ�?�< �b���m/�=_�T�e��Bd�Ei~����ߘ�-{7EH������>��p�L>�z���ސ���2��F���A��}I 0��������Yai�]��iεLB�u��ΕA"��3��^'�I�S�}:˖�+�1r�J�6`���@���iLe)�3��o"&]bI�9�c�|o�Dˑ,���&-T�-^)��.!��;W�&��a�sZl��Lr���Q[����m敄㴛 v�-UI�����3�!��N敏�u�$DH�B�Ü���U>�~ϗ"�W��[m���zO<���o�5x�im(��:��Ր�	3���ڷl��MFv<�����,@S i�N����m�w�rt��5�w�m���"���A�q)���w�!����r,Ff��P����Yg=1��k4E�i�r<��8ugc���W����8D_�<!K8{�u���̀����Հ�t9����4=���E��?��t,;�s�%���}�A������4}�&�� I���[�-���K�~�}�$�z'��ȧ�+uM;o�:�@hQ���f�b�� 2eYGBiu`G��:)�[#� ������=�/q�μq����w �e,�y�]�P��v�]7eA-��X�uË���%��m��lN���@M��Q���D򨩐4/W�2 ƞ��D �%���hx�Ƨ�2��i��w95E��&�7�v������a�w�	�� �)��Ku[_��Z6��C���J״������F��I�����.[8�8+�D����,E]!w/Ͷ��d㘳�I��=�q�S�ZU�Gm�5�b��y�oZl��!x��I-�V�3��9ݸlؙ��D:��"��H�'uX�<�� 4����=����_�u�3���-�U[����'㧴L�OV����7��������b휙�+�Q���p &�7��7L��Z*�S\Fp��ֳD׍z�3�Q��C"N6�˜w̠�b�_wSqd	�N��:�P�?���~�)�y+�r%�!�dރ �#��>Z���9�����
��B��sMAq�Z2_�X4D�@_�&�7�D�d�|]G�B�+���E���q�����m8��ůÎv <��MG���(}�u~�n��d�&[�.�FSTM8 ���:�,.�'12����ʺ���Ff��`��CYg�`���{��	�<�M�i%ڌ�Z���G��c�MB,:�|�Q'N�x3z�ݵ�,���鷮�}#2�vJj��-�>�o[CO��4���Q���p����$^ﳣ���}S�n�0_�r��LD�BIY.��"�Ե@]fZ\+���V��rxN6 �\�u�K2O<�4p�}��(������e%n�3rL�u��.Rv3���S����Ҝ�~�1�/�����C�vRϡ:}��XB� ^B�(����"cl����J�vo�_�	��z��s	��+fnMYDsuW�k+@ze�3�`L%?u�.�x���:(��������YGϿ�$������� Q�
�f���<gHF�a&fS��$J�W��N�2��r��I`�Q҃�}�ZƬv#^8��o�á�Ӫ]C�d�uI��iAC��m�ՒO��`�|W巶�ɹB��9e�P%�ld����u{��r|Y=��ֵZ{�m�~�Cͷ��}P&�R���n�P�I��.]w3�@�LF�܎�Ѧ��f$gx�ɿP��%�lg}��7	5�i$눒��~x�G8��Ꙁ��x��q���OF{K�)5����]���+�
� y�P|߮oL��o��X2����ry('t��Gt:��'���cm�Ssݦ��5e�V���d�+ᑐ`Ɔ�W0K�B`>�3�8����64�Z��D܊��Di��#��i��\��m�4{ >[U�����@4����<�m�݂]eD��#{3�~�E'�>��}���Lb���쬔R�3�(������e�����DyF�Kq��W��iZ��T br���]�j���]�I���8�{�$~S%����!��|h�p�6cz!>_܏���4����ߖ�����Gi���\j�­�47+��MT�wpz�۶�2�I)��O�e�<���Z';�0����i��q(����XLw
�Jx�hd�I��w	�MY�MTdm>�3���A=H���hP���4�/0�7�a�xJ�i(�!�s7=~pC�^��&l�o6�� {G�V�[5���ڳl�M�T6���m܉#���^3`��M܁�l`C�i��\.�y�?��0�ˢ�Cߋb�� �8���=_��y��m��E;�M	�<�F�u-�56A�d<������?=��ect�u^� �S�����<3�� Ÿdߜ���,##����[`�'35-��G�bA��f�
Ĝ��Í�kh�Yѱ����O =K�G�b!���!`�FM'ŋ���j�3�j�;�0�"�\13I@K�_��+�^���W����$qԒQ}��m��Һ��L�cF�E�\,t���%F �P��w"w���N�	ܷ�u����4a�躀T�(����d�.��?�/�4\w��1�� zPL����Ӕy�h�'l|(+��.^̡2�u"�͟�����+i}`�nѦ��-��9~DD�^��/!��BKd�^�U[j�o�2�P�K<U0��n��MxD;���//�J��lL{�6��	1���h��@�2�S𐱲Z_e_$:�?��<z�e\;J��0-
mK�B�~g���k�hs�����%���؃S�8�u0�F����(���=ތ����Z�V�7�<��Nu|���i2D�1g�8��g�܋g�.(��/:۾� �)^�W���%hx`{����wZ�(��%8��6PDfRӍtg�m�vzvFy�G��f�O�����bg�U�F�﯑x�	�@�^i��<��i��<�.E
1O�CH?[Lɉ��cI٠�3ЊXXC��FiE#\L�U��U�;h��/�3�Cf��nl
h�b������%׎p7CR���]�E�蔫��n�(*����|1���!4�qʶ��v�<�w@A��\䘰�d*�"/d�O�e��c�*�m��*A�^f��&�~e'N��q�_J/J��+М@k>KAc����,�H���$���l�=��)o��v�N��F�A`��/4y���c��J�H�e*��Q�OD�ه6�f�x��V�o���2,�U�5Z�C�<��-�a�yP!3�]�����f>{Ɉ��=�4H�Dc���	�p����Y�6R�佧��{�h�I�6R�pS��-p�kG����-�Z�>܀ZB�.QWN�d=܂�8��^b��g��P s����KE�[�]/�O/��ݬ4F�"����=�^}��˛c����N����6y]�$#��	ӪA���W�u��"���ie?�1TWm�@E��m�r���4�<���dc�����A�w�5�W8OE��cY�|�
�%���^+��,G�������H���<x��KX�aƓ��w��,h2�㇕>�;�o?-1�zo^�-yꥱ�U��tW���Q~ q��<S�O�Ot�F6e��/a�Ux�q�&�<�ק�P�@/#-kh�l��@���*+���r����ÂN���9�j���%����s��������H�2�a���%]��_���!�R.Ø�=F�Ee0v� �C�TBeV�3	���2��z�kB�����.چ�* �����n�ATo�_P�J����r.@J�[��c^?���4 }���f6� �_6�NQ�P���Y�V�#�!�nT�����!�Y���!��d}��V��Zrl�X1����@��yB� 2Wq�)2Bul���8��K[�UP �a#�������&�*�ȿ�I���V���m�YB�:��v޿.qJ=Ղ�[�B�}��։��E�4��BK��q��O$T��}?����N
�'���ޓ�S(�\��Eq�]lA��m�O�f�g���E�P�Ņ�D�DE�8�L��d��9�Tt�p�D��&6K�x�JR�Pb2�;����$�Fe�g�]@�ͻ%u�å���]���]-��|w�Ču��T��@Śf�AY � ������з����T͌Qy��'j�2ᾛ�%9)�E#��>�ga��ħO$nق��ǘ9y�d&�Eq���
U��v̖���"�p  ��$3s�3��FgL6������Sa�3N㢾����M��AP"��όexCNp�e�u_������nDK+���f�W1����/ΗzYhg���?35�أ���Hd�K�g�F�_�G�0�_�5��-�G �5�|!an��i֜��V��@k�o������ 2j6�V��Pm�� �L?��DY`�zmpus�d�{��s�	Z��l�(Ę�6��Z�PW�.��MP��b��=����7�g5�	���u�\[�WD,I�&���/=���i�<�i�/�[�8�G�P��.N	20þ��<�\��4��&<.燯!λ����H�cٱ��lh��p!T�>�뻍E�<�:_Nl����ě;�V��jM�O�ջ_���7�x��X�̐��R��I*�K��(�Z���g��z��_��]�͚�Q���x+�%��:a$�x���qŸ�}�/]�Y� ��}$ z�(�iĠ��C3Ih�r��Q�J��#�p��-�1E��X�!��#<	�����>�)��ͫ��I�r�W��hJy�H��*���fw�ƚϓJy����O���pSX��Bw�t��(af�VH^p��|tZ�Ņ���s�'���t`��h$�;='[�<6�^!�WS����LYL��c�I��.)^�z`+�}W�kV�0I������6���`�#uu�;��:U��k�#��i�$!�H�cF3�K����J*NVlӍ2p8�Ռ�3���T9 O;j�D]�Y|i&�'?bw��E!5@���
L�^8")����<�C�ڃL�[;Q^B���Y��_w�.Ũ%�j�f,-�z؆4����&�
Is^
�]�가�I�~���0Z�g�f���%��yE
�mT[����i��A5�ٛmBdu��R�f�����R�?��?i�Yr�:H���4��c��!�V3��Ϻ��������M��E����&`V���nSֵ|����|��Cl��w��-� agR�EO+��k��w�ɤ��
��e�n�{���c�g;'��S��98l A�$3f�`�����x�lKА�Q�D&9�d1^p����*���~��4����>�j���v�b���D*�F�TX[��D��K8��Q
����Z���'�C�(*/�(XO�����H�ݣ*�`��y�
�[/s"��"�r��X�s=8���@�-^a_"c���Fڪ`Bo]��:���2�L@��;�D��!E�<4�DuV�r4�^��<# E���/�R����͸@gLMZ�z��-Gt����q3���
�%����T� &#Ð��W������a��rl�L��ѼeǙ�Z\��&|��@�r���A�tRO��I Ip.�ϲ�͡)�:�  L�'L�'P�b�����DF�h�N��z��~��$� ����N�.�\/&�K��ϗ�[e��#��&	Fr&d �D�c.'�)xd)siHLg�+����Q��E�3^�Vs,��+��IUD����b4*kO����X��^��~p�?��J_��w �gH�Fl����K��=�j����84%�z�(��)�ź��4���ﾺ�8��A.�j�='�p
$[�u%����J�����kޥ��Dm��S�U���DyM�{���,�S��2�g�D�	Ċ�۽��1{�!�"��s�gU��]W�hG��VrDr�)�S/}��Νx���V��\��j�dA�����%��bƶ-Fe��x����GμH���G�XE�<����'n;��d������L��W��|�<k:���&�	�]tܯ&�T�NKJ�8t��(�>�����Z��[��n2>^� ��{U�0���_�Զ�&�8�N�!���`�}r,���t$�V�
��բ���e�`����k���0W�uO쪻8�i��u���<��s�wUq�Xaϕ}eX!���òԜ�����L�q7������>���>1��	�_)5�SgWI_=U[��C�4v]��%7�AQ�`BC��h��� 9����o������9�dE����Ç(+�¥@{�n�ɉ�H�cu��+T��vt_TPk�r�]�G��:k����ͺs�ӴC+�X��%��U���Cn����3�H������)�[ł�-]��mO��!*MDVh.W���тNG>�"G�T��A��Ur��L7_���[]����/������2ΚL퓴����?l�_�0W��X�N��~x,�C��j���	K�� q��ٳ�����ML�q?6�j��,�� ��]��C���(-X��L�l�_إ ��Z��%"@��L_��"1}�@|�jonǢ�i��Z@7&_�6�i��	PJt@.�.� �I��w�1Hڄ��8�S��8@�ce��*�ڿ-�(ƹ�:�쭐2_,9I����D� ��k�����e.͏�ȵ�F��vʂ�c���d�! ��FG>ĝe[~q{���y/�X�:�|�YEw�=��lI���
k/X�%���_)��c��T�0깶�9Ĥf�`Z]�9�&���#��lLI�m��9�����@���`k�@h,�:�]�N�T�Uu]Y��Q�.H��l�At� N��ݞ�!�����%��j���0�־֞3r�-i����nc#�\�Q?��'���eL�m�$ ���A_��`׿\\�8��ޢ��Y�����2k��;�eż�H&�޺�^.��(@d`K�v(>/cB����*i�@3�.j'D��N=���������s{�.Y%w�v��X����s���}�q{$�{>��`�E�J��嘄֑��I��Ipb~�Yc�Ч����!$���7}�ہ��S�����e���raJvɶƕ�����q!}H�AK�F�B���=yE�1�^;̭����k\R{dD�����z�:*����/a:r���!t��/-414h���]4��f�cP~�kᵃX��o��aq��7	��W^��z�,����]?)c)��2���`��)��4��.�ͱ��� �$s�a=�����f]���� �@��
'Ԋ��	�邷��(�I5�-,���R�kR�ˀ!�YQۋtP��z�_���J��Uǹ��p
��n���v�~�YZ���xcY#\�Z��Z�yyo{;Ƅ�e)�|bW.�3���$b4C�x���9�0嶸Z�H����猽���)b��"pGGA��Ч�U��j�>�����2�86�TPUs%����� 8�����f��;�&�r�+/�KZ��u
^s�کz+;���\�6��J�i��Z\�;�v}��J)1Iʼ�g\üzc"�e޾�G 5WH"�K%Џ��}F��[�p�ٲ��_U�?����1���׆b嫞J�U����"�� 9�h�{��'�/(:Ђ�GTЪU7͠P�@@c��>��Y*�$޸mg��B��[.�1���(�Q$����wT
���g���0��??U����24P[� �/!�� �'s���Gc������~o��'��cr�� y�?��]a�<mV�AV��K�U���.��a9�yjـ
��V����C�+��\��&�}��k*o�.*wx�������������KpL��t�8��v�D�E�))�8uPn� }�oF�! ]p=<��u��h�T\��u��K�YzOō�~�$:�2��VjoVdڸD���w
�teU8�q�J�i8�Z{���'�yt�b�_�e[S�R]���ϰCx�Xtn�@�	~�'xl�i�C�Y���"O}oK*.�9(Y�8Q��!��"�XP�s�_z��ct�x҈�QO�p��G��'v�3�By����â�o���-�b'�0�a^Xh�Do`g��}~ 	�Y�d�5$��r��г'�c�K*���1����Nb���
��$.���7��*@�A_9�E�6���ć�;A���N��V0ʹ���>��u��C��̜�l�M�@�jt�Ɖ�=�죔=�?0���z�+vi�h����U<|�/þ�c�Io�窯��9sۿ}�39,~��
���W��@$X���`Eg����v�$=r�α�u���@���؈�D����w���ݨ�}�Ńs>���`�c{�P�<O��pX� ��܅|"u�g����h #͑�Ύ7�_��!N�� �q�p�0�<f�G�������e3SA5%N#KA��/U*}�s�3բ�rF�A�"������gᗪ����I7���Ř��s�V���뷖�����_Q-�fd�L.���]�����7r����~�V��������D��?&mz�/I��a���3�b~īc	U��<ѭv�'B;�I��N[r<�z�TS���v<5v�#�Hd�@Ό���_e�@I��N,|jBr�{�<
��0��J���:�m͹ ���k�h��e�Sc2�H�ax�����g�Hۖ�hG&�� �A��:��={��9A4r=�w�Z���b��Ͷ���-n���ש/�jIb��~0����_.X���:Ӛ߾@�{���"���$/cFu�i/���+��M���v[�rR�7�c�tkMZ��&��3&:m�Ϯ�>�(�K+��O��/��*,�P+��;r���^��0g�.o��\��G��#�&�,91���A�H)o���Sm�Q뒿.^�b�Ze?�8V`%�ҭM�n@��GP����rza���jbg�U��2��2_V�� ��Gi�~�7B9�*e1 ge�;�?��Q��yd=���O*&88�#�N��i���D��&ӫ\/���B"%hm�#AI Q�\R�9ejrh��ߑ��B0-�,�n8L����(�)vמ�3GL�Į�wP����x��!e��}O,�7��/��JQX�MQ��8��)�苟�V��a�S��j:�~�8��Ե�W���<��v����R�����1܂���9�C�>�����E�FF=��$�����^�%2��-=!{�fLb�B���"���5�P�7��)��͈C���,+�PF=���S�Y���'(��h6��;VsL+�Rw}�pP�q��g�Yf{/�N�jT֓�&JN9��S�5[�B�Ѡ��Q��.P�cu�u�(�x�D�Õ�����{{#'ܶ@CfU$@�K�8t�M�D���zʻ���^e�����X�u�l�W� 6����8d�����ö>	]Q���%�H^��hes��[�vЌ#b
�3�\�k��$�6¹��Ty���^CM�Ŗ*s��^%ә��|9�����%5o�H�&.�}��2f��M���15p�E��ȴ��<b/���%���z�A��51�����9	���2M��kqN��V���3}i�hs-�Ą���u��eϞ���,��Bu��yO8ģ�H�>l٪��)�@�� <�e^�eR ZC���f��7��E
�b���mL�l�GZ��4��4���m���-�!3�s�n�Cⷒ�I�=�s���?
"��}�o�������ȩ�46�g�TY�0��et��!1�=Ά��z����Z,:��XA�'���(H���]������P]�d�0���5N�!OC�M��;�1uJ�����vc;�5�����n�TT8_7F����I	*ў!�����ܨ0�3����s���:����vH�	*��7�����̽��37Fv�U�u���d�E��
�s@E�c<[K[��<�Ǟ.� �?�t' Y�^��3�%��h�\�?��R[S.�m�P^7O�6��y��/L�ߠٯ�ٍi���F3�F���S)k��#��M�$�C�~f�qO�������&�A��MT���������1=�)��I����gg<5S�՜�9\5l$�����|��l�rq�h�X����?f�J~� h�JQ�X)��=��.QNG=Ff�yH4�7No3��)Q���j����&{PBD)�?�J܇M,H�*v����>�A�{���g�*��P�Bq��Ұn�OY�M��K�Q?�j�~�����2����X��QӋ"\:�v����hz�1uPO뻎t����D�i���#7��*h��@u���C������3S�q̊@Ɩxק�#kBri8�v�N��}!^-����	���-��\�ؔ%����?ҕ�_+�Th�I������X
l�cp&h��>�p��/���S�vp})덺�L 9'd@d��Bn��>YF!:����U���g�Fi��2�v�w�9 fu�n��#{�L,�P�c������	�7	�jP�6j|��&{]��(�و}C{�>�T�t1���%֍G��g6K���#rY�#���ӎ��q�t��Ѐ���lR�sp��*���<9��O��ҧ)�������^�A�sDѦqs0��6����n
D���,eQ��2�q�N[���H	���ʚ$����F�|�d����E����1����R5�Dن�=hAF�f�6[dd�]g
v��<�;[@Q$������(�����]Z0⥪��d�1n;F����-?��a�h5}�Q�n�������ʟP����=B6xJ����= �Rѯ���$Mwi�l�^�{��b��-u�"�kGuC}��'����������o{~P�����:8fi�0�M�[@@�h��+w�z�7`(0ږ���f}w9.�����:X��w��sR�4�����
�m-jM~�yϢ��Ǌ�� -�:��IIO�Lx��U���@������27��w^��g��$�xoi �I*����%����n\�e�>6��;:���,�DǴxBl7^�gs��z�&5�%�87WC9����Y܈/�j�z+u��?�`Ci��&q0��ܯ����2٩�u�s2����T��9���No�?���Q��w�˛7���0*���T��t��W"}��4��r��?��� ͑ԉU�gV_��lIIe��|Df�D��7#{���?�D�
W8��4[M2��.-׿�0Uo#V��O"��=e 'r�7�]�A�13H0Z�sH�H�s��*X�j`	�^�Y�� �x��7'^�1ɺjAP��hӄ��G!��I8u��g��\��% 1.�_���ua1�����D	�<�L+mݠy!·%D(� ��Ԝ���3?��3$�<>�0��;~ur���<��\>��c��9	"�ݷ~��z���!<R��J�]�E����}ޯЧ��H���H����e� ��w���P�i��̜h݋�NBFm� �ed <Z�����EmB}�0֍��D{*�pг���K���1��i�*Szc&Pr���D_��[��Ow�v��X>���p��eꆋٚ�	1f�(		����r�A�<R��ca�)�ͅ��t+��^�6X��b�5iԂ����-I�����<���B�]�f�ܷ�\^��"��m�����n��"�32gh(Ћ�n-2�4��l�	��C�pEs�׬�ᔂ�Ï1��cV���f�v�MKG�G7f=���p��C�~�=���Ku.�~B�;���iY�Ie|�U���O�]^�i����U��Y�]<��Vi�9���dW����(9}��Dr:|�No=����BD~�5#��ݱ���-��z����J��0�zŉr�fY�����ķ<�O�67�l���\�x�gP��䠽���M��Q��JQ���hc����5Z��mw��S��f��V�"T����f�7/�	;<����P�L�mSPya#�U�@d�҃a٘˒-�,C8�w���+��F����[������$h)�4ko�#��i���w�����ҏ`,���j��K		F�m�]?�=�g�'��OΆ�M�L�{�ޓ@������
��"��h��P��W�����bd��?��J�I�<�uSCN�>�漰q�Ϥw�����8d��/T���u,�rhnLq_58�+�J��aRʛ9���==���UZ���H��#3��N�P�Q���Qx�t�/�^���^Dx�E²V�P6a���c��iz�r}��s0�N
al�"٘jk̺_rp���GmMז��qjZ��*�� 4�k�|�z��$䈏���$)�o7�T3���Di����(���W����)�F��ѭ1�
�E���4��g܅��[k�9�
x*]���.�m���1��N�gԍt^���k�mH�nו�VI�	7���y�V
��Z�jM�r��)�.�(nc��S��3O�-�9N�܊T�|��F��Vy��}��0�C\��։��� J��]p�\�W������=yO0�*��s՚�.�9���,�Z����0�����C�aq�ɨsiD�����E�y$ԂzF��7a���@� P�|VJo�&�$���[t���=��*��>ܸ��� {��9�W3M�I{Y$�6�6k³��3��Ȳ�Oi����f��`0�C4��р��Gm)j�j��o Q�Qi_Oh�+g.��P�ǟ�0Mm'����K�|1�������lá2�b'1 �C���7X��&���:ǆٴ:��>-�6`Yk�-ې��m@d>7����!֬[1?N=Y26�%g�cu���"��d4�PQX5��H }@�[t��A���`������Ưɳk,Q�����^���1bT�꠰cҩ�lUf�όJg�۬-'M�E:2��շ�_^ڪ�!�"DN�r3��E�(���sܝ������{Oձ�6͗D�~ɿ]~2	�M�1"��~1�6�g����h\`��m�p�FO��ׁ¶�p��ֱ���x[�Oyz���@Ӵq�JN��o,-��愎�'�W��{����k$	�)�ͳ�嗩��fBnX��A�y�m��������b; �\3�!ƨF�bU *et�g�� 8V��x�Ad�=�Ց��IHnY}�Z�
ٍ�'#�L6��!��B.)#��!�m�C�8n��/��(?��� �ɒJ�*�ߙ�0Fp[����� ;,㭸�rb�+���b��g�n�-���Ґ�@�[�{��P�}�&� veWɽ��1�9X������l
�x�>�l6��l��r�����*���Qa�����bf8�{J_�cK��:;��O��~TX<�'�]ߣ���.��� �oML��.H���V��3D8"d؞ϯޝ�xl�*���2�P�h��+�װX\ژ{r�2zO.!�F��(���Y^*]UQ	y��ؙ f�����j���f��m��bc�ׅC���j=��e�����)h�5����ƸФm���i6���,��Q��?������[��Q 
�h1"�(��5Eq�PX�%y��XR~���	��N���J��b�5�DKI�3\� $JZ��Ȼ�?����ܻdt���C����.tϷC��L�}O��NC��bߟ��٪~��N�R5i��f�}󿴗�)C�>���U(�o�8Ŭ�h�¥��ȍr�N�ų���(��d�[���K�è�\^�'Q��\Eɼ�A��ɐ����d<�(#{$�5&>�N��tq�/�V��d��_3
(��P��an8bu���5�)۝c��6P	8�^�e��[��E˿H�g����L��Ҩ{>|�Tj�h!_W���|�4�h�u�����V�/�˟w�κ��h����Ţ ��	];�d5�	��	�2i�s.5R��b#���:�Ph��WL���@�唆�"РV�:�D;�V<���G)?�w@�h�[s�.��=M͸�S-��TN��H�{�`bL�M$Ko�i'<*YY<��M����)>��	�uDH�����)Tq��#��
I�BZ�,u�P8pEQo�#P���)$DBFm��$��Ch8��~o g8�}��f�&��z��rR�;1';��y\G�xC��1�]���0)���Bԏ���	ii�)�h&�\�X�f������I`V9F���y+�����$똂�'2��7� ��6���*x�`�5�������M�pL�.�E���F\��8#
K��A_W�0	��D�
+��o$�ߴBLƧ=7��>�2���tb�<��"ſ7˕�C��驵)� �-��W\��z�O�R��g���6��I`�=ِ@7D���bq�Fg��$�0.�v�(?����}�e����L5��q���o���+�RX����*[S}�3��z�����~K�c?����oqY�L=�}>�����s�8Q�~��@\D
$c����5|�w�gj¬a�y�P�w�e�T�M�=b�z���[ ��M�0�v�uږ��?�B�:��;u� G��̤2�$k{�6����q��`�����:����K����f�~L���CH)�����E�5��eL�v�E�E	ɮ(��8G�=��t��+	|֝L��ݙ�}4=+��Ȁ�G��g���#�'�U��
� �h��7�� �	�,0���y�/�χ�)6z���z��	�UD��r@��R@�q�@s\a�B�������G%.
���xf �w>�暔''� Nv�KӘ��'8b��4e��+�I�mȢJ[R�T&ZӘ����u��6�S��'���' s�"�v�ȅ����HQK� ��v<">wo9:����E)%0����[[ID��T#�~��t�:��7/��R[�	�-92��{���{XL��$M[M`<#���޺���pr9��#u�qᗛ��\v���q�8䭠�m� �#i��C�g9�ͤ���!ُ]*QZZ�b�H�Ҫ���q"�W�vϣn���W|}�Cň�|A&=?��|h���ײR���E�����ȕY�}�����r%_�dLU+�7>�A94��9Y/6A�#��-NE�����ޏ8�cr�p� YkШ�˂���ĉ2׷)�����y��6�\��UA�r9���c�����yR���u�S Shp�9����'87n��y����z���������uM��w����ͯ&���C��N'�#]�-��:J^86&���@)͡Cn�Y\���<�����gҼ��EO���D�҆:N�g�S:��VЊ~o��`dY.�N3�8{BS�� ������^Ĥ�x�Ub��A����p����ƃ���Ȅk�Z�1/�]F��uл���ۉ��K3��7!�w�I؞*{ݴ�	ۮ��-q��%�@K��l6��NJ�_F:��[F�}�L>D��}K8SL#�`��+�d"�Y��Р�)r�&RkHf�=�}>���o���Խ��ٰ�-������6�v�c9��K+�oB�M�������O�II�4Ƶ!dN���lqp7��e����,��1��[@O�z3�ږ�U�j�9�m���t&�)Ūo�K�t��P�R�N��z�pٞ�{7e�4��Vmk�T+涔���I�&��8� I�������6`��d�Ʀۑ��ck�����Fmݸ�Au���q��=ך�u���}Ce{?����M�|�L�(U���H��z�G
b��G�[������Ӝ9W���d&�Ia�.-��&&�Z�m���B�%�zY�:R
fm�.�N^�����I)u��h��`Ą���P����֕��VhF�����vh���y��)�����A�33�� 0Z�a���UBCN�e�kۦf��'iXr���0�N��5A�+S��y��~���W�x����� �+�m��
Z���UWË�ur �1H.�����6DH�%��V���GiF�� �՛�Bh�(d�`S�:5��v��^�.9>����;ųF�#F-x�$�}ǖS ��0S��F�޵�-g���k�*��#�%0�=�~ʉUrY�2������y#����Q���;�t�ѽ�H��>��#V��#�� e/�v3��>��%6�3戈�7��[����k;!(�{���9���Ġ~�Y���v/;�"�e��s�����@��1���vg�����E{=��+1�jQ<
�΢��W�]:5Հ���1�2����m���gͥ3�vq��J���)���4DK��t�5�c�2�	,oŀ�eW���T1�,=@��fK����!,8c�:�W�I ���Z�7�׿T�my&��G}�Σ�'l�#k��8�s�Jb��[��0�'���د�Q���3�z���t�����~�3��y��I9���ᩯ���ޢ�c�"��P�;��H�a��2:�'FG�OKV����c��U���M<�3��fȚ�({_�F���M,=Tہ?1�=���9�ض`�ȟnpa,4�y������I�P��T��ܙA;ex/=EI5o	"JA�:<�)eZƻ"SFQv��)��6�膶?��׮�<&A��)p��X0X���'x���~��j�j�>v�ܗ����Ȣ��>�c��ٛK�۽��\0�/EɓT��P�je��3�C������~��O�/>���ް!�S55�7�^e�w?p�aKv<QV{���G�B+�����C��U�Z�y�]�ڇ��;��54lE���&a^�J��(��'����o����V���D���,N���D��D\r�1uIN�v4������3浫���m.l��C�:��S�|4W�I�CY����^�����!���[/>�Yet��g%��2��g3V>�L�$c�L���6�"^����e
�/������XDR>�!Y'o��C�F���0ـ�ȓ�ظ��<���=X��*	�������*,��+l�~O�!+w�E"Ŝ��5<�a�k�zY�&�N�@�ݥ�\�&K[13�5�,��y��8? h�1Z�����T�{������ 
6AC������
�-9��F]}�.����C
7�269a���K_Q�Ћ� �Fλ�)/�&ǳ�xzZq�7��e� �$��,	At��]n����<ĺ>�d�C{�-}p~�PϼpխIl������}w	U[}=D�{�5��B0}a}::v�V{\V!�q��	�C�À7^�찠�b/�� v���Sz������+τ�|�r7e�&��f���׌�z�X�N �~�AOKS��
'����Łj��8hڱw�,�WTj�1��R�h��X遱�Wnxz'+��-AXvq�{�� A8�[ՠ�Y��$SfU���v���	(i[ y	��ܙri-��s��|8����A-���G�r���2��f OII8߭@Ћ�І�����s2S�6Q����a�7S��vȔ�"���ў4�yQq���+~P)f��JKg�=�;��۠������,Fy�[ӹ�$*��q}�/#���.XWc�����[CJ�D��̓�2�s�S�;r,�9�l�Q'����F�k�e��|ȥ��r|֢�ߚ���P��P�~1��S�=���m(q�3�� \4�\o*Q�����-���^�e�p�����ȕ��1F/��F��k1C>˧P��e8�F���!���OS�����>�4dz�E�j�P�w��Y�2���f��A��	!ɶy7B"5�+c��Ĵ�\�%�ˣ	�s&��{����8�i���	�%�ϓJ����UG���Z�����J,��#O�w> ��QF(&��s�˫��Q����� �&�a�3η`��=#8]�~�89�\+nΧ��x�&��M,������@�A\X���*����{�o�/�e��K��WMS�	�@iI����$�V���M��ȓWOW��t$U�����y�G�Q��}�^8�ec�M9� �G:ܝa��b��B{�"W���3T�/v�v�%���w�[�cE?F�=��})2��)��3co�����%���J�S�/ơr��9���K�R����"�~g�Ξ�l<����a=�R`��N-�3	?�AN"S���pF�,s�s�{�}M7�%����?=����<м�4���P8n'��mD�8���K/8�Ç-�OT@Eg�~�G{<C+�u�%�[�q1��n�x9����b�/ �X�d<��."��y�yf7ZK�	�1���ԋP�����ߣ�pF�G	�葡��_��[�	Dv�ߡ�3�L�XV'��xY�VW��$����U��ά��ƾ��eM
����ߵ�;��ڢ��b�M;��&�1�427|��Ue�1�-�D�����S��L<[�\�}[lDW_0m���^�}"yq��
Gݸ�i[�?���O7�� \%E�?bYO�
�$���i�; �$0X��P{�E&� ���˕��`�ٛb��RO��)����S���(扦5�L"�Jt�pL�&�w���U#Z+�\� �f�^��T{AZ}g��~T�C��E��8J	9_ k�p����jg	H_���4mJ�M³I��I]�8s�(�zZt1W�'2b�U�Un��A�;hz�CO��RXtXjIz���:��7�q�[��9����V`E>z#�����k�C[R.Z�7h<�����q��M�{��EEFt�@���;�?�|<�y8�쟕X�Wl��(4s�\��:�.Bh�o��Q�c�"�+F |N��ْ O$��k�G�28��b�֠0{�DpT���g���O��좦���8IH �@zɊ-�G
�:���o��"�|<�������eD"�p������� .����˂^H�~7'���7�0]����d�8+�6���l�׽DI�� B=��|DQlA70kA��b��F���T�"O\�'�+ͅ��s{ V���߰��';ɹ��r��X�ؘL����7�N$"ڎ�b�ځy�݄`��Ē�͡#��GQ"�z�7�O ��؇=[���$��2"e����]��r�ɏ�w]�&�B�	�R��Ǚ�jӠ�������ó�}��C�
�����!�n�)�7�g�wjZ����< zhhb/�V2�1�7^�\y�ɠ> o(k`,zՌ���2�A)P��;�1�������_o���ՇY4g�	������ʚKβDK�4R�,�qŐ.���^�
u����5<_t�˿�~��;0����f�%c�UZ�!4���^���ϫG/A]B�劶[F�`���_چ���&Zw�s�N���f&�5�#f���G+�ה����j��9�^�Vl|=:�&&�)o>�u�˹�P��5������!ЂIW���K���U�7}�J]-e��/`Q
L{ n�k��.�������桗��e����NB�-k��P��W�������M�+��f5t���K���O{(�w�ǎ���58�n��{-�NL_Q�g��ݨ���ؿU��y�l�;�.v��!���՟i�b�� kx���L�J�c��m�Y{��������,�e����&������*�I�L�k�]&\Wb$ �T�����j��&HG2#`�J:U�����!܌.�}�D�ʄn���;�E�r苫unجT������]ȣ�ƣ$_Yl�7YH��.�C��Y���L0{�������xv�������� ^�J�8w%�De�V` ����Z�N���Bt�����)�E&���k?���:[�ހ5 �6�~�"���ĀA&�uB��{�m�!K/Wa!�O1�y�X��Y���5 ��Q#��sz.m�oPSe��4�<M?��6i2$<���h��5�����B�����w!�[y(��ԉ�A��%�6��I�9r�ӳ݌K��ڡc�U�:^pi?8&��P9�~Af��9{Z:�vڰ���z=���!h���*�d�_b�,�/A6��8�TE��h6}�yO�ED B2_�sS��;
͈Ք%?��^jj�p'��5jt��U�n��,�vn�3����j��tν���E�)�y��p;ϖ{�^�2�B��D���'����� �w���f�bu�+M3-�n]����Rԍ����`�̰6p9{ؔ&�WiN\(II"З�A�a L����x��}<7WW��a�}����۸z���s&��@t��gDy_ςŢ:��ٹ����a�2%q�ҷ-�×���X3Y$Hɀ����w��F*@q:�l�G�-!-(�*�g�^
*�K�#�,,�,^� ��aF>N8y>���Tm9ΔB�E��uE<G"�w�T��p��UM���#~�u�mm� �݂���SY���y���A���0�:�YO�c=����M���q5����)hb�N��1�]�CiL��F*�y*�����^2doDcn,xC�-5�t�G�ð[t�udE<�&�K���4��6-sȞ����|��5�NA�`��3<��1wp�O�;����2.�Ġ�`��< w��t�;�j�+Է��A�QV�ݾ]4n&�8���9��l|ĳs��Y�Q�l�l�}0�Q��|B5��x�1'7�c���[�A�	#��]N�����gA�1�{���1�\14DU52�?���22$��C_dX�����-�_�#D���W��qV�����z;%�[��kLS������Q��������,Q��.�	sf��s�i@aڅ�止��j�(N��=�ڪ!�7"�oF�!�[�ɯ\$����NkVc��._����__ ��]��K�i��������䘩%�w>M ^����V�!�f]m����&�Z�3a�J��F��}ɠ�� ��2����?uUK�������A8\/���8.�hI�3�cYv�v�6X�n5���̊@�/���i܍ϞtN��|n;�����x�z��'��\�L���R�;~��fC�����'Ar�����o����I�K�2(�Zs6��6��W�K��{�]3��4���O�9�e�&��FS#��A��bl�T3�Q�t���J�ޝ����Ų6d\�s�"%k��ñ�����Y�gWF=���@�����rJI	#�s|�4��v���'Ό�N� �	��� A�P#y�+	/�����^�!r����r>Rj9�@&a��6E�؝Q����&N^U����B:M]��&hb������ѿN��i�+�z�����yEI{�05<�&7�94{�<f#C���˄�$�ö��g{z�� ̐�e\��"Sru�c�ruQD��.~PRs ۥ8Oav�ǔ9�.�"����b#:Xy j�s�a���*׌u��_��ܨ��~��xU]�=�KYv����d?��ȭ�Z׹�^�v�}P<�i
�(0_v��5�'�汘�����ʧ -z�O��M "�Z8�6�:T�� ��rD[A,tG��
�j��"����l���y9��s&�?���Iܨ�0�ɣH
��`�k�,-���n�uL�ٛ������U/�FZ���c��lT�4�hA���~mpLKغ"Ġ��e�3���=�~��!hE�i]� �����78F�I�"��ll�EgDs	��&ф{���K��N�e��?�Jy����qDR ��ě)�3�E�5�瑚}V�����R�m�
��
��l��*�D'1�p�R�Ķ��M�S0�^CVч�=�S�,�(��jsE	�V�;�D�TA�@�{�ۄ󶅰��F���0UOt�L���lѪI9;��=��1�iv�L�C���TLص�It;&�S�M���4:]}��:����@*�gP��F���c���߮�����M&�#Nb�29�L�~�c<�v��hi��kY�D?�GF��P�uL�J8��Oi���T�mWY�]kCS�ͺ�݌�=�3�{��`)���y(	���^��G_G�y_�4V��D".���7F�qb�[�8�o��pl�Z�)(u�P5��l�¥m~�Ӿ����b������hʪ}g��(
����ٱ�@�б�e��Dx|ӷ������P'�4�i��}�v=(����ۈK��ӫ�_��`���G�v%s;`T栄'd�AW';.�x��It���S�H�˸�{����eϧڲ�Ө��h JS�'�p���/l�ΙV[*�=Y�J�
ڰ �	�پ%$n01�����}�`6���`*��i�+Y�`��"ə�2����j���n���"Y+�|�Q�T-ý�������=��m�E�XY:i25PҖS?-`��MQC௖
���f�|~u�o:���a_�rhaEZ�pK�L��ȼz�t)Bq������wR�
~�� �F����,Eӆ�oMo�:�����T ���щ���C�<���%�?���U�zӱ�_����ڮV��9�t�s_��bm,�ɖ��iq��WA,�<����rl/�!e�<t���~�)t��]~��������t�OǱ���Խ�
�(���>��(�/�3�ު���������>�͇'?<Z_��hԏ�������8T����DA�˟"u�s$�q׳=����AZ�L� ��тzysEQk�<��L���& !���E)?�<g*b����C�_#�4|e������ [���2�ύ,̭�>o]���c�;+W�J�ʂ b�*�����E��g��Ų��4mo�Nsm X����Te�7<�ϴ�0��\J,��Ǘ�gŵ�ӵWz�Tdx��|��;
���g�e69�[�ȫ*�Q�Jٔ�8@�n��it�.^e�GU@�w"ذG �������gu���X� ������mEŖ�.�P���0���f��~-��4N$��_`���.�F�P�ao���oy�R��"�z�o��Ȯ;
��=�z�Q=M}a�Ox����D�9�:�2���=�`���'<@�@B�a��@Q�!�#�G�|�Y��Ņ%�d/�xj%#�7�eT�፤��UM�IRSI��aCk�c�
���y�ɚ2���F<W{Ɔ���T����<R��r�N6nk5��[�|]�0�,e��?\���B�I};�ܼ
A�m���Qw۾f/�U�G*��-h)QB�oV	���m�.�~�N���ϻ� ��<�D�S��Cp�P�@���D�|%f,�z��A��4�t�C�ſtX���[�Qo�7�������.��ڹ �((���}\:�\jf�1��R�!��'�'	�w ��L�kt��Y��l�rn�{�,o�@�U_g�%�����w��:�s��V��xN�_�Gߥz�Xy�۰8�#W`��}���ʛ6D���Ή�S��ZgY�.��8WMMk�T��KC�9�K�QI1�;��_���>3�G@������"�}�Y\�ǜ�������5��/�l�O���u��6'T{Ӑ����o��+~�ډ�e��� P�
1[3�����  �U�����Wj��t�L���x̾��/@���_
�)ˀ�>B
�X�~G��^��z�G�R?��jG�ݤZ��4(�u1~Ϻ7����y��nĠ��S/��I�V%����U�H�{Z/%Ώ���]��N��C�tS��R*��MH�A+gK�X�@Σ���v��3���	���� �Z#��ts����X��߮=�n�n�e������v��&�Hs3�-~����U% ���5�z��m�]��ԲzD/So� �nWpD�{��E۵�-g�����A�E+�ek�̥2�]�̇��� �X���)�b{�C����2Wߒ����


� o	潂]�t�����	�.�Mz��Ь�cЪ�+�a��?��0���z]����c�Q���$ވL��q	N3)S��>E�#<�&P�z���6�."�Q�ߟM�i�
��ܫ��SYw��&F�x���g��K�t���$_e�I@���k �*5y����S[dE툁��<�p�������S���X}sf?Sm2|�D����\a\��r����;BB���㽄��TV ���E������*z��>��,2�[Ode޿�"��|����Y䱫�'����Z�]��1$Ϯ��9l���9�_䜆_��$p:A0�e�&�R��X'R9��X0�"���l7�M��. 		��������U�y�:��|�?i��G��¸�l\z�f��o)$��P�q�}��jw>���ϸd����>���&	zτ�cp��� �g����=U��	�1���~]�Ă|L �#7�D�ݫ4������:��Y����:AcU;b8�ze��%
	