��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX� ��V��P���[Z��W��.^,���mfŃ������s�T4��Q�����\�X�	oWݤ
Y.�zS]0M���0��>�-�Eͣ��16�e�>��>�@�o��(��t��xJ`0�)���%t�*�%7�!7�H��zY�@�c�~�`��3pW�����m��'���ʼ�
;=D��;��p�#Gp��(�����/'���"0����8�fYt#��?����{�⇱{'I"Qˬ|0-h�E��f�q����4O���;b�$�q3~�o;�#:P���N���w��7��́�Db������u��ށ��*�ڌ%m��R���\�.*����[���[��:��
~�]�rPF�2��F���v[l�{��[b>�%��c�9i�ڟ�؏�+ʰ]�89,C�-����q$T���U�� �KA��X4���r Q�_����R6�.��e��ܺ7˽�X�ۧ5nW�Օ�����+�*XJ�Ag�_�1u����m�>�Y��Ry�����U)�M���p����fH��M�J-
d� ����\�S=�N9Dx�`�3�zu��7ݞ��|�gk�/5,��Z�+֚�����>�k�;�t�:�]�3P��8ɿ��/q)�T ��V���V���}���2�Z%h�5gQ�-�L���~�A��`=2F�6'=����&����g61�V&��T�̭1� ����},{�%�� ��=:�D���z�pD��E,D�4�6T��*!�N�yve�����K���%G&%�L9L	���x��*�`L�ۼ'���Ix�D�9�3�m��+�b�Mr\6�:��n�kELLV~����Yos�ê�7tJTڷ)��e���f(
�r�ķ$�b�S�,(�7C�/��r�7�|ݝG�܉�P������d
&XEn6�*�&F�W�Р@S+2�^u�9M�Y��I�}e��8����
G!�9.��Ş��g,��r�_�� ��o����e�ܿ']�����(mj��(P|]���v�L5�IϨ��.2MP�q>��lNb�S���'�7R����3J��f�l���Q+��p��h��	P�#�O(87n��'�K�JqȴfĖ�p�����[-��i=�R��������l�]��<�8L/yՈ ony���L�V_w�2�֘�����]ϖ �m'Θ����iK�i�%0h�c�<��&ec��[WU��?[��F_�-�&�Uf���'���5��[}L��U��o%Ƌ�W�ސ���1�����j��!�a)St'1~J�� ܱy
g�����(I0�U�(��=���$�̶�oG�\�P��mݒmT 7�U|Yl��o��3��L��s<u21Qa IV�P	�lL�Ř���� j�t�\��SŢ�:l�����h�����/����9���d-�P�Gv�o�> �,��ZκƵnRp�k���'��t�f!��&��hxz^G��-��ո��FG�2Fuo2��\��y[�>���^�KLs�?� �@����cJ�����~xq�:7�[�|�3��DA�J��Ӊ�s�ԏnx�n�r�Ȍ6��[Nչ|�-S��0Q(��7�̫� �c�JR	�ix")\4׫�4��kP���k��c�.��54zl��G,��4P���sfx�Y�S<�ӄ3B.�~�mǗOG�,��D�=I)�)!yxKG����w�*�߫�e�w��M[D�H���T`f��x��;4�7@���kJ�b��t̹c��r5�ԋ^�O]q����^��Je���#1;�Z*֤x6@/}d�XS)h/'	�r�R���<��G�~#�Ȏ�:_v���8�J�U>�1N�b�^��n`�E+.�bCjCC������5�/<�>���ۀ�j��W���,�� Ε=k*��4�y:�����!	I���V���F|X�;���R����W8HR�Q5~��Ȓ���.��w��h�lx���>f��?GNc���wҨ��*�������~���$�(���U4I7WT��V{�7bl��0��Nm��K�]��3��A|�b\��{J���N)J3��*s	7v�t���Q_ܗ�+�*�?z�L���79�y;�k˴�����`qb��E[[���@��׆�3���Oh	��K�,����FV>�j_����VgI�y�e&���_F�kx#����%�p�)j���y�4+f��;����0�N����j���H����:ՏB�����i,�K��r���Y��yi]��B�eM'�����)��/���N�>��7�5�����ń��cTu����s��t�8 �%<�ۏ �,�n���`�[��H%����j;9qs��` �j���kL�نA�ɻr;D7�ƴ
nM��$@g�9��Gx��;�[��?���_���O�cY]h���s�X�!T����2Gk^\��.?<t/���ϧT�ԛفf�m':1��N�*B;(]}G�h�?�]&����"����L�mS����I��f��=���Zfp:�`�����������q��HB��&YLR�sg�����J�V[��QY#a����r�<�+��W��:���[\Sð���u�|r�4�����S�sL}y�N��+� N���$���=5'{�3�[}��1�޲��Q=�C��A� =�G����\���q�����1�{�T�h|�v�)���B����8n��Q���P�'i����!��Q4��1��(�Q� D�T}M���L�-~���q�gi��)��q�]�Z�İyՖ����KI �Α���󴜶��i��a��<�������U�9�fNb�Aj�A7�e�?n��N<���G��IN�/�x�8~#YI�.�e�>ِ�Ꙁmz�<W��1A��[P��oOr����.iYkh�����{�*N�KL��6e���,���.	(m��g}�(�B ���DK��Sv�R��%0�^ɢ��͆�B��)�xNRr��]�>��,��%ޘ�-��*��n>�"�ڙ1�4��pyz�_�$-hWycN��FB�Y=�х�L3�>K��Ybqhq�`?�ev�Q7n�5�����B��h����0�{_L�'�g我��ҹ:�ڱ\�\�R��~�f�Y'�FV<8z���sp&]Y�=�[�y�qXi�Ǔ;�S���=[�]@�_Yhҿ��E���������_k����u"���zދ��nQ�W�p�Gt��X �R��rܹ��y�r�4��>M����ЋS�gX��:2c&ѳ�ҋo�?Y�AS�2Ô��f:�m�����x�(�C>�ϛ9Mz��6��N�X�,��[�_�`�l�/z�[�X�0��,o���\SxlQ�[Θt5�Y2��h��1d'"���R�ʢ��%KD�t"�3+u�6��d���NE�G	V�.x���n�.�
�h7�>��)<�\7*���~���+������1��@s����	���j���p��s/5�S Xp�|�R�hJ�/N�`B�������'Yày�|����������vQ�+tif�.� ��c{�(�0D!�����79�%��ES��J���bZ��pW��]y��/�������.���6Ex����)Sz�����'���㱖�Е��hd��2���m��o˓`�Xg	Q��&�������ZG�O[�|�3�����/���+rBs����8����A&�lr���3<k>���X��VBS��m�3�eK_Hސh�M�i�B�-[kj r��Y�]�
����	�a:������D����F�!x�N�ڿ�tT��[Fa��B{��Z����(���2s倧�6g�CK��$�7o�i��ʎ���:~s͞���m��<g��S��y���ʨ*���%-D�S���A���V��J�Е ��,����+��`tL6z����, d�t �󧴹�gZ2T1���KYR"Sc�lC%���M�Ѿ-�bŵ}���i��P���z�����`��~#�N�����4B���{8���j*љI*�{��omyY<�Zd�\"hS枷�:}�ȁs��l)z���C�m[�ig`ں&�|�LT�����H+Mz`Y
O�����=4��d��U[@��W`!?v���� �"��=A�ʄ���'d:�ea��������[���d�C���x0�x^��]����exbl93�a�f(Iم2[���wNHDC;�EU��*>f�3J�L|5�jY�9���kf�z~BG���jC�]���ў�wr�#��O��)��F�������t�d8ˆ����G3Pft0�� y�1��X���;dt:�"m�R)oΪ��~�^�4�l �+�9���벦>�j�.��};�¦#��40H���^��,��K˟�����î^�i~wv0V\��I�ș��x�8�_�~-����h�}�:Ez���Y�����!���DĴ��8��K
y����۷��u��gPL� Ҍ���/`˅	%6g�"ΗҚ�N���i\�+��;B@)�i��{���I�io�棤��Ľ�r1U�����x��$��~���wh�9�a�%��D
k�Ӛ3�w��T�:1Ϲ�W8���}�h̓���U���V��M�=�Ra�|AG�S\s� �֤� �����<�D6nF�R0�8"������� j��~1�`Ӌ���!鄊�A�yz�q�<�A-�8��)�����&i�,P�2Jv�eP/��ӗ�=u4�?*5:k���d��wp;'g��7���V���{�D�N	��X�<���d��՝H͖i�^̙Dq�p�]�� C'x �g,��T�6��ZO�5d*�O�r�vz��	���x&��D�X����t�X��9R�}��b
�ҽ� �ӧՁܹ�o4oޕى''�Oy�����cH���?ֱ�$#�/�y1E�rw'z9�6$�Pe�����zU~�S��l����܃��H{��#ӻ7�
kYP䍸��O���l�������J���<�cVT�!gu��xa�e��tL���x�0_q�G�J�vN@ &�����ԝ� 5X�G��%Vţ��[ �C*G���z���U��C,O���O�L��P�pl����@��|�,���174������]�:�
_T_&�v :��♊��}��,K�{4G�;RjϹ���;.՞�/����/;r�����v!�cI�Y�'g�1&�<!�W�n K牗�w���i왡��]���_�\�MZ��7��z�Pq�F]�B3�V
9K�C�相�.��]�;$-lX��g� ��̳]�p�Y��b�U<}��à��Qr�G��;�G�h�&Ҋ��3�*������0o-�Y�\"15=0��
P���9���Y�'��VTr���;� VS�w�fnZ/'��p�,}1�P������M,��W��ݫA,$G��d���M8=�Ә��I�7�ZZ���My��WƆf��E[�=���p=��9I�z�&�L-��u$i��qZ��f�OD�w\3�_��<L�l��C ,K٪����%+�������gP���A%A�#����!Dp&uq|��/�ű����{�|Ĝ�J_A��)��P�6S_��Dd>1�>�g�f�ڰB @��cy;d�a�`����ҕl$�	ޗ�ßʝ��f��i�΂U��;�8�O6}\�Xl��|Mi��fg�э��-�i3��h���0�Ǔ6h��%��b������'�beN��+-�t���`~��~�a1�t��Et��$�4��s&˷uk4�ҍ�3O�vm���I�[�)6��D/�:ϐ�Z���Z����5S�T�2b�ݛ������M�N:�q�)���BX:N���O��	Ǵ�g(��ռ��	���J�"{�7���5aI�G!�ó" *��-)C�����1j�b���p�	���)���K�0�H�����X�[
���rPQߙ�)����sLѼ��w��r��t��'��c>��w5��d~�,5!T�?s�N�OX�6���0�`&�cT��1�����.L�x�^�hH��}N�C��R�)�&w3~|sI�����|��F�S5�+�A����&5�m;X��c˥ �"`ѹʲ0ZC�w�>�2����o�Ր3���[_��C�d[B�XȜV����%��E����@�7�H��6���0�W����ߥU5�����?��6�P��������:���y�b!f����=�f���VZ�o嶥�7C��\��_�fdYA�Âh�GeȬ��ԏ��g�p�2-3�h���9��BK&49�%pmq�9 D����걗��݊@sQE$!	�.�ů��m��	]fe��4"V#˼�|y�h�	��r�*��ŃA�� ܷV�Bw�G�ʝ�h+D��E.�z:Mj��H��M�h�iH{�UL��_������m@d�Θ�j{Xk��r����݋��-W����'��x��S
�iKo���G�W˗���c�����Q=�t��Ո-ב�qb^�+�t(a-4el�k�F!�O�䗰t�,I�9��6����X��P]q�g�s���#�6=	�S��G��m��2B��dO�g#VVr��,�Н٭Z$��%�1���L���� U<��u��ۀ��E�"���а~IGoΨ� 	F���j��]�e�߾��:�g7L�#Va�2�+������&Z�����ڬ�q�i	�eS�_��|�V� hͰ �>h��I�E�sͭ^��ܙ�aF�G����g:�JCk	��u%WI�I�졗��Q���� q���~��m�uL�@��ǒ�@d���B�d��a�TR��x�j<���?N9�k&ԭsRu�E����j�c�!�Z�Sm��	cm��~a-���A9��|���j��	�lm��/�h�H]�:'J�'�cOk�D*Ni1�Y����n'�FI��d?$����Ay��\m��ƴ�pv�`���5�av]�Ǐt�h��Us�Z(���H�=����m;�Nv_C)ф��7����(�����	ƫ@k�a���UΜ��������@�J��Dd�i��J�/�uR�V l�XS�7{A�����2e/W�QX��n%"�-�������Ӓ�/\��+f|��?�SgBX�ɍg{��v/��&����<��Q�G��^�����J]�m��X��"W�|ڪ��%/�g��y��fO�ʰ� I�C����g=�sTpaY%�����:yj�G�u�W��=����ޚ׆��y��8�y���yj�ڕ_�a�t�v���j�ؒ�7�,�2��DΙ�5q�Ź�&� A�*��*�fθ���<-0�Xx��٧���i���F������pHR</���K�!Q�M�b~_f�qrď�+�R�ri��7�<�W^rS���|u����hJ��:Y`�j��r�e6��u3jT`�Xk�=�w(4��ִ��:'t]-"޾�\�0j�}b��S8�W��=mr�S�E!����@|�=ۈݧ�<�~Yw֐~PH>u|���c���W���ݤ�ׯ������HU�t��ҞH����[�3����.���u�$_��C � '�~�m��N��h(���As��ǡh{�*5��Yx��0�_v�`/�h��DNi��AGk� ���'�T�qL��gL�2�[/_��4j�����SS��ͬ.��J�q�u��׾��pb�iek&*�L��r�F�ky���N���x�\Kh7��y������x���[����Y>�N	0h7YO#�JI_r����Z�u��۟��
[��`�7l!�"d�rg�m�i���������^����\�N{rj?s;:�>�@=�����>���k�.���)W�x��q�3>����$%�:�w[0�41~�j>91��(�5�����)?���ς�����5�A�eEC�Ǯs���*}�|���4�Y��>�G&� r�fs�N8#{T�5U��~1�l��D�z|���B�ҜR"�����n^W+|�6��W5+f�7�+���ej:�m�:q#>��%�U���8�`��O~�R����[��q�֡�0,�mz�-�R�g>O���W8��J�hD�H?h062e��:����&M�VT����z8F�SH�E�S�s;�h�� ��^�3�a���}[�j�0E�+x��2~כ8Uߙ�M<��<h�jg��Z`��(�����7>7̶Բ=�Q3Ē0Q<�pz�]/�g� 
Ȳ��ߔ�����)�`��� �_��uH6r�W}3�겵���a�GX�)r�[f��и�� z�b�(�[[�{�w���r�����W�Y�e8����+\�g�c
�~�s�R6D���kV ȵ�D0!�	B�k�����L�J	n΢�c�}�Mt-���>�	�K���&�ӦX^��=ͮ ;�ҭ���F'Jݸ��3������c�\�bS�2��U03'�'����5!�J5*?��
-}�����ѹw8��Z�Ե\�?��'b�?>�J3jc�Q/�y���f')u� BVu�//yæ,�v�9���J���k K6lZ5�����`YC0�X@ĤfO����%������f2��U"1ֺ"_�nΎrm��W�� ���(�:o���ٞ�Bc�k&{
	"���9�����;����ƪ���N7��b�`���)*:m�8���W�%�ᅬQ����tv�D�8���0�U���T�mOL��J�nP���`T��4�hqϽU���t=�Om#�J�.��f+jC7@�8�+�m�w>S���NF��n�p�������m�s��5ض>ʯuВ��l"�9nNb����A����_f�`|:�M�1M�xe��a12�S|1��{�L\��M��
kz���()���@X�!F�x�䨫:2O�W�=ӞAq�g����fY2����^W��d�-yz�LˠJ"֐a"���-3�΁���*�g���bŵ<6�^ڪ_ͱ ��n�JIٜTw�k�a��M�
��5pw�Vح���b��U�瓒,l���ʹ��9;I�8V �"i)p6;OK��ץ��P(���P�(s�C�!�����u�����>ȥ����k��%P�G�S�KK��P��*O���+��[40p�?�����*��ut60�ǟ������7������96���>�Os���'��h_R��h��u��@���d����Լ)�����/ɂ�ZϥŤf�n���x�#mF{p�`���kx�I��BH�
����w�x���l-t��˿��E�?�����(j���j�W��S��xtDP��}'t��Y]��3y�,4��e��!�P�+L�N����]F>�4�M2���B+-Pg2���8+X���L}�*'���h���+Ce��ȆrNDp˫����b�I���{׃�+��n+aN�We7��;�'д�_���^����6k	L3�|K嫱����ĵ1jxm"�{S�����Y/T8�gu.;&�&(�NHɴq�:C�!h�n�Ra�bdL�k�&k�4��7��LH�3I��
Gɋ�!���mxs0�9��P�A�m�MX:i=`pd�����q�?�~,9BJn��TپmTJS�᱑L��0���O�BW�6�B��:��ݬ�c5f����p�y��n�,�i-:�-)�{M�'oM�8>��J�I�f��O�A��aL��J�N����0u�킬%��g҉�u��k,�v��+ڵ�M��"����Т"$�˛�[I����jm�UD�f8ź~��V�A{��;��ng��M�&��!LjR�۾y8����$kt{
���DFªn�d���S�����$���+��ī6�P��V���?�C�Q�iPk����h�󜒚�uş2����kȤlU:�v]P���x���̈́f6������m6��m���u�v�m�X�j����E�4��V��a.P�^���=d�������O�l��{;0�"��^M��$xZgJ��|�SU�r�o��e��i�Tk�c$��Y��0��D%���%+�[飳�H��1�Ȅ��nD4�bQ�cL�6��`۰���61�_��0���92�φ<�uR%l�;)�13�����K�C���%�9E�-'�	�߼%
�,�S����<�N��v��*E�Z��F3q����2���mG-�k����25=nK��w�e<A��}�UֻH���6��,��\�ڔ��.e[M�"���5���BMK��J���4�:
��������z��|�JW�ќ�Sg	�,�g����+��:�q0ҥ��_%v�^��k���M�g� M��ѵ�:��r��+���؁����06+�����BZk��P�%��UǍ0q0���xy�=ό�=m�@~
�tUy+]���k(��L�/��8F��m؉�����J~�*O���
{|>^��=�&��?*g_];jO�W�č�$�,�Z���{��oe�T�[�����4̘6�ā?��@u�/	2Tܬ�w6]q�=OݝO"c���$u�Y�	�������#Ϋ��f��EL�I�'��k�r]�K$QCM[gֈ��3�����x�ƽ_�M��I�ǫI9�預�5��m�|l��%80'�Ω���q�)Q��/!�uNtK�&���N��{>�Gk��b7�> ��K�}��p�Iٕ;ga4x�x��p�I�[�>��6�y�_[��[��F�=L=�i�<d-+�.��燪!nj_�h/�Y}�{D�kו�H���7I��o�� �Gk$��6x�N�a)���y>ѡ�4F���:I�Ia<y�\;�R��8-*�]s;�7f@,Y��`;*
�6�pV�PQ�a��|�$}N-)0b��
�^3�	Ǉ�4��؋�ڶ��T�)��ʷ�E����_�8@����~N$8�'/����UwceU����c�|�.L[����!C��D��i�:��S��%������K���	s#}
��T�f��-j\����R7����QQ����#"�>{�g��K�Z,���)&=!����a"wִe�_"�Ls���ye����Q�nr ��t5$^��^��Yi�����6�,�!w f���u�sev�d: >�R����㴀��r��N2���A��Lh�Z���;QZ���[l��m T[���F�f�v�z��b�$�O6�>�ގb�1D>��`�G,@���r��J���]-?�|���ش�r֣Y��	�����$�z�_���`���4�0����s<+=��>
�}c?��	k�Eh�������Ed\UG�|�0ďK��7Z"9U錘l��F��F��TcL��]X��mB���쀼c2�p]�@�Z�h�<Ĭ��Af���9�B:�k���`��E��-�*+����=��2�K������)d����ꂮ�*� _'����|,��JE�P9�K��Q#�c���t3Ge�v�o^ �#�2͵��ƣ���"�$�P��K>��������[%1�{�' ]�_9����$��元/�8�b�|
�����7�.�ġ�a�~ӭg΁�]#�N�Q9'D�L;���AXהAfda�A��B�$��U��d�ӄ���+b�Q�,�>�]{��]�4o�="���Nz 2G׍���@C?����l��Zo�?UK5Q�/�WaLz���L�g��+C"?�r��?����k�Zm�,�b8C��[#�\�/j���Dk�����:l��oA�M$N,6ף���r�4_-9r�JQ�.h��B���r�Ls"��!T���{q7�����^-b4��Õ�_�xK����Q�ΆE�jV��2⮦%�D�	6�6Z*���tR��i�S�'������ �,Q�n�B�2��V��<Jpfe;y���Z�۩|OPSU�G�FXB����WhV��+�`��e�j�:Z*8��O�DJ{F�Y3ߕ�z׵s	{�h�>��6M��}�ٴ)fy��s��l�����Cw6R��gM&��;gej6��րhY5�#����}�W@>!Z[<cd��%���M�?t�S�L!�B]�&U�zT��:������C���#�q�HG�m}L�� ۑy,n��ʑn�lr��^�@�����Qm�ŉ�m���Yو�`A�����1��t �0:�T��Q�z㚐�&H#w?h��(y+��{�_�ss��i��&gJ<�#d���{(EX����	����oS+�&I���|A��k�%sSh��Q%��� ���ܝ36$��%�}|��� q�;Ā�;Y�iY���U�����P���{��ꥏ��s�H��<RNpr����cNHS���J�ׇ9�.����0�a��4!����'�I�<�F�+`-P]cc�V�sh�����R�is�y$��u��t���ñwF&i�l����v�.�9���+H�<3����uũ����3�F�b�n"�;����Q��0ud/���I=���H|s�l�*U����e���
�X��eZ
۰s���Mʿ��'?G����C�5H����<�o���fxV���Ɉ�u��x¢w���sY����R���ڤ���wR��pq�u�����@�Im�2��{���5�#P�_(���^}I�R%���F�	H>��Q���gnO���@0��m9��ݨ�����
3���B��W}p�A��Af���|��	�-�3WfE�1Q�+5[���`��h�<��dս��ZEq��Z�?��|�}!ӆ�e�ٌ�gVi��9ٛ
�q����� �W�^8}u ��9�!�-Mz> A��{�i4�Pd/�X�5�ݮ�z�5T�GjaT�$��+�Ix�� ��Xⅷ��B������,>F]�q��dƌ�?��vh�|1�Ax��&Z�$��)����|/s�+����l�|��s��(b%dn�S�4���N���0m/1it~>�'�[(Z��n�Q��0�Ѳ�P����blIܴmtMaKg����C3��D$Iz�˚�!�������l�sFb%���i���}IP�Go��!�/��EH0�[���#�"�_�-:\D�Q�:�Fb��i��5rjk�XfZ��D�K��qx�5*�{�kQU�5Ix�	t��Ɇ�mZ�%�(D�3D�IZ�>��p�Ǻa�2�7���ʁ�6�(�����e���sၼ�39'�S���(ǞVq�����j�,f^��	�c�j˭��Dk�)���IX�m4a����y�4�<A��5C�q�Vmr3y~ �dy=:�g�i
�MN���#?:m �N��覀4)��)�IKQمv�����V;��7V(���`�x��_ؑ/�8��{t�a.���y��}i�M�7�S~b���5qy_���.?�85-�_��R�T���ә�rn��(���GCTi�qr�6;��N�rC��4۩���1�5�Ŋ�)m��`q����V�0��(B��BJ�7��Wk�����ځ�����\�[���|�M	�JA{D29��Q���Q
[M�(���^m>��N��q�뗉hٽ�Ah�W�J���.�dOH{�����fV�]��8z����x��g�Yn�*t�H�͆�̎�����]����-ci{�G��[��0�~~L�j��n�?��jz��F�9z���/�����~S��AU�=��=�dKJ_��|�|s~?HY�j��Ar��&�� F�RbBf�=�/�(2ܑuK�y
L�Ԋ�����v��[Ƌ���J.�M�h��� �?l.�����Ѭ�Mj���Ow|S��!��4�n���ʸ"��!? �A��C����h�l?wP��l]@~��k���hz)5,��_�G~����� �
^J��j	�7�i�ے���0�Eu�,^m�щ2PZ15;\����:�X�R�c:.�/h��ؼ�pd	���Iߦ����l�E�Q�j[�C��M�냔x��U����2ʍȼ�F
^�*Cϩ]�O���AM�#�H�����9s��Nܨ��|�;�D���]�`����Ճ��_�|�F���u����帼�=2����I�xƨ-�O���#L��EN��r��4��-0�N'���Q<�����FZ�:���,3 ��U2�zT����]�jw�JŹ�yx��/d/${5��$fg͝1���6��'��N4���P�rO�b��29��H�u�)D�|aASڪ��֨p�0B\���� ��2�@�u�RDsg;�G��n�`t�G��_	�o��E�)���`��V|����� 8�i�о���B��e���sH�(c�yթ��Tş1��|�2� "�׷d�BW��ܙ�ͤ��#~�E}4,4#]KE%��"���F��)�-j9�1�U�K�pܸ��������ZSFy��J��Zz�{I��B0���M�Xvn�D��2o����Z����K���	��,]��G���F��@������tfR*�:�M?�zɒ���t,e��-3��i�5.�m���-
�f�S{���lr��pV�;^x�ci�E�Y��#��i[y����Dּ;"�sI}O�ڍe:ژd8%m7�T�
�|�+��"4`�
cjHZE BӀ��5	��~�L:��{��EL��_.�x(���jb�n�3�}�dؘ)b{��0Hy�/�9`�����Ο���oIa�I�"`�`MwM�͞>�<HcW={���1ьE�y�#�X���� �7J>�Qw,�d3�)�B��!��8��	�v�3Ϩ�L0��O��͙a]�EonGI,qW�9bJO�th�M��>3�c[�q���˷��9�y���$�b�!ɥ7Q��I�8gZ�$f���%�R��~$C���So3T� �[X-;n�z�s֌�XҙR�`�C�s�bs�KLl�4T���-���G�N��]�)j=a��ֽj�?k�$�B3�7<K)5��5��a�RM˝:>֚#��Tq`��mqCA�g��:�_�C[�"B2������T��w�-�p��r��e�E�����l��L@R�����d�B��[q����{���)U�^"���/��/��Iv�r��g�v�j�\J�pQY�G���E� 
s:�z�7��̆�Y���>]B��u�	�y ï��uP��R���(��4����<������"�hWHU�JE������+�݋�YW[�Io�]uo��]s�~oΝ�u"O<�j[�����:B#���[mI\��0Oˉi�C�
�2H��viA���/f���AI2qv�2`1��&��y�����,FV�_��9Pl���jW�SfQ��uJ��Ω��Dj��͙���_�pc����]���'��߮g���2<��B~bS�xM�l<�l����,a�6ǀ��>��s&�L�Y9n���O$ve�Ѯ���q��ቕ��)��YiŞ��z���û�R)S�r>a��&��U�7Sd���� ��A��e�bJ@,��DO�	���x΃:0P�����O"B3�OR|O3�d'����!�����ͦ��f����1���P��Vq0�nő&G�v�o��F3$����0��	�Rj��^��s��2=QF��`s���+����q��� Ub�e̘n��hxɿʽ>'�<��0�<�uᵏ�0F��������ƞ���H�X�wd�Ԋ�m)e�#�LBh���3}��b9�B�x��Q��Xs�%,-2e��g��M�뽛Tl��B�z��H���Վx}�#Z�O�����������z�9��ʘ1)Glh��s����t�G�MO6+���2���'������Ap;|��� yQ��e�N��Xӵ�E�>4mtݣ�wZ״�ꣲ����{�Eث� +����}%Rsc����Y�EF�����3�@֨ts��5`d�õد��j-[J�r��{#]�#D�X[���� P(�>��)��P���LV��ꨋW�)^�&���=�CF�V=�̉s]nkҠ��>�2.����͗ԟU�o��������2�_��l�{����H>�?���N�+����R���VLuM��{l��4QPĭ=9/�������=�i�g�-}�up�a �1�ݥ���q/n`��Y���X�J�ɵ֛�'����c�'0��t��w�>����ɚ;��5�F������A̡�媟8c�n�bgC����� :� �@>�|��ـ��H�}T�ɍ��[����U,�$�N��+��oU�0F%
�l.�U�ꀖ�~̨�G2�;��F<�m�h�/�Ư^�c�:=iĔ�������]9�Z����������Z�u�M�U�����Z��i�o$�p���""a?�
�� )􌖌Yy�k��@zC�VP������&�-J�C�<F[r��)52P4���M�}V�+n��]N1Gq��1H��7"���������M��8Ͼ2���a�>��`FZn��4��*-�Ō%��yk\�J�����k���d�����2�c3�a�j����ĭ�K-�n�#"�B�s��,����v���y��}�+�rc��-����'�:�{]��1�]n���\�fGH�l�.ˁʭ��,	�O�s�"X��8��閜��bu��Q����A�AֆD�����x+%������Y�R�έޢ��F~�#]�E�s�E�~��&��+A �A(BW!7�ȫ/_;k��kT�]�x)ߓ�k,�T�X���w�ډ����i�{:g��@>�4�P7S���)�엸
�
����7tY��骺�����@��`��ޛk�Ir��]�z^o��ʽ��|��J،��%k��?��ٜWB���'��x�|rB�y�o'�.�5)o+�3%�;Zf����gm��F+�d���NX-�g��4����AL�P"X�,m����lz�l�>OẀ�<���.!�o{���-,��o9���՝K�֋��x{Jm:N�{���P�3��G�'8�&&f���$Q֭�R��;{����S_(pT7ͤ�nK��$ �����")�:��2DR�8��r��5�]L�@�v��l#f׵a~f�F󶲓� �9T5DT�q^�i}���br��n���d3��c�9��Q�5^쬛�i|�Sƭ5nc�6��cJO$#���+��i-��!��������a	�B�f� \��h�1�PuT[E�և���]�\�'����oi�	Q��=�5�C��{Gc��'�J��F=�q/�`��o���ʁKk(*�SE����j�׀5�h܎��fy����T^Du�)f>�5��-Z���c�)amR���n�*��Kw7���T^�u�J�,4fQpWB.�A6@7�"P5\r�'���os��f�i��?�/]�!�&�l�<`f'���Q�&�{jXT �ʦ���(�g��S�Z�cJw��S����1]>M_�-�lxBI�*J&�@_*B�	�dS^Gg���>ze_�.L��H�3�CP�:� ��ȷcU���en�A��5�c�қlE(b�K�N�+��8��3"IW�"���葑�#6@ѷ��}�ZPH���3���r�Zm_��(��%uAB�=I�Ô���8+6�o����J��c�k�ޒ9�B���1���x�JJ��~o���;&>�{��64��z��L��z��Ԏ	9(�ң؟�{7�s~����ߒ`.�K�㛪ζ�Y��um���l0p:
7p:���S�|��rU��hݐ���]#��{(��х��f�Ý�U�ڝ*�|E�����pGd��TuU�U1�
�\���W�<O�Y�F!���=��7_�Ѹ��+�(�-'��&�	��ň���h������cڮEX-ꌀ�2xχ���\kmQ���]��n���{1k�a!�\dFk�(�wܕ�Pğ����>�3���i�K�J{�|�wo�x7BL~)���u ��&h9߻.ߝRc��1vɒ��z��h��OO�J�l{��[�9��RZ�yI�J�i
>�r�>�v$`h�U��m���gl�N����_S,^"�|��_���<έ,�W��&����*��s�|>���6E
G�z�
�ӡ�_��G���i*t��g��C'ܜ��iY�M��j>�;^X��F3�iff�|�Ld�3��45S)�)�Jk�W��A����7=n�=��{Pl���� ՜��I��S�&�Q⊄2�>�\��I5v�D�׳h�[�7��L�z��	zm��O��5|:���A�I��dm��<V�1��Ժm�t/�`W��+�ߵ#ī>|f�����ÁB�T���)/E�l�Ag/�.Qq��g���%-�[��;�h�PF�,	R��"Q�X̋�C!W;�A�RA�4JH*���5G���t zy�~QOnH�m�	���pj��^��I*j�C��ֹ֑���V�����zL�7�t�*��.��*
~��\���8\#��	��ʪ�j%��p�`d�K~�䄻q���*4Y��F��'�n({�fq�R��c6l��.]>��������6S`�Jv�������Z���Y���2ۯ�j\7e��G��o2W���8�ed%8�Iد�d����h���@�6��p��Dn�[�"�i���2<�:�R�� xMJ�'��|3�Pt �0z�f:��f���lwx&��o!%��If�"�y`T���i�tݮ�9	ưC���˛���3�m[�)?DK��$����2>u
��OF�e2~c�����)���3��q��_������pc#��8,�4�ʨ�'#ђ���s �s�������}%6��v<�wgU\;$��R�"m�p��!���^N$�ىV�����Bᇡ��W��B�GnV�
�`�N`Կ2��ޔ�y�����ׁu���o���a�H{��*�+���b�q׈�}(8}@�1JaV�;*1��}���ٲqQ4�6�r�����6M8G:����Ug����g0��B�]"�Y�i�^�}���E+b�C���W�y+��K١�3j��o�� ;j_��|۶�Q���GXdQ�kz���j����?���3�RˆuX����-��P(���'�tj*r��ܫ���s����C��g�����?9����N���cɯ�S"���H�B��M$���}A�|�BD@*WΚT�b��U %@U��=�p��EoW{{��ڏ�$�>�
f��|�B�.Y)��#ܬ�On�ݡ�bs����P�xy!^J�_̀"R'3QJx��>��]�����e��G
���bץ>�_z�>���$�jT�HB?#o�{桌_�{!Ot�h�Q���O.��;_D�}àk5��ػ�
�<1B�k@��7��a�ŌQ�x��D굝Om�M� ������B����7اB]_����h����*�*K	�W�Μ4qC� �c�A;�1T�l�ƅ����Q��Q����Թ3^?-F��6.9�z������
HN=�d�~,����s������+x\S���a�[X��Ulko+��h��[��!ӛl�<%Мa	8*�!7C7=���tx�L�T��O8�򏪤��M1� y|'�M��δQ��Wb�Ya�x�G;�6X[)	wWBz�4I��(�eK�6�@�y-��/��)2��D��fi��+�I$�YYpS8��h�����J;��L�������1��Ǔ��o�_�[���I���XZ���x-g��H��wnβ�����epM�7����xgT<�t_��I�U��u���$�X�NU�;ײ��'��_g1O?���X����d��PQ��, .��E�M<�����$��\���\��D5F��wr�zĥ�-��ۑ�Ȃ�g��{ _8V��q)؎޶d���֔LA�8��=7 �p�	���݁��l;���	��,�A"���a�������~�V�$�X�3�a������>ㆣ��Q�J�)��Š_]{=��K�P������5H䴦Ň�Ŗ�K-�A��X�T�j�6�{E�p�X�,z�qr�:��$����ak�R0A�Rx�PŹ>��d�ߛZ,N�v����F��ƅ5�̲ړ���!Nn8�P�?&���9%��k�p���8#�]������m�d�����h���#;�=���S�����8�+焖cJ��^\�&4p��Qeh�؃)�Um�
�ؙ� orz{~��Y�_��g�1�m $/v	Ȼ�4��P�T	# �h`�$����N��Z%�6 ��qc��@�A�h�pC��Gm�M��0�-�����tl~4i�� �9��-��W��3�����5�DӃ��)����D	 U����@�N��a h�*&�"���O����&)�"f��[�E:c2`.o�P�zb�_�kH�4�����-���|�Dh�L��UlaE|`}��o1Ꮼda`�E�;O��p��&�
��#��!1�:>�`���GC��H5J�˩�L�l�2f�;��<��r�Yh*�,s�?A�2RB>fz�>���[�=�?~"�i�+T�������]4ϙ/���'L���1h���J��+KJ���t�cb������F�G�`�t�A��:1�	ҰW��0�
�}�����ן���.��掕���-C5*Ȱ�8����-!�CAI��	�]rud��z��J�}A��y�n��$9h/	���T��Mg�1:�3.�'%�9P9�[Is���l/w��J�x<w�_u�H����8=�Q.��e��������J��k�M�.�F�*-!�Vb�@�fC�J�^���ىƮ�:[R.�h����y����Ғ2)�P=��ý�݆�~���>/Y�ܝ�K�"+c����˗������j������;a�.oj7�qL`���/W�3�*p��,�h&	$�d|�Z?��XF�a��
>��_���_M"rb(��=M�zZU�($�����1?���H�Ͼ��1��ǚJ��'���,h��?�oW-�z_�jIN�\�ف�f���'�nK�Y�����`�Q�or�ne>�x=�NZ�+{��<�\�ǋE
�k�6��m��_§%��K�G��}��-ϟ��u�I7ֆ
�Ȣ��fj?9���_�j�k3�xI"N��oM�l��̇NljxYy�e��"� 4rT�X��7��+�]��x���RN�W�k}�G�ZK5t=[�k�-8��D�������g��x��hA���\~��F�Ѕ	#�)/@{�Uu�̍��X�c�5�{���B�����z��aG�\��季1Y}�X�O��k���vW�(�:�B��zw%P���{�*�q]  �h��6.����F6�X3�Mt>!�L�q&��=��t�[���q"R�U����Z�)����@��{ӳ!=�A
�в��fu,vH�:��$�;�G-�[o"�ℷӢ:�pk�gAc";�+ L4�	��qhtu�����GH��q.�������fX�y�ڠ�cSWs�#L:O\ot�]��/D=cb�b�By���i�$���[�7��������?\�3\��/�Ӫ������2C�������	��h��
���{7��@_Z�D*�R�Ɣ�&"���ĵ�ȗ�.����v@h�6�AsvO30XO_��/�0b��栏1�[b��)��W��Ci��b�_�V2�1�-�sr���)`2�0��<��R{�+��2�@P��gO��#�@�'o�Λ��?��3���6����ٙ{.Y@�"�$i���v�4 ='�CQ�N��j�4vI<�S�x91!��� �õ���U�宍����i>�wќy�Y��?�Wpql(?�'q�/�w?�!5b�M��z��^�?<78�5R'O^�I՞�1��P��Vh-� d�mN
<w!�`d�Um�¥u^,��9X�U�Q*v��qI�XE�ih<�L��Ө���d�A$,	q
�r��liMo=�I���u�)7���)K��~W�tEo��F�l��%~�I�r"f,-TΥ �_���3_&K�D�ɔL�|>� �8�Z&���uN�]��M?�;鱡��i53K�g�3՜�[#8/��ڀW�"��_��2�4ܢ)ǄR싲OI���8�����G��J+HL9��VJ�8��p��-o���^F(i�*V9�8������t��/^��8UI�s�)����'����w��5V���	4'�[䠙�S|[���J�Gq���	$���j�@˿p�\|��6�xO4�Taǻz�1:(i_�y��)K#��ܺ����̓�q܄��ǳ����f�$��0��:��I�"��}s�= ���lڼ/&%�ŢV����չ�&׮�Ł��!'P%6�-� �s�*&�52���0A�#+����M�T�6dZc�GrJV��h�����^AA�xa�1��FC�vC-��P��$bpq7eq[�%�n�}�]�C���}$8Il�_@ߩ]W\p/�>�	C�c��X#S��r�9|����E=���.��)�20�^A�71��[G�Hv��T?QB��|n��A�N%���|��4�^�>���.��)(�<��ڲt���r�
�C��HI��qƕ��xB{����J �����_�8_UT�l9��L����:��@��oK	e:���&zI�f	g��X}�۽ҧ�m$���Wb��^��4��g%5�G6(�-˳F{WO�����ʇ��:kNTZ ���6�T��%m�vи�J� �_�j�N��`�ĀH�B=II�X��;8��֍�Oe���X�͏*��t.B�hRx_�2�2_kG��)M�����0қ5������N=�]�K����t�\��'�IVt>��í�B�[{vV��C7�=A��/��/�Ȍe�P�z��ޝ�����H+��@(�l>})�'2&Y�8��>�oTG��.Ĩ��!�흩��yϢ����i����L��H�/i��)�s���&4��灝L���Cj颍�x��R��h:�9+L]�*9C�"�	��u��;yU��N|a}�mH�R�x �w��:r�+��X	0t{g�Y�E���NNz�� ����V��24?����0�*=�*�6�;F�X�!�9r:�1��O������ ���׌���fg�-@.��z��݁�?I��sc���UXˢ�{�0��W����AD��F���-I���1)��x0]�wW\�ˉ���h^P,3�J�c���59z`���?{�����|8��?�IGY�$=x�2K�����a��aJ���{k)Z�RY�w�k��R�L/>~(X2e���'޹�T���pF��,�-`�3� ���`J#ά����E�[�cj��R��������7_�lR�,R�}}�,�/�����ZL�Aݐ^�Mdxj`S	T'��^́ �S�U
�DG��FBN�e�9��C��.G���=��]��b(Al����?�K�@6�{�wt��9�T��������5����t*ANMp�v��Za�n�a���c(�@`Y����?rLT��Gq/}���y��u��|���1��Z�c*;'�j!�)DW'B��i˗�kӟ�{m���fN�>��1ߨ�c�.#��b#w�R�'���j#9����FP��V@eF�6��LW�%�,|�@nSS�[}���2Ё���Gra����x��
�
`A��=9����8�6��y�9�
鯧ΰ�]0�\�$L��03�1LO�)A�C�_�.,^�q�d��I��͍:�pͅx�j�sm�*8(�b��yȟ��\��a-������+���s����JaA�دK�L6k�zo4`���{1�	���Vte���yaUU�.�'ײbeP�޸�]xӥ�9�<�a���09�0��b~�ctL�����Pߧ
�b�E�gu`YmٻdA3S
%yij܌�6y��}.Y�6�i��Ȼ�yW��~�d5R��l��J��>Di�(��#�:�"����F��r���7瘣u+�&82)ȑP����1b�7����!Y��:D��s;�Ѣ�\���t�-�>�?K��<ބ�HC�m �����Xxv0Q��B�G�U,��R����ڤ��1�����rYu���U�u��{3����6t��1{���Q�"I[l���,rO��9����_bc�[�*I{�闫A
4�g_�D��E��ȇ:/FAfz?��$�-�Ӭٯ^{�!���'�#R;���ّ���)�W&h0j7WTۡ�)�: �_R�g��@:(�p��p��m6���4<p^R��^R
�0S����^� �PC�+�}�81��TȈ�õ�*쫒$����35Yt�ܣa�)�����\E`��{�_��4w �M�n����v�>Ĕ!�ˮf���F�����U�".x+��?�~xE�ݧw�wf˲�<S�� �M�$�����b���;�9;���6:��7!��I<J��W�!�FxҸR��)���j�1�qEv�BU|����/"�Ԟ�9���f�Ck�\>m�|y�tJ9���o&���\�׀�I�P���^%��q?"�f8�p���F[�l�2p��iF��*�J�o���_�5�0
��l�tC�I�γI��K���.�Q�L�kPE)�c�D�͵L�'%[&���f<VZ��*r*���MYmiM�,����c�ޒ�y4g^�{�r����&�ۅ�����,�#$;%���82v��a��DK|��x`����V��y��4U�?���_r�K"�D���6`����}���3�s�p38.֖7D����D�0���ZOU�u7�E�y�г�y�h �lCrs�����5�U���jQ�F�N]HP�o!�6K��y���P ��$%W%7��gRr�PY�ƣ8�P��Ks���A���f07w�{���4�})��z�h�Z:%�y__�Юͺk	mEM�^.9*4��{��q�-J+ls˽��^�����9�8�@o_hH5t��Vj��Pe^��M�P^ 	�Y|)��Î"�K�yӜ�	�Dg�|{���x���H��k`�-�G��84ۢ�W��ef��L�/1����=;�K7�nE�p�qem��Z��*�5�[��_�����سk:�?Ľϼ���d��O�. #�v��D�!`O~�m4voOv��uI����%�JP��OsűNw<ʖ����1�I_�v���s���x�<��4l�h@ɺx�]L��+!f �g�q��B��b{ARᇁH[i3�Z�J�qU�3;c!1��֔XB���Q�L,. �	s4�*n�vQ8�}�N�	��|�Z���9�4�̄����{�	)�7iP~��t9EZF�y�x�~�S$'�F��k�����$��H4@��*�b*`�:e>�N�(�M�Ǝ���J
��L����
�.��U��!��d�5�>6����baZ"y!.`��^�&x�0��@����T�l)��$��黕����@c �#ڠyY�,O*v��w�3gtQ�7.웾!�Oy`'���_0��#)����L�9c�����e�4_^���� r�A
`��̒PD��|!��3~����+��\܀Ac�>Z)j���fCW�(�Rlf��I�&��f��ɼ��Lo�Q��i���c�R���1�K�ɶ�|� 4EҽpsD\��lN�>��Ç�X9���b`�V��i~&��ۆ�9�@�-��=�9�U@2��o��KS	.-P���ʃ��9�O�vΔ;#'ދ���4�9�8]w�H��XcG���+�W�<�P���w�����㙴C/$�XP�6��1��
{L�#p� �����N������{;�􏤽��IO6�:!m�_3�X�(Hl=i�R������Q�dFD}��<��Y���,����蜑h[w-]5F�^�i�YR���C�����M%���n@�t3w��0�f�+zo��@�v	�ڽ�,��:z� �u�(w��Q6���9�3�|	Ws]�O@O~���~�Z��	��%
è<[qr��R����U[�ʖ��[���'Q�h,�6&���f$cút�d(]��՘�"�$��4�.��7��nV؂��%Sev��T-Ub�8��8Ӡ/lS�B�'�<����ڶwǌ��	�|C^�`enY	�EGǩ#\�\�:���pJj��M��E�Q�h&�H�+f��(�Kֿj���]��E��}/,ʲC�9�� W8ǌ��*�5fT�|���{�ݳߨa�J����;�����b�G�ȃS�$-VHJ�8#}Amj�@?�6D��D����f g��R�ݷ��HD?1y��a.n��6ea�d!��U�s~�`��_��hDe�}G&��fRgn�G��m�[Pe��\�W���x_TV��J�c�eU�n%%�|;+F�ݑ��	+�h���䡶e \�Q���F�ĩ ��o�҆Ԓ3Nv������r��*�ΐ|e�="��U`�IT��Ho�h���y�:s!�G�0��9c�u��z�����7�/]�G,�Z���U��Ǵ�r��Im#�O �b��.�"�}T�)�^�#f�7��},F0q
E�-gYاx֓���%q��fjYR"���J�����@tOV^}��G �93�T����4�n�����:�g�x����Yi����O�xK�[l���Tw�.�����CU��0'�`��!2-ϣm��v�:��T�qe���I�(����w�!I���sa�φ{�J��R|*�P!5��Ss��Ԓ��T��$A�ɽ�Dg�U�bf«���@���;�T�1h�'�M��%���m	�����|�#��`�m0̺�a@[�H��"�e��uɝe?\�%�7�j�c�N�5�x7dg�p��_'ʆ�Z2+�?�'��P�(_l�pc�fWh���}�B_���5�7U���;���&����ѤUF}[�pqNi��o5_�g��$�!��Ѵ������7Ve�<g�6�ǝ����6�1�pDSW@��觬zB��G��҃�}�y��w즩�j�����.�B3�g�q�P��E���a�������c@��V�W��H^�HSgkh��?��*簼5\PL* �m�p�)�;�Pm��<'"/Ώl������=h2�X0�W��_�[弙z��o�ʈ�'����Iu'ȯ7�� 欲_Q��q��_3�Z��~��@���Ϫ���9<,�w����Ĩ�P�R�6n�j�UU'��o\z���1,��%���2~q:JN�⟟�m�դT����8Brl�=���P����:���!i��Y�>d��}��j�l��To�ϚzAW�{�g���V���B�����.K%X�s��n�QF����	5u��Ɯ��?TV���C��]Ni����|�pj��VA��O��qR-%�h���)��d���L���`NvQa��4`!q���y��A-V�9����xo0&�o�(��oR��s�ɖ���H�ӏ�Un��צ"�����Ԣm {7g�^*�2V�r8�ʂ��*3���W_ +��PJ�͘؛��;}�mO�;�-�&8�HG~b_C��*
�_�uN7�J��D���E�1z&񔈿9,�V����h��}��D�k��n�m��w�ꣻ҆)��/��;��"��"��aX���F@�y��R�6xk�����4��6(�醲�X�LX<.�E�n����޳�Do��X��n�E-�p��x��*n�ۆ[���(�}�is��;E~��M���q��A�՗��T���Zzk~ ��2S�G�V��l�� 
?�r���(������P�M�(f�_�����I\[a$y�t2`*H��}�Cn@!�m��f�A�^ʱ��]w������U���_��v�US`]P+��ZK��y��R��i5��`��<p�e!b.]�.Ձl��"�s����C���� [۠G�ǳv����-���M�(>0�j_�U��F>�$�=u�(���)�6���KdK0d����2A?�]�)�1���QSBh���;
v�0Z������B��<���bEî��[��Q��C?�d~�j��~9C./�"�5�-�_�FY1-�f�I�����y�Re�bk1�^�)c&���������<6`9���^\�<���5\K�D����m*ͅR~�U�:�t=0GXj]�{�T�-_��L�]F�K޽"W~��3�� �q���ז(���Y��p1���L_MŐ���RE1�9,���]�i�d�����{b/�D��!n|9b��Y��'H(�1x�Ϟ,�fD����s�l�������5g�gQ=�0�a�8�g�mea>�'���� ���msa
�j�U�xّ��~�	��V47��dZmz�®,��HAz����G?�`{�%���2������Ō�
0$��NE�������YS���������x����.=�#���C�}�s��؉�תHBS	�y4��Bò�Hmm�so�'>@$QA���u]����3��k��e���)�%� �m���%d<���`�v��H����:[k:�9ƽ'�v*}l=��H�	�|�&�A��ĕ�vh�M�%rUw�u����֊�M㽁���iӞ#���/]�\��^=�,w.$"j·�lE	��y����2��!eQFB갡:C�>��|{o)A=*�Iqz�?���L�_�������b���Ƒ9'p��d�(/���>=�/�����|զ���1>�LX)^C�	R[?~
��8�;E@�3C��I�I��@�_'��b���LPܮ��Nf?.���M����4	��D�
l2��?������BX�z��d8����/ie��0ʆS���0��}h0�x���U�(�NµK�b$�l�G�ߜ� .`��Nu-��y�g<�2��	�h�!�b�PFz�Q���я�Z��܉)���q��V�ĺ�Y}TE�(�\t�3�h0������$8����݉,jMAu<�=�~T�6��i�"��Y����/HԖnѯZ�4�� ͉խv4 ���6���n��%� �ߺ�<S]�)�2;�V��y /���z�m���8�J�`3�!YΫ4��SuH�cÂBO��%Ck���M��}�,ЏB�
i>��b��,4��4��lQ1U�Ӑ݇����N�+Ur�c��(����j|��}�q�+�e ��)�j�I2E�����yX�AL/��q��g�3zߓt
%����������}?�^VĆ��{߯�I�w��s2�z5V�_�U��U��^����d�L�q������)��o��y=S��~�_/m�u���k��F�&��~>�x?lm�1"�f������JV�un��fk����t�	F���H��Jb|���{�%5LB4h�$�p#|�
�(w��**6�P��@�,XPa�s�T>��W�q7�,1 D�'���l��Uj&��+lw
����>�N�r��YJ5�&��c�7��]OR�p���	��
�2R�i-���m���ժ�)�J
��uO�]]D��SgJQ�0׹
��TR�t�N������)��(c��	�R�m�ʇ"��� ؝�4BΒ�L:~�}�����gY����_ׯ�9�(��̡�v
ɜ���_��&�b�b�;y!��bO���8��]��K��m�B�
)�Ҟ�Q8�
9 ���`�R���3��� �Ύ��Jw
\{l_!>n��7������we~{�����~�J�����n0�$)}Dw\X����C�I�m���Oщ��s㋡?�l��'>$Jgt���J�,W���#�e\�� ���댦5g*�	>�z�ΦHr�]��î�ʎ��.u�Td.��<&x�5�W�`�m
R�|tF�U]�(y(����C����~Bt�hg��e[6�����+�ϫ���L�z��r}�lZN���>� ��
u~7�hn4��e��~w��-��5�0�
��@$qQ�������xz{�5�;�H�3���ԸbD�'2�8�����Vҽz�KU�Vw*���Q��'�9x_�����V�q��uoq��ܬ���^M�<pJ]��]���)��>�xa��K3_���&���(��OJֽX��$�D �2e�cD���M�a�5��c��������lo�s�̖*��t���UG��U�K-��>$�4��%|��%����;��b�~�X���2�s�&�n�㿑=o.(�������@�������\T�B{�>�{�v�6(�v��,W�z|9Ց�r_[��������ȥоLpH�x�d���2����u�4�0� Y�&x�*֘)LjG&:s�;�����tBσ����N	���¾��d�X�<# ����zcΎ�Q�t�22X�����[��&��G�]|�+R1E%��Mˊx�w�ٌ�$�����P&��7'��<]S�y��B�B��sT9H+���V5 Ewxe7}�t�/it'���u�9��	1�+D �Mԅ;e����-�A��3H�NPٔ�[d���_/R"j!3��]
�������p�э�Ol���߱-�9�&��Γ�4�C5�.q�,�u6�0�b;�s!�9�*���Ʒm�����"�����R���L=�mu	1M�����];i��ܧ�xA���Ͳ�3��:ښ�R�ԨbP��&!b2���֖�p]�0J6�W����N�Q�H�յ�{���?�jÛc� a�>��wu(���(,���'pK�tu�"�;����7�D㜞-%j/=���ѻ�����%�H%p�#�VǱ�F�:�W�����?���J�e5��Vc����Ѣ���h�&�D���N�;e��������%��d���xEl$�Y-Yzu�]
�z�Zg�y�}\%r�wŸo�b�#��\?��3�ܭn=��}�7����^�9ɩH֓H���4�[��P>�<�q��~	~��k�[�F��c����0�P^�M^�cѨw]z'u�����#gV��q�Gb��	�:���t��G�L�<��Ӫ�V�As����Z��OW��K�	�b
\D;?p��	��zJڤ�.W�	���L�U�;u}m�K;V�6��GZ� E� J4��%��Zz�
}%g�6.m�n`�A��b�Y�.	��~�)b!�t���T.#�J��gE�˹ jaQ<�ꧡx��J�G0k�9P3Є9b�9h��@��RTE���9��6��*�	��C��'��j7���*|������.����Hj��; )
[��G=�1�V{�8�!��	�w��#
�v�q.���e�ɐ���=8@�V��܎/4Fė��|anZr;R��,�(C�]k0Ud'���*����s0�^���d9�����(sn�Z����Fe�:B�dW"�f���Ps&Jz��~MF����xٻ�V��\�J������dy�-�j��5'����6�ɉ����\�x��	tuW�6��R=�
�����挻D"\���}�xI{>��w*Oz���ܕ��>��7�0\��SjC�;�٘ć���N���za�q��]\}tS�r�F��� /�s� Y��`jf��xS�MD���5p��dK���Ҹ�dy���i�if����5����&�ES��?���$���\�TX
Ǿ�1�VRI�>�员�/�h�Kd4j�DF�V�)��&
\�k�XL���aP��^U�瞟��%�6_�>%j����m�%0<�w��Xԅ,l��;R�E��o8)1�)Y&��4su�fҀ�|�� H5��7�Ԡۥ���URҗ�u@$�=�+���UC�.k�v�G������������F�a�؈��[�y�^t�j��ǪB�@g|���L&�C5i��\���f���'s��S:<g�-��YId>���fpx~乳��DT\`��O�����CS�?��0Q����8���/�S��~��Ց���:��k|�� ��c�*�cO�=��`A�����e������D���ծ朹i&�2���-%�9�z=!P�gE���c�8����-EA�K7� ﰸ�lƳ~��,��:�=:�}�қ��A�~�V�0ZR�Vp��L���Rس�r�r�60�E]��!�uCp�����J��.�zm�~�*�g��[< ͞��q�����X����}��AQ"�!\������}p &h�|L�G�\|ē�����Hř�'R1���'Wҙ{�&Q�c�M���sôb�b�k&�~{M0�	?Ń��ji��f����=U��3��T��4)Z-{;�nW�+�L�s� ��-1ڊfcbBVxdOk��U�ŚffU��HY擒����_�F�}�x���o���l���A늉�s\��em���7�,��UtGv|t�{1/eο���i�:1���D�Us"h0q+д�M���S�fdҀSpeѕb<��w$z�M��� ��^OZ�r��Dɩ��x�^��5���h>OI
 �Y�@�4ahÖ�]�@ޘoBל$	�t�Kn��B���R��s7��v�4{ξw�v�N�v
x렞]AV�s3�����Ēw~�Y;[*���_�z��>oc
������,��)7. ;M��5���-������Q�[��q
�����_�?�Ιb��Z���
r@/c�-~�m�ϧ����d�0�^M4�5�8*�[�1�B�~��dk��J��C�/�z��,X����'���YaD�������k� {�)�D%da��ݭ�$k��!B�Cp8�R��ĕ(�%���P�b̯������kg�W��b�4�u�_Fj�1���Y���O���R�����4�� ��햒�xC[�kAyæ�n%�܎酜p�����N�׀@j����UK�n^��������t��cxQ�[�\�-�
� U��n5�'����!̦2��s�ۍ���{�K��ؤ�Ol��,`��$*T\��x�� j-��{O�����@:_�a���Iq�	��-wY�q���_6Nx��L�G� �t�P(mZ�u��C��:B�ۅӛ-S�`�����6�ւD��n��x>�_���w�4T���$��G�����KA0���)�U��ܰ<�(vb�4eI��D;D�?�7,8�����Aj0-��הqi
{�N�j�I����!�5D��n6"!Ga��rg�<{���0�O��G�rH��U3�*"#XF��:�&��(K'���k����O��Z��G����i-��d�����"�J{21Uh-ǝ��"���x���i㏙SK�t�P�q�����7�ʵK�5�'�@���t<�5���2-�`�t� U��m9���,�y�د��Q��P]�yd���_���0�j�6im�	H�j>�����˥o�%	��CP�-3r?���.<q��0H���=��>���䒵�O�{*�/��6���]��hֲ��W	9q?��dbL\Y��A߮J��DW[=�NR�u`��_��� ���,�Α���,���ý.���&'�?㼜�����Y�
�GΕ�.4=U��aJͼ��D�Os��'k�6#�ԣ$�x�0Y�Nq��#�	n��(�^�̉^,�-��0fқY������ޗ7���K���W��G�W�[�]M�>]����g��EML1]��]巪�h����[}I��h�<���3�Ct���82��AW���㒸���g�YS�W��YF����V�Ý9��������|��ᄮڹo�P<rɭ'��Bs7�ܤ��(�c�	F�Lȑ�#���_*�l��X�	*��L\��R�*:!�~�aV�T1��vV{�U�g�eYH�0r�.AS��7���a�L��b�E�H�2S���W��Ȍhg�zen|��ޅ�>}E �m忨c���H��n��L�$A�]���z��~v�(��iy�R:����:���Zy�'Z�̏|ݞ����y���ڛaۻy�4��U?3+��>k�<T1Ba�*�L�ԕ���#��M�i�K�?y�]$�p[��T�X��pz\>p&���ͫt��ƙ�<����J�p�6QDVW3��P�%���|s�Y��´���#���j*{���E�� jj����*� ��Y�J�Fo[w�i�
s��� F�D�+~�i��t��Y���,���:��P�������6P�t��k���!\��7��I��؄w	ʩ||���9݀B�p��"ɹ�"7��F���FM*c�� )���g���b�	��хQ2QdY��b���
� R��I6�V5Bj�zO���(��܁�%��9�i�pXR�4�(�Lw��o%V/e-5ۉDm�	�A�2��RY�4���b�D��@��/r��&�w;В�y��~ȏW�k�q�$~axo��:�b&k��5ZK�J��m"��.��3�	�g1����������r�s��,���@�z�A oC�d9�hp���6�t۸/�N�4��aƒ��	�sǖ��ؕư
A�>�y�����5�i��
���Q�w4O��m\%���>oy�5'��d��=��S�7��L�X���+
�J��Y�d���m��Q�;��;�jiPrb�<�)��p���ݧ﵃��+�l~���h�Ͽ�� o���%�(�5�2&�R�=��3��Ǚ��q��S1�S�>��4 �d=��{)���cH�EɎ�m�����.�ܷ��@Og�\��/��h���YA�
���g;��X�>��\���ʐ��ܫ����E����s�(�ȿ��$6���s��|�rIbav�_6E�X���y��ҫ�]{�v#+�\¨|�ơ�rz�F�� K ���Z�oI��̲_�E����� �5\�g��ͪ]��}�k�O
�^�xk�}oK�T��:�9Zi��nF����>��u�2U��L���!�bڍzf���=ܨ�6Z��_�nV>�7���`~�8ρ7�@�{��wRvR�z|O?P���M?�QPi%��Y�َ2%�cLc�T�D7܋�d���m1�Us?��+�XX�6��1%�k�;8��2��[�+-���f��g#	�o�����1V�g14�u(��=0��-�ן�.yr&]���8�YI���Ė�,V��ޛ;1��1X����+@�s��-�w��H�$q�B����hخXD�_h�-���<���jHe��[�<N(�k�����c?�V΋���F��j�Y�I�&޶u�e@I�6�^P��9A�T��`Z[-S�B;���O��nW��t��޳w͹��n��~	�Wj�xi��d  d��ԝ��8@����ӳ3���	��H�,}�=��{�-Y:��J)o�X�& ��u�M��� 	9�+1Z�6~_�i;vJ�MY#c��P�N��CJ���	���J�mң����(s�Z�!���6��#���вh]�g)��AW�>,[�'�)-�Κ�MP錖���(X���5��!I���0�h!����$�@��r�=]��"U�mq��w��#;�Q����Y	Gx&��l,g��6�i,�{z`��`SF��w�T�,��F�{����8Ǔ�,�?Y��ɒe���eͤ���<]})t%Y�9%��-+�F��T�`�r�n�����
	!o�l8�!0�!X3���I�ד�@�u!1�xگ�hBf�|�N2�ohZ�s፮��\����i�	�8<���Ә�p���sf������0_ߔ�u�����n?�d5'�VrMJP�B�}���'ʆ�ܫߚ0[�/�\Nlv�L��1��Y��bD)�?�cTY�@�j�`�ـ�����6��f5�=�U�ƶ�嘄|��-M7(B1o��La�G4!&��yY�G��F��=�<I�w�	'<���3a�F�+����o=}<;�`$쒘k����I�H�=�m�?:/�H�D�-�PGS���3WI޵���9��|v�Lh�c����_�r"q8�����?��9e���ۄ�׈�^��>�3��t� ��S~�}v!}�	�"ߙ�Պ�y}zѐ/�OT�Q��W��b���r���C����=���l9�(�7|Z���j7����}վ���m3�	���&ka59,���T���Ĺ�g�Х�(28v���!{��U���z2�7�~����p�	3ʝ߯�tb~<�>sAH�%.�I[K�+8�Dg;�������S���~�.KTX�Ղ$���$k����Oȁ̛�\�.�(���R�5*�/:��Y��hdM�XN��`��eu�Z�� �C�=3����V�Sr���P⫳��C�-��}.��r}D�g+��[��Y!d�T�8�w�o@���{~~��C�G���N ���<��c�8�gTR��iar�^����=�n8./r-b���/_�>~F�Sl��!d��B�d��n�v�wy ��:�X\n>a��jV�Fԣ�6�' �2��7pQ�����p]Қ�����c�.�vC�r��w��'����/&F�H��8�4gh79���
G�ü�ݲ��g������P�o+f�v�KĆ��XΓ�O��NYӮ|�z���L��7�R4����/'
��
,B��b#��N�%���L8N�9�Q�:�/���WתR���fq����9_q��B>v��@x}��K; �f�q�P���΁MK�c�����*gc��׀��[��;��tll���{�C�Ƀ�d�2��7��M��(�H���zFp=ӟ��2�5Y	D@��?�<i�c"q�7�mj���,��s0Yŷ�f6�fy�5{V��[ڴ�YJEq�{�@3W�7#-j��8aCѷ����-ׇ2����%/�kUO�_L�u�)��Ae|u�0X�f�z�[7XS��V�!X��`vKx�xV���z�n�]/7��'�]�Q�1����X~�,jΌ>Զ����c��k�շ�L�L�<u��)a�㻠HxZ)2U��lI?��i��Ws�����/��X�u�R7@��6A�&���F�/�@<�\��H����Ĕ����qVz"�Gy0�r��d�A�Z?'���W~{��e߭�rFY�x���t��<8cP��Aߡ5��)�B�J�2��6�{뉻eN���-xd�k�.X�7d\���H�n.�e��Q3�gҰ286T��$����{�~W;X��P=9o�pp�. X?D�}��"��' �8�G�it�Q�8������|͐�죿�*q��E�l�S��y��r�k� �P�n��S��S�Me�,�^e�I���[���*��"�DC�6���U?҈�]h��xR�X��v?�)��8⪪VkR��QۖN��(��..ƽO�R�����)��l�V��d�k�S��L��YJ�GXe��&��$ApdnCdO���/+y��ɘZّ����& CÉ�;9���рa
vh�4�D�v�E��V�ͲW5`s���R蟼���:���n�ȅ.�ګ�d� */e�Fɶ+<�y,�4�=� X�-eA����l�ܳ0[�T��{{��%އ�`�ח]mP����a�-w��P��nV�0?2��n-��)g�n� z��a(�c2IȰ/b�8�d&��A��CI��\��-@�Ϋ��+�'k���)z�x缕�gW��<�