��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�d�]�D�D�ow�P��趝N��� �6�����.cIbp~����x�����;��[
x�|�'I2���ѭ�M��s�6gd���g;4�7� F�����2���J�ŔC]��1�r���s��[�j��B6� -���#��*��z�N�q��Շ�yq�f�4���|��la �0x]���u��T+i�.���F�n�ҋ��?�R �W��AaQ��>�ZW��ZXix�t֘5|L(wh��{��X��l*�i�X��+�����w����wb�\��ɧ���eO���vu����Ɂ���ϋ�ۡeͲ�nB�^<ͤ��F���F%��V�n�J~�z���E��{����|�G���=�>���f��$����sDџ�8�tn�;2����<�����td-$���Y�g�{-P���}�3�\%�ET-V|��>��07�@��g�.�4B�@��i:-�.l�̂Qs�u4C9�����W�������`!t'�C�3�][�x��$0;E;��sw$0�Z�sEj��${>U������4�e+9J."q��;��z܀Ǆ
�ʦ�z����ƹ�����
�L#e�˼����<%YP��Dl�KC�H����H�}�.Υ)u#��0��hP��A4��s(K�pb��d�aL�V�4��&F�A�E��\�;s�x+��`�� l��3��u�-ZA4�QX1�l��In�}虎L85@��Z����I�nW��`�%�B^Qe�{1ƒz}~����/���)��Ռ���i�%�Ã��� 7�A�n.����FP�s�;TGr��d[���T�]�w �B��?JiH�h����tI3?�j�0�Qְ��vQJ��'L�ŷƙ[u:�K��c��n�ɔ�xN���ju��r�3���n����	�P_����Ԙb�\�5O�OP�(��3��9�f�E�	c�֟{�	T����QW�������f>o����jg9u�w�OIB��à�y2�j��������gB��c%:� ��e.���C^sJ{�@�Fѷ=&��S�QIi���T��]�W���x��#�����T�lc�|�`n6K�m�~->3����4�8�٦�h|����p.0�%{j�l��!N8�e���9���uu�X7�*05t^��6:d����;��V����4����K�x8�*�P��8h����f�4���#nW�	&�ݦ��aҬ��p�=ds�PA��\���`s��@+�锠O�u����g���AVO�#��#�0��a1\x{��w�'"O��a����kD�d%�>��|��f��7_L��WLq2��^��ּ-���1���"��'8>��Lx=��[�� U��wcE<m1�|�I�?�M��c�G���Ňw�z�?]N��m��O=F
	>����@r}a��5���׏Eˉ����>�$�3��Jt����~�=��&��:$`甍�,��U43��ǋi���>=�_M��d�V �S�l�/8�x��oI��s�/8x*,s\�;P/���^Ѝ�$���ܴBȡ�w������4�n�V
<9�c��;|��zV�d�;Q3���V��z�B�&
r9�s>�]F�D<e�i_�bˈ�E�/����<�22�}?�q��z�� "e�����mÞe����%���!���~Ϯ�2|Z���V�O�qoEE���wG֠:�)�P�Ĕf�\斐ˎ�a�BE �U=�_/p��F8p��D�p�M)�AJ�$�ǄՂ!�N�玲�2c2�i�<J�D��Z�Z� 9I/��$�
,G$l�����~0����i������YY`��G8���@�z��b�����O�8,\���p	Y#�A#p�1�
"F�|�H�˖��ǙFA�l �W3��3&#]t�\��r݄��%{��>�����^��(�-�	����>����ˠ~]"6/�Al�����q�ɍ�j{�{u�m�>6���WKl�{�����]�J���*��iiǱ�g�w&�¦G�s���G8� ��#���3�6��?G43Et�:�������1������ow��A�_1!���eD{L�sB�\��K��m�*��x����>�Yy�Z ��WP/�}���R+�\��L-Yw09_�������G�	2��� �R�`0���h���ͷ�.@Q��'x۬~zxr��7n��h�W��J_�J�#�%i�{x/��#�K����D}K2�OV����<z�	��a'��kN���v�S�6����ڣ�@����A�J��*�S����[�o7�?�#�DrD]�)����f�O��j��#�v�{�����[�������]6a9��{x�M��Ho�F[��Ae����Đߔ����<Z'�&�k�$�s(�����ʭ��+�՘i���`�x�\Ye�!� ل�2Or?E=p�	���f����
�j��z��3����<�4�6	A��sZ&�q�_�n(�>�5�.��d���4���˪H.��lo��#��Is���ڙ,��Tp�l��V��$0�=��D���P�%��H��)K�����Oh�d��A�#�z$u�N[�]��z�*E<�	{��Kؘ/�������a��Pd�5VcN$����a�o6w��p�W�d��f~p��$=����B2�(��۔ճ��Yê�[����*tq�Y���)1}�BLD:����\�#�PFR�!!��T�7��%m�q�nGع�)����&��Œ�/f��5�Wr^`�6z~��⟲-�ǧ&��D�s@��8�/<*$���k5�6�� pa`�訋�kp�|�I��SS��uw�bD^��Zk��W���n(��SC�{���,|���t�ZD����QF����r��?:�q�m��Z� #k����c��B�r����+�HDq�гR@�d�����nC���P�7{����w�RG��R��[�P~f�V�2�.��F��������DR�֦���i K5�^�Nib�	bI�(��H��k
}aBQ{Xs���@����~&у��k�q��5ag���(2TB)W�|#.ʸD������+�;U���Ew�̋�N��넅��՜F�C}

�m�mݻ�BQH�w�F�I����a�#W���SQד��@���D@B,���2*NE  =J�z�~Nڦ�2撅h^@8؋C������+�l(���xIť�=OZ'dSly���p��S�0��L�Bl���aWWD#��_� \���fg���Ϫ�d`�1'u�<���=�	u蝋�#��1� �d���6���kZ<��ݩ���}�� �"�:�~8��"���b�lw�y܊le�2���@��e��?��Z!���^)A�v�>�Z�����������Zt8����daC�4yĸ��f��ng�iU���i�`�$f%	�Rl�e�Ka�@�ѩ���!:L�ŭ���ؼ߃���D؊9�s�Q�-���6�N��!��u�-y�f��;\ Q�*�j��!Ȼ	�?�r�n�*�ˊ�B�������P�hϣp6�+8���TR����Z�U��c����������z�|m�)g�@ n0X�<-�0���x�U!!��4�(h�R�{��{�B�9X���=��'^�HQI�eQY����;ݘ�t9p�.LW&�1�&	�)/���<���	�5��]ǂo�z���z��͉�`�`2i��ݕ����~�sG�?�8��$�x� ��SF���z���Ez�B��_��{�v��O`X�,�r�XT� �kG=Do�"Z5�U���Z���q!��*ǫR���~��7t����Ui����D��3��a3�4(��*����76S4��L��q����o��$8L-�`�W�]Q-#��� I!��K�\"�@�#�lkKd����Xݾ0xQ�`8$R���mm�%G'?����O�g�+a���¢s`&�[�IK������f�cJ�=����&BP��V?N�֥:|����_h�v��(,ERt�Ny�q��D�d�<zS��S:t�N�Z٦~~�c=8�ӈ��[?Bg�	���f��#�Z#�h��u��6 ��ư��$�'�NsL �~�6�%���Ih7��K�SjMy+��Vr��v�4��4��%�C�R+V�@Y%.�����j|�'`��pj��XΗ?3Ǯ�@esp<��g�4����򀖰���V"�K*�0���ol;\+�]L]�z�.hf�?��JA�.v׵$�d�opQ��$�4�}�U�ٓ�6�`QJ�T�g\�cknǫj{����F���K��
��d2nVȯ{�*�LĶ�Ǹ�u8d��Rf��]`�����y"8���?���@���V9U֝,�`:���A�������W�|n׌�+9'u9#�G�&AG��sw���/�f7K�?�P�K$M��$e������b��쥺��9��������Ry��6v_sS��@l4�}����n\p2��/�x�&����fc�}"^�^��F��{I�b�X�����R":�@#���������A����>ۯ$0�Ek�1"�:�J<��tYe%&��M�����I�ڍE4=Ϟ�C(�J�y;O:�K��T����c��y��2fޕN���eb3]RT��N��m x�h[�ΰa5��c,�2�������#�.t�w8-��'��߿�M4K�bZ�*7�4:ݪ��.�ؖ��:�|	]��|0X�>���\c�f��I�b�1b��Ғ:s�����v���=]S�yh�3�hᘳ#�ma$J[��{�Q���v/Ð���ld�t���3�YƏs�s���0��yA�$��t�<R��uQye쐭���Iᣯe_]���mxN�͞y�~	_�&�x�X�`�9�6�!���i�.����"*S��v��K/]ʭ�gڻc\9_(+��J�|#L�:һ3�x6��.����M�Wc��3����D��2b����B�ڼ���s{q�롢��Y��|\�ܐX�h������7�fXԺ�%�|�训��ۄ�-TL�R'��.�SkV��R��	*A�d�Y
U���ŚX9�c�ڹb>�xׇ!�+�X� �?��1�4����5{5�(i�d5��,��i�Z�e����{����5"�;,'�J�6��?"ʆzY��)n
��z�p��6	��Fi�Y�^�4n���чp:V�(���4��S,]"��Qd�HL���������'�V�O������e�����Xr���:c[�Xh�?zA�/�1�����IZ�K��+Y�`t������e�x�˺��YMVrFQ�����܄�:�f_Ʋn�]���JP�x8�_Y8�I2��%�/r���9�a��G<�7U J*W�Ś�(N��ʡ�ڤ�b��uć���B�f���8R�����o�7-m5e�����|zfdv^.�*Nç�/N[d�5������
8�o��h�E~ �\��W����!qZ��B�P�%L@|�3�����=�s `��i��@�m4�^ݓ1<�y� �7ZxOl������'�>�+���`K��oڻj���OW9�c��'{�r�vpث�JV���A�''E&�Nu�$��cX�p��^��hoP*/bU���lф��;\������V�r���Ֆ��C\�>�\6�k|"~�����Z�ii=�Wq�i
���֬�fmV�l��\�r���[8���Ӣܒ��$�e,�n�)Ņ��%�q&�e�N�^܆˳N���n[�K�� \-3�G�mX�Z��[%g�L�_��; e+�����9w��R��;��I)�f���A��}����%I&�5jq	�is鏤 b��vK�.�
�H�H�6�u�MF��t��w�)���J�l��h\�vf~�W	��V�l��B��?I��}q���94�m��u�`3�פ�Yk}�w�ŗ�OV9�kb����S�a=j:Z�z�;�V3��9��U�}�zl_�� $(�҈Vqle�{�ԛ%�w��Q�>��(g�3�#]Pnj.���~�eGơ�](H ��6�7?qA�Bfj�k�dA�������0��C����5�ފ�s�X���Ct��\K �W�#��MW�)x�y���t&��'�g������u`�����]�Q�ַ����b�_CU�5�@�4�f-�%������f�0^�+N�7
.Gi�-8!�خ�%L��9��㌲϶o���A���ץ9
�/�cc�������!���,v�|Y�sА�w��]z�[4��@�\(g��3�Rʡ&3
K[ߏ�ws~����"��ǀ�N�=�������a��lr:t��O;͜�C~l�Y0cw�\���ܰ��xm@����WR<=7GExuB~d�!b���#����2����	�����#p�\��еK��	e؊�o_��E�g˅ː�^� �����i���0%T;�8�MZ�%=[��$�g,�^cM�`I�|��Y*=��z��e��g	��̽���c�I��94�����i�^�3��kf���x�]�t|
�[�40��T7d�mH�=x9Eo5�D=@xR��q�};��������\�\�<eIYs���p ѕ���)QFx�(�0	��#؏���	�G�ҋƤE�6z�MR_��t;�@a$�����X�-��3	t*�ؖ 7|�}0AZ�tcoDL�xv�	F���l$������!�ϩ�v��4(YH�c`�^���W��P�k�M�|���dd���ʒKc+H����%P.�}~����/.�Ƹ�r�0�{�fu�L���~��*���<��_�������3�固.ʭY�Ӧ��L)�+��7.��%�ݬ��6J�|����,P�K^�����';D�u0w�-��-���r��Es��w��:�W�z[G�;��G�,��k�LS6kwH"�a^㞔W6'":,�38���*���[��:���֣���b��Fq=�Zd%�ߦ"��1+��e~<��;a�t��8�me�-ۋÆ^H�cz�_�,gݘn�Ĩ��@�~���^�=�+^T�E�78�h��L�$��i�w��bFl�����w1���'�e�����{|p�K�[W(�W"�Q�wkJtJ���e�O����EgndQ9٠5��z�`=��������VǬ�Z�C���C�HZ+�W���\$S�Կ\`-8r��;r�<42���]e�ɻ |���"�5�)��8v8n�d��'>������oH��"�3�zF/�_B9���&��	o���\D���[�i�����G��̬�N(|m�-�zr n^�*7���ꓰK��<���]~��ft�K��@�0�a��%?g|M�<��T���l�#϶�$W����A�As� �}I�����^(1z��\��XY�a�r�w4tF�Z����_'�3��$ۗ�`�6���Jٜ:cL9*G 3��ҋ6 OJN��/^����*ˡ���h���r�EC(���/F�����ChAOE��߁��Agea���Ē������\bV�W����)X�ġp�y8��(k��f^�d̴�;��@��x�˃����!%�{R�r���c��Ba��z+
7�/�"�]�M8�I�?h�w�nt�'z# ]�X���U�}���.�愅��tdjX�p�!���3����Ӽ�/az/:��
T�_(&��4L���k=@^�4�>��?֣�?�p�ӌW#2��!`�!��zMQ�uW72���*u�y[9j�<k����qAy���h{�c��6$ߥ	��(��7͵��{Ec�V�4�uw^�n�8Fi����,ߩ�8��,��ƕ����눅��6�.�	왯EhsB���pvR��qme�ڈ`.Ij�T-�.�I
wr����r�$Ôʿߑy�0�4!�4�@#�-�NZĒIn���4Ҫ?
�O���o����y�n�8���4�l�_L {������g1�^KTw+h�f��eQ�7�R?���P䒪w%�m{�<�Vh*~�&�}H��j;���� $d��
?��9��ߡ�T�noR++M:u��u><�ZMWs�-��5��v����҈s�Q��a ��G5���A��&+8M�q+���^dN�Tږ���VąT��yG���l�p�e����ce�`ݠ}�qq�$����XwyT���!�z�-�h��?�-����	��H��T���Ijy)�:}�WƠf�u��5X#�0B��S�3*�;|����B0��_���~�dKu��}�R�?���<���2ś8��q�/�ۻ#T]��;��l�1p$�~U�&��٥e��(�:ai�'�2�Hg����]gihV����������o�����?R֧�捈!����[��:]4<,��cԱ�t��@8��t�x��C�����6���ȉ,�o�c�y��j�����٫�u~���������zid�<a����H�/˫��?�Uᤫ�e���%�kd|��N��k?��Ɏ��{rX����1�T�D�V�ғ�ѯ$���i�%�J��=6;���p��H�-��ȬE�AgM�j;đx#�N�+{�v^7���9�	ٵسN}3�J�Of��X���Jפ�u��L��ɦP4�Sz�w��70�r�	'3T�rV�/O����( א8V�����%m)�]wd.��e`��fw�
3�����1��<�`�����x�ݹwX=/�`���Q*/Y��G*q�@TY��Y��o/_����`<Q���4�,���٨@,t}a�C*q҅��D�� e<�bڞZ��s�����ޭ�DQ�q�{���ܵr�\jW:-]�rT�`)���ȡSzα�H)����8L��钙� o�d+�|b���*䥦-�n���:�(hr	���U'>��Ư��D%�M��,4�irUt�M�0
��#�erq���y.>�$"�H>�#�*N݉�cA�2��1^P��iI��@��\��"Y�x��f��I\�/s�=�20�;���g�n:�K�S�$�������	�΁�b�$2�O/�䜍?{��CG'ީm��O�F%\�C�R�^��TA���TNGq@~P�q��l��f�&_�P��X=ly�~���bEb�XBd�B�m���&�V�g��x���e4�ܙ^������T�S �[uТ5~]���K�&8�͡o�|�ƾ���&��@�ḇ�g4]�	�?$��8�ɩ�4��`?SEZr�Kg��:�3�i�w���� #Y"����5c�k�WC~�zC�Rȕt�W�q�pfU��Ǯ����8�r��FS���V����b���e���G�C��_G	�=Uv�Vi�������p/��n��"\��w���������gO��>�w�и�Y��&9��������H���#�+�w��p�eP&�Y��Z^>�����<F�Y�Sߩ����i��P?	�b�޹]"!@o�c��0�
����
Ox��m�+�$N؇+���dN��	���ʘbД�cEe�Pv���+ 5>�E5�O~I�L=�*�_`���"eޥ���_Ʊ�I���GR��P�'-s��in�z��qa$E���L�B����(�����E��y��P~��|��`aN�Y�&r�X���S��R$�MAO	(���Vu�nA�,^x����J�V{0�f��AZ р�|KPXLl���q�L-�>Y���w�?B�7��dI�_g�ƕ}6HBC��?�a�� v��x"�K�}iMqyA�����7�cMOm�#��nx��p�"-dv4&G���'�Y���D@�<k��Ĕv!`�5?V����1��C�8�v5���e���5�s%R�����ז�w��%k����c��$�
%�\G�f�ʽ��|b�~Vc�J����ƛm�kt�j���y����K���I��w��ev6�XZ[�����3��0�7|��f�+������j'�4F�Q���n����	�˞�ݛѻ�윫q#�首��R�(���3�߰Q%'�_���2�,pݲ�2�qX�����ʏ(1Ǣp����u!���Q/���;�o����ń�5��[L`�T���z�
�?a���[�oo��H�g̳���]�7 H���$��~�����v�Sc�^[�Q���Q�`��hR�`�$9���,T��$�*Q۫6�,0�N8so"�����(O���m����+�J
3�%9Y�O]�����(�^��E�jP��7Q:)��WK�W)>jm�^�Sz}��K��b֓R�Zw���{������-v�`��m=S����t��*O�"$��w�d}��'m����}�0��ʢbx0ȭ'w��ޙ�愘�4i�v�7�<�!� ����$���\s�lU�|F��'���^������O_�H���]o��K@ 7'A&�;y#i<����@wڢ1\�#`�6GO��㉖p��/�\�����B�Ƴ���n�~i�V�(]Bv���]��~�F�� Հ?L0བྷ��K@
)r�7�����nVqծ����<h�4�
�����F�ߞ=�����29��G�kO�;���n�+d#_�(0�Mw�Uh���(sR�%����� ��3to�,	 �2i �������sԨ`�`@�A��V��t�1�.?��[򱧬K������ي	�A���}Q���$JE��s���a�e}T0��A?p�g�ז��d U�p7tZ�*��a1]	,�[�a-V���<� �`rG��E#I�����9pj��oޗ�?��{�H{�.E�f��/.�;#�X�2r9H�T�Z��E���p�����$]fy���{�éx���|WI���rk�ݭ�_1u���w8��Q/'[S�׫�:3��ߤ�]����3m�-���k��S�ݗ_��7��!fWs,�>�\h��^��Q�O��F��I���U����,@�r����&)��z_��L^��f��T[�+& �y/;Nl����� �ㇼ�q�z�`�(�"���dG����P�[%�H�X����C��Y����32�Z<���C�	��0G�[j`��@M/��ܺ-�7w7���SSZ[���D�Rd�ALM��qs#�� l���E��ȭ.���%�����������]�`���62��G"�������O~6�)�ݣ�rY䎕y�g�#�2 �
����(1�(�4*�i}4���M�<����i+�fؓ�]��:���\�.G�M�(9-)�ϣ���y(1�_�t���b0iL��/ˋ�%�ZLmm"�.�{�>	P�����y��V��OS�:W^b[M�ة�Y���@ f�`}���%Zt�;-����V9�7���Ue���X��v�꺃�T�1�T�hK�p�M+B?��>�ofQ�\b��YiQw�0����K7̢�"�o�F3Mm-����J����c�seW�̙�n�'j���#t�3��?�qݪ�<���b���; �!չD���K�J�
�್�"t���E��qz�t��1�CpY���\4,���*�.�;ձ��E63��5:`={���u��:��#��;����[�B�����۝h�x�3�sE
�h�o�;�m�؎��c��Z�g��L�F#L�S��-�I� N�NN�g+ju�C�����4�Tbq�+��ʨ�Kb��_�5Ֆ������f�7/R��I즓j�r���xiEV 9�r�Ɉ�W�O2�pu�S<�:�3����/?;�-K&s��P��J*C�S�z�8�]km�*5p#Ih����8�������걏�`Z�Y��ɤ:�\�e�Q���E�<�L�ɐr���A�6�6�n ��S�æ-�s�l���-A��`෭X�-o1�D}a

�ZN,�B@����t��AD=ڔA�7z?i�u,v��}vA�~����V��Ec4-ě`H��ҝ���_^�Hچ���P�(���
�F�^7f��
�3Y�ڲy��eU�
��g�Pp�BX���3HZ�yA���0F��@��"�U��؀�^��C(" ����i!�n2��O
��u��Z4����yN���ԣ!/G������$�9�{������<��Vy"J
n���G  �gْ���N���"	1�}�#P�)������i�
m���j����v:l[h�=y*|�j�?�J,C"&�11�{����^��k��(ԭp�"�d��*�S��T���mf�+cB߸9��a�Ps�9ˤm�� �q�UK��o��yֈyd�<\f�+��*5ӭ�r�_nVE(p�s�4�7X��	��������]��ef�� yr�����pu�}!)[%nFlM���
��4X��Q<�����]Z-ێd���R���WGnü��~ ��1?��~�wD{�6�� ]�5=�S)H+��$�B��q����~�0�N5̨������D���߫��[��'nn4ϡ�^��#���	QA�"W��9n���R�\�\�=%z.eU�2�����0�^[�ޖj6����N_hP���.1c�1Uēfu�&���R���^r����g@Lk�a�H�3�V��Q���Np���QWLk����4�y"������J�cs�\�+�6Մ}��QM~���пxÏ�2�Ʃ���M*J䍗�]�o��վ�sj��qAyj����Q��C���ұ�PP�3b�K�j�Ļ���⍢�0#7��!���.�i��{^�Fh��Qqy� <�%�n7��|,��Ʀ��=����4�I�k@��k�Tx�H�ρ��؆e��*��F���?���$��	t�h<1P�mH��-�2+:��� Ĩ��=Z+��2�!�ȹ�s$�|2I3]��=�jME�M6\�7E��:��D���t�LN��]�H{b���V�U������*Y�+�`+tE�+zz`c�MP< `+�@�a�"g�I��+[r7�D��9ҙ�q0�J���pda�̂�S�طy#�1/�r�u�A��`eT���)2+��Q���W=cqP'�YKi�*&04��y�"q�K `��
�	+$��r�H���-���!��➏�턋ؼ�dxDt�t���2��d���1<s_�O����5�,S�D_�O�����c��l�V���W�s�dV�T9S�/��P��ӨW	U[D�磞��0���g��;-o���^Q z��X�f6tʻ\\�˨ _[ԥ� �ڋ2&;�:��4f�Q����<+�=�oK\���h-�[@S�$����b�yA6J�ƿ[Z�%P����.;�Q^I<:��{ʅ�UJ��B��^�^�bYz�2��'$�
����I�Q�p���4��CG�(qT��A�c;h��k,cG�+H�f��M ̲�h�M���Pu�]�0��L�m\}诎�dEO�T��NsU'�,�k~%�,_p�����&7��1��{�r�fҧ�?����T��*�x���*#�Y��1V?���'O��ւ����sF�^^l��?1��� ��|��徭Vwq�ey��{�L����K�1M��uQK���ϡC����8�7%K�>"�?�(��>�<�Tȏ�fw+��E=`-�)���g�TM��7@�˾ڜڽ���3����!����4U��BO����mR���Y�_FG߀%x������7c��М4�KC�ĕEuGv�M�2�Z��r|,�c�NB!΢<�Ð-T��z�	C��A�j�.X|E
D]b{��&o]Vj6�ꚦU�muW�/�We�;a�9I�{��f����&�P���S{}F%"��"�
36+{�θl�%js/�OF�m!��N�,kXQX3�ʷԕ�&Դ�`���Q���V@��k)Q�ذB��_�7���"�[��=K���!e�>����"��Bg��c��&�����uw�d��Mm�{�@3���g(2 ��IäVn�+6�5�n�d��e[x%G�����Q�c�*L��CP��j�s^�ý\Ɛ쏣.L����{�E�\�C!	|� V�a
ң8�@��K�ߛ��x1���	d_V�&��J���P��dZD�;�׉���1��{�S%C���C�1��M/���N5�(�nW�ޟJ
<�{�%,��
qG
3�����7"D���I�͑ߦA���s�-����4:Z�Rvd;�{���j'���4���<�A9��1ל��"�v<��P�Nx��� S��S#bm{��
݀�ϡ͵S�
,�P���)�sMř9h�̯Z���BFg�8E�� v�&��LY�rr���<���پ�o�9hk�N����ۛ4,����|԰6�wr���x��μ��pXkq���Q����k����L�&�gT��A�����U]���M�2�%'��I ���c����6�K�3����.��gt���;Z_�+q<������O���e�㛎,��z��rj�!2��C��/��@�E��P� 7ZU=�"�D��+�G@+q�`��Ƚv3j���r63e���}IPU��n7la`��@KRw�W�Kץ�iT����������q��_>�+�@#0�r�%r}2�����
��T4�v��=��ˠ�_�e �� � ���Y��)@�/�.]��O{�=R_kᖀ=��G���gͩ7z>������]r6��������	q�i��y�9�:VϽz0�`eą�"��B&%�A,,x�a���?�|�^�y v�lA�H�s��r��W��G�C",��K4�f��t&Me����nQzݱ�f=�n<�Z���1.qxi�fz�)�{�ӹ�V����P�֮�S�(�*�&��*��.#z�x`} �wG���q^������~W^���twE��g��-���`��r̸���d���?'B�����N�����
��T��į��?F6���'�h�k��E���{��l�Qǖ���E��s�O�n&��� ����E	S��zn�f7���2�d���	��m'�Q
����qJ1��.��!��js�-8\�g��rB퍍l�P�����6;6hW�{�f,�яk:�U�|�:�L�����BD� ��+���:ұ�W)+����1�?F��B\]%��*�����gF)�a��7�VL�oNeݯ��@$�`88{U),8�S��,�`�+�=Fp�*��qϤ,*�SA��^<?�sA��
X'"�����ٛv�Ovi�Ͷc̮�v"��~4��m������lW��o���[1�~�����⼅�׭���1C�c�<��^�F��X���/�
��d��&����' �Xƚ� ɇ*2<�R��/�W��(@���Jy<�
��la(��S��c�D�ϥ4������z�z���+���_����
�L���Ug�̹��<��Vs�`��!6Q5��)�bz�)Ie��1w��X2���m����Ԗ$L�2�\E=q L�FA�[Cl�+/�Z3�]�J��.�x`sNl��DA�{�mմ���]����a��L�EN���c&3aƙ���d����x9����SR!d��b]�����˦���|�åԵ'S�h�m.>u�Hf��Ie���}��*g�$H0��1c��);/=\^���P�2�!&��l2�+gD��v�o)�I:[�7��Ѷ���)r�,yl��46V�R2ob�3���N9�f�������Z��{/G��26��4����E˙����3��ܶ�I��u��*Ը�J�r��`o�c�^[{ Bݷ����Wmi��Í����[�ܑ6��\2�&��}�(�d��X��.�Af~e�?��2]�K-*��U�X$8�d\�UB�)�Q`����>m�3M���|���;5�z�B3�j��� A�Fg���X:<rL��_4� ���B^�}��BO[N�lB�&y���s�P����E�$�v�?��+jmD:�:��&u�ح�f4R*$��+�Wj2�BTrzb\u��w�����^�r�W�;����섻1bZ�A+x�:�I�����Ml孶��y��g/]H�%K.MZ�G���A����ÅC3��زW�����w6�W��`Hv��[�=D�1�|�G�5�绮�EwG^�ê!6����g�'��]���%A�O�9N:��@d�zO��!�� �!����Kʫ�7�T��
�$���p���,�B}�D9(��@ƫ�O3��v�k`�{��" �:芜6l��S\�#v���9L��3�/���^	��#Y��ό�n���
ǒ!�S�#��S�Lkk��S���X٭N��ś�}�J�1F�)|��d0��0g�!�9�=M�l �s�xT�E�6��G�y�`�YTkn�!7���`�m�Fz+��fx���O��N�^��C���r���� U��O\D6�P� �Z˧���}�#HJ+Y5�ص���Z�^DÃ���Ҝ�������N'���2�3���,\�' *�ߩϳ��;�i��07O�d����kXv��[�x4�G�x�x䴸��z�B�e��;�>y��Y�{ET��m� ��#�#���PI�(�]��路��
#2�c­O	Vu��$��F��o��
�.	,+!;���W�x,��i��� ���G�DQ.���
���|��I-�j��"�
~��NV mZU�LD/�1s�'v����'ѕr��O٦vJ`�!�'$�����&���G<�گ
UEb1Q��p���P��7ju.��(�Bk�THׄ6D�U�j�L��v�<�6�p1Ewx���|��m,�@	����_G��7��S�i�[�å�7+	���:��J��!�Ӆ��}:�NP\o͞�Ck_t�SqB�@�"jv������z};o%�-�
E[��sXp�s�D���tJ�>Ɗ�s��Ay����/�ڃ�I5@��Y���\�a,K�\lxI~�잵��e�.�֦�Yp����3%Χ���=��ތmUTɦQ��*��)R=_�8�./s�P���4!h��nb�����u3�3k��؟�d��~�g�|��jH�sĐ)��Z������d�T��`�<�k���7�o��ϑ��7�`ͰG�X�����q����3��Qh�"u���,ť�+��U�"��i~�/���ٳ@�E$�l���2*�j�i�����N$���+�[c=�����,oH�����Z߰�Z�S1�7y�����X�ؾ
_�p3�qP��':�n �����#7���-Vk'O���NCE�4��2����'�xUu�,�J��8^7��in���Z����X��stO$*�XD=�=VE�Ek�#I�:��8lw%��Z��N�r��7�AC8%��w��2J��ق� d�5�~1�l��K�1�X'Ri��ېUeՒu\8ç[�5�D&�S(Q[���{G��h��H���~:LN|�IڅD[�	�jh_|�W�f�͒坙�D�d5�����<��C1;/��F�����Z'� �[`��!�58�Z�#�~����Ik����7'瞠�|2�A\�R�,����u)�����lB�İfJ�����U�ii2�
��������H�H}��8�Q'9�ɨ�@�=��B�0��d�JJ)κ�R�{�@e]/ztu�O��7��1�L�3�h2����}Ql��� �Q��z��ց�����0ԕ:l�΅"`֡ׯ��o�#�'�^��E���N��Z����Eg\�N��9�[�h�g^���� �����}]���P)Kq�-2��:�g�|w5M>N�S;�����p�9滟��/nKe`$r��-�ky,���������I?h�jH3�;���:5`���Q���0�wؾ��߬+,f9������I�'�}G��u-�0jT���K��6���
[/1Ml���3���y� 	~*�BZ_�.�! 	���m_V���X�4��E �PH�!N:�("2�'����G�Bŵ�+��^�� "9��G��SI׀����|�7�Q,m'<�y
�@QZ����#`�>w��~~�e
��|��[����O��)��q��m ��B���ml��Wf�8^�dj����>bM��f�M�$�X�n�~qn:k�m�?g�uu'��%���.VZ�dW#8b%+-J�byG
��Sl<���D&>����%�Zu�ς�=�A���l�u�4�0���ŘD' H��Z���0׫���$�I] ����
5��a����ų��!(`�/�߭�/���=�]�$Fc�G�g��jz?�Yn^+�yT86w�Z:՟�L���õ��(�c�;+�x�&u>I�?8Ph�ð��2w�3^鳔����q�e:9#`�ī��#��k��f Yb��ˉ�G^?\7;��lps:������uӿo�I�d�����_��ԩ�`kރVeR:w'�ýN�b��J�+~g/FpI6��"T�F@�~d��E�!���m�85�_��)@�/\]�����`�{H��z�T8J�֠מ�%�z�C�nyt��S��7����\����ZB��ޘ�b����S���|�FM"⨂�a�q]J
���*~�yW���)*���)��L��f`�k���g����+1P�4�=_>թଧ�w� jGI��["$�#ģ�~2������@݇��8i�#�s�[�U	&����iK��B*��pG���Lғ`E�<Nը��ƘyH^\��n>����esɕ)���wR(���Ep�n_�e�-q��;��.v
����tq2��O�,��7*bb �YF���=^�0w�@I�����-V�Ir�wT lht�)�R�yV�ʐ�v~~�c`�q�>��e�~2�1T��y���K��i���g<��^���f�?A����\��X�<9�W�1B�7����Y��>�ٽ�e�H��8��d޵�d$��7�`H�w(�\z�ϾT��W�P��}!_?,���� ��SϬ�E��ϔ h=Z-�D�Nq�U�2��V�'�F�Sg� �b%�=�8�P0;c�K�\ݐ^Y�L�/I^+ 2y{���R�!��f��}!ǃn*-Ը��i@��(0��0�IK�U�6) a:]*U#MwT���:^Z�ǽڠK+ֱ�vQ�,6�e���D�����o�� k���`ٟ�%l�S�4.N��h3�)�Ug/�Q�{�R�����f��i��Tl<��h�ғ��*\~H�^f���Q��Hy1W��7����
��@K�*�S55�o1���C^f��^�1� ��$P'ʸM�X�*���!��o��5^����vC8�G��\�L����{C�O��SM�J}��{Ю�{�c���QaM����FȪ	e	U�>Z�����aBq�o�\��H���3���+~Z�n�[q=�B�s#�W�p�KJ�)���#��ǸE,�ۀs�+�j�U߲�E!���5��2���M7Ҵ�'��A�G�i�"�|V!��[�\����IS�:�K��TtHj�0����ԥ"p��2{��R�k%�sY8_�!Ub�������}��.�-�	;=���	�ؽ�Aw1�Ka�S(��o���y>�_7|�(�Y��
�S����EA�@�`u!�C>���Ft�9���l΃���$:��Ԏ�>����$��C����-�~�-����X��\/�M��=ziʹj��-'W����y*�����̰�$�V�X�N�#7�:�S���ɛi{dt
���u+�	xB�5�,4?���Z���xDdc�����v��k�(Fh�;��L1 R,�1L}�*r�Mų-]�.�4^87��S_�����f�~�%���\GR2B*��� &�k��rh���{�*��GI*�e�����ѩuPQ^���/�aO�Pۥ���u�ar�8��]�#��#� �M]��H���Q�/CmEY��t�1חV߾�(�<� 1�{;�y����,�0+�����f�!)���Qk܊����e@iۋ�EQ�%�`f<~
shv�(6⠍��$p�X{�7�Lg��y��/ؘ�h�E�|�2��_��������k2� {�`�Y�9NJ�b%ϡ�]_���:Z�֓Gjl�n���])PR[o����J�%�U;u��� o��k�Au���>g���7��ù����9@�7����4.�[��5H��#;�yeqex&�����+4��Lp��m��@�*ά�Z���>��]�*k����ޱ�sV������Y�L^"j�Q�0с������b�3�<PrH&�-�0,���?��w��x7I#UPӓ�Uf����L� ���>�f	��^o%�G*��;�]_q�hJtD�qY$�saE'��:Yc.�ucD�*E����I�qQ�dN���l�� W�<� �vL]�4Z(/���'`��!�\]�b�n��9ʾ�'���� (eN���H���P�k��_�^��-RX����Q�����e�ooO2��.�[%�4�"`Q��׋u;DG� 8lo�����9u؁��k_!q��x�^vi�\�Y8Al$O8YQ�Vv̘�1˃o�mb'{1`�i�6Iy��4['��e���ރے�#�D �����g�3�f�K��3�1D�>��1R��g3�0� :��E�=��,	)a���Z6�{q-�9�I�+���A-�bz��V�ۛ�)ğ-'{/4����v��.����'%�Fp�Y���~t$S;�:l�4.�O�鵧u8�����?�[�v����aY��-�5��J�G2���gsG=��V c��c�D�b:�n�o��ix��SU1sh	�.}Y���
�[�
JT��.x�<��-yg�p�?�d]D�Q���6��0
K�S5��;�I��5=J2@�|�W�a6ؚ��8&�\�g�mpt; Q���LP�����d��8�-|�S�e��5&"��P������b������smsU|�����I�)$���!�';C�^;H�6�CV���B�e�5x��1v��a�Y�?�w[O.�9	#r�h��NmN�bi�'�-P�<�]yE�W��X�g�B��?v���1�6��u�X�z�XL֖���� �[
PE� ���C�T��
�d9�4�!����艼:���\o&�c��/�{�|	�V
��Km��,q
'�F`-�[U?Ns/}jg��D��-;�Ϩ>N�����*��F9X׬Ո��5���3��b�-�ga���&��SĦ#�t�D樛�:O)bb/���R6�,��)%�܃����2�Xm'�����V5�.P������_���8e�]3Z�r����0�́�_��$é�aە0
���\;{�!h��v#I����[<���d,jo�rU���Y�����{��'���׍{��������>u<�A�BZ8k5w�C��j�e�.)��W�w�,���  ��Zxl�vz<�<��i||յ�GE�;�?���[�»��+ͺ��9݀��#>^T������Y(�wix�qǗ%^[C�LsD��]��;�[k�,D�M��mG�~	���Å�q*A�H6Oݳ6t���p�4��a�z|�g�S~G,���XD��J�:�ŏ��(�Uk��ݽ{e,��Ao��SO�)��|�!�h���!��{�4�~nҬ�D��7K�4�Ma� �eQ͈RE�{uT(S�?71}� S���_���:�T�򸥍�!��\�����.���a/���Ӯ��W�_^��2�R+mÖ/C���PFD�|�os��s'�u;l��5����FE
%dx����<}@��[����!}�� |��te䎣#��@c�M%=z!��X����[���j���n6Whspg�s�2�&U�u���α�x�t&W4�9a4�K�:���SIs����K#,��p`HH����j�@H���-�F��Ik����A=������j��N�[����R����k�}�.��'#t�X��7D���:2I��
���D��j蚍��{k�Z��=��b��)�뀃c��#I7���F�] �8s����6����2�9�!'���u7�4�4���N�X�����O9dC��2n)���F��������YCmM���;59XSS,��W�~��
9��������Ϧ�>����4Zg�X��©�X��5/>o��(���)_�����@e��`��ddp��`x`͐�e�3K���҇y{��^������A��W�SiM��F1��`*��
���sⱏ1(�� ��τ~J�o�I�j�41�Ŭ� (:�*	8C�����L�p>�s�R!��y�A- 	oB�.	z{�iSi	F�k̖#���LA�hBQф�dx<�VSE)t-fz(�j��&���0.B|݂�K��
�/�ZO4
�Q1g�/V�F;�AS��݈��o��m��Ҋl)L`��%�{9����oE{��/:��C�8�����2��y}���r��|^fS#ؠ�~e��`�����:�[�`���o �Z��5y��(�M����-5�������!�^�x0M��0����ɨ֦�݂E�]��N�1����)�ż��[ȫl�6�s�("�`o�� ��Jď�G� *S'�K�ej��e��N��������l��Н���{��H��ud����cTXR�ra�N���1�;�k6��]�HKNfb�=}:2H#A��ب��o��M��h���4�Rf_A��d|%\�������p��k����^�8VM��r|�U
$eNR2gS�\��o�z��&�$i��6����p`�������oO�C*sӜ����+r(�Q�2���uݱZ�.��z������ >[9�=\1ZEb?Ք��D�g(��L�e"�bh�D�8�<�c�X���TXp��� 692J��ZuQ���~rC�5i��X����c�H3�W��؞���"}��;'`���[-��߮y:�W�"�2��B���w.7Zد��By�n�
��I0�Y�X 1�9p�Y����d��1�C(�2�&Q���ҚއQ��~YE2�#,�[c\yɨ��R2���W"�.����6�15X�WM��Ճ6�^@7���"Gޣ~��u���2�q���_�u)S�/��k 	�&���"D^��=��,A#zR���L��jPS�f�E�W�Q{�?�r����DRC��u�@�,�r�,\�����)\6PNB�~���-3��c�[�C��h���B�s�~��z�V���4!8��Z���ڲ'���wٴ���T�[�į�D뤱O.��P����Y0�y5��;�M�t¸?�_�
�q-��CнP9�A!0�����r��_���I:z���"�Z��˿D�R7z��~$?�o�ٌ�3H2�W�iF�n���
%!�ܡ����o�n���[Y&�r�\��up،-�y����"�y<`�9ߊ4��ԏ�E�~joVu�[K��+F�_Z��F�K��%��|;�̜�y���N��PHm(/m��V7�q*l�i���Q�F#�%��h'�G�R��o_LE�Ȃbe��X��pMmaTȝ�z��2SΛ�?��Y�mB�UPr�b�X�o1F�{碢��zxI�̑���c&pT׏4F�*�4�r���m�o�J2�`��� ��2k&�³��
E���NMM/"?lH�ZE���Z�-3G�����ꇟ�puxj�7�ϧ����5TM�D�<�������6v���f��e�]����p;I���&���9��;��|1R4l��>�"D� sdl8��)�H]2�|S5��*a'�|��>ϓ�	$֔�Q�v������9S�g����$����+���,�>� =����.��D<v2^i�S(q��Eϓ��<hv���>6m�&�դt�*p�E���O�+c[&��ǜ������Nx�D{c�	 �T&�.~���V$#<��2#����qq6��{&uiR�Ũoll\�b��'��z��N�n�A�E���O�8أmI<��z/�"�V�����ݓ�,�(��|�����O�����9��7���ܲ���lGGo����J&�b%�m'���%W�µ�p�T�w��F�'AR���wb�7�'�i�Ў,�¢!
'��+��Lf�EÏb�:8k2Pao��J���U�͜)�u��(�󈴨#PvLJ��)y� ��2[�'�y���ҍ��-�x�5$.�v~�΋@��vG�Gc˰�l�ӡ�WV[s~P��T�xl�9��2�D�?��ҡ��ל�r��p`����[��u�7��)���L�ux�X���\�<�{*|�!a�B�j)�p����o�ɺme����*	�5��_�]����yU9¶�u��/�)� �to�W}��|��6���Z3	�s��w�9w��d��Hwb�QO����'�µ$6&���OصS`b���D(d��
�xۋZ���C(��G٠/Y3�t�c�ē&*gY��� ���M�*Գ�.�{@��h=8�B����?R��Y�ܯw�:H3g���B}+���T�bZY�/��S!E�������Q�:0v� H��"=e�)(�Y�f��ס��s�8F�KģQ���qO���mW�q:�^��e\��s�wݲ���%�x��
�#��^�;���))I��Bz�����s�|�8,5����AɅU/��%6q,B�(����b)��&�z! $o��9��(����3�p��(�bKk�&]ն,�zb! BH�:�ո��!��Wz�I#�v���|�f���c��+�0ؠAopoB8μP҆�ﲔ�/�f�o����}����g&i��P����|��v2�͓Mϟl���`�ܾ� �!^L�8(#��#԰n4���ֲ��6��ˤ���vW�:�V�pHN�b��N\�������wu�#s��౤��8`�`�ן�-�C� �g)h6I-�˓�,���	���+Rʮ��v�
�
����>9M�Z���?�I���^Cj��0':
���<2 m��Z�>g�2�m��Cu�U��X��0�$�|��� �������c6-��I���A��z]o��/}��҆ӫ��8G�;M�C]1i� ]�����x&.�������Ʊ����7�D�)�U垠�ܘ�cIb�E/��4kÜ-g�î��4	{f(<�Kqʎ)��&�2��?!�操�*��PK���!�nr8˔�Nlܫ �$�ɤ�M�ԣ�\x��_�q`ɉ�;�$G*�H�e���:�1H��]���n�f�l���*�/��P*I���S1�T��(4�����/���zi�;s~M4��3�:�_��N*����]�w��֘Ёt��s^,�1�Ssi�F�a���%��#W�fڭ�*t�[P�<�܌��6#�POk��xA�}���A�t�B���Z�šQ�%?��9����^f_��Hݡ���v����]B��2�PTIН���v�x&p_�Ω�l��[��,�-��d��EhƗ�Pë\�?�e����=���,5#y^�`tJ��M*��Hm+�V]�����\�n�;it�)?
�Zz?'���?�n�<�����5L"�x�~;���2ז���WJ�Y�1S��7��	�~�ֆ����8�B����C��Du��& �X��/�Lv�d�|���Q���91״1ܫw-���6��{��.���z�r�9�  [ �y^GGA��G'�GM<�X+?�)�~&79�
[���̒�Ǩ�W�.�>�ţ�Խ�㓒�:��}��"ڡ�)���&8�i�Uj;tO5D�E!/�O�a�iPT1#�)>$���
{y��a쀼���⁝�)9hV�o`dh�\�!�o�N����i�F���_�d"��S�\��Aq����g�ׄ
@�x�p�l�d(�E�bo+��+����x�N�
��ZX��\U^�R��Z�1��^�;��VVa�r� X7^d����
�r}���N��j�>S�f����J}TI�҅�f�qq-Y5j2���$�P��b���ܓ=`�wL�:���k^�t�"g�B�;%�# �+�m_,���_��S��6��<��~�w��d�	�P��U�a�4��h.�VQ���7b�v����� ��s���׈�v	�c�PY��eO"ؘ4Z��^�;� ��C;+��@j�nJ��VS?/��ͮP�{OoZbI�	��%%�P�vWt$~�}���{���[��[bE"az-H�C���=�<�������18�q:�D.��5N�$��i��AWH��5ϴ�?�|�.s�MN+��U�yɰf�,��<�c�����G㰹���2�nP0C��S�wu:�<�_���J�ef���7d(�I��[���f�s�N����\o�/p��`-g|�����REO��#"�FC�8���Nd����I�G��C#m'TW��-���&f�`�DiիP�C���1m��ˆ��-w�*.�.�A����]7w��)��~����&Y��*`��{8�\d���)��z�tiݜ�?��|��3O0qm�r��;��Ԇ琅�;�x)rח�GhX�n�](��������,P ��E7�#�f5΅�u4�c�x�G�4� 7T������N58H$a��/��5Ⱥw��%	aLk:�<�����@�	\��v-�8ߛ�9�7�b���~Ո������.Lg�}����^��v�����x,���8�	f�_��|)�����1d��[����|čߥ[����z����c�V���i�ƹ���~�h��.c�����z2��C�<��m��;�Y$V=R��/#r�2��ɊR*��wr���a�ѹyp�{_t
�8B��3���ݮ=i���ȝ}p䈠<~w|�h���,��[`�� ��o���;�]MXsFG�fm��$EMF�%��I�9��dG��n]����59��������Y��k8'5
����� َ��QD��)vwZw�g�5������'1�yIa\�}���N<�
5[�x"�I�6��i'Q�;,6svc^ZM�hMx���	H0P'K�TM��";x&�Vu9�NY�(S�1̩��s����&��ȽUz+��|Y��hV����u3������:���p.t�)� �� ���}�)�nJ0�h�%�t�NA��Y�`��\����Ⱥ8���H�����]�#x�����m��z<AP�_���n��<�����%��+>R�Kn�z�����VR
��˰uG*nc�MTw�_�Cx*�jh�z��~��)�K����-�~N��X�7{^��Jh��_k�1�߷b��5�e�G�5�vw��*>����V�Q�")B�C4�<���u�tq�{���4�bh�bk�w�4$lޑ�B'�)5�O��I�E
b ���5��5*���11r�%H���z�i������Whq=�D��F����p�sVCB�a6�����7⨕�����8+4sC������i.
�,<�+��3�����o���.�����L#׷�*��|x7���X�f�
��=��������8�[8h�IDu�υ)���0P+�*^'F�8Ƣ��7$������7�@}K�MU����q}ĺ,x{4�2��뤆U���r�2�vcS
�����c�r�{��$y42k�٣��idn�$kA�1I3n�Ib~���O�������̜{.��ek�}M��u{��)�j<�=��J-�[=08��
���].��nh73����:�yc���Q�~�l�2AV �c�N5���.mo��5�����LO�Q�?fC�Ar�1ȋ���n�[�Ų�#/E`ā�_�'�<��t�>~#Qf���r�}��L]���x;�l���=^b�E���`������=�nG"��48~q`�D�X�cQ	{mK.���v��C]����
��|���\� VQ13=l���q^���o�--�̜�IM�ѳ
j��$X��q�+_�C���eR�1A�+�y��/�&n��|�x-T𡻰s�[�騞�Ъ�����3�˝�maT��y��\ܸN��Z�6�(W�B��il�~2�W�l�Ho�c�D�R( �$�3�y�S�
*6$�������zA�[���j6�ϴ��R��Ò��ū��d�$˝X���x�����&���p�~��	%�u���]���5�^RA}9�/��낙׼!O�Ёe?�Wʎ�1�N��]�&9<*'/]�;`��(��9l�Օ%O��*��J ^�5~h�?-=68�ܧ�!�V,y���İ�����Vhi��M1J�N�$["{���LU톝\�@x6���0��(-���-���V4�M�M��Ȼ�"�N�n<\��|�Z ���}���}���SVj$����%��L�^� � �̲�%�����[:е�'6�E�j�iS0�
�
��u� mj��)PW���=��t�4=Jjj��{kg�1���X��u��+z67PKq�7Y�%>��
v�e@P��W��V?�_	ۯ�q`8`q~��`(<t��2>z�.�~�N�0@� i5J��VjtY9�We����g�昿[���d���HK�=�dr���bb�G��<�.�K.��b��܊�K��$��4���  G߃�1&�*o�/u�� Z�׀�TV�v���j�_p�4��զ�������TtRO5h��@�zZ�;ʄ�Wi钽ҝ�HsW�ʹ4�&Cʈ⠎Ѹ��р���R ���q?�,$)�;�\�i�yT�Y�4����`_�;U���H|%CS#�?�O+�<2hxx��B>^���Q) �X��7]౒��z檣����\��U��sq�hġ
�p��+h^ #؂��
s�L�
�^�����D�;��Ʀ�[��M��U{��NU�#��`��� �!�����Z��2p�|�p;W�y��.V��܀)xu9�bT���i,�Guȗh6�<M���Ԅ7Y�"'U�������Ҟ���l�Q!ʚ��}�����]�;��p�h�&x;�=�ִ<�4���:��N_��w��O�x�����^��X�=���~��q�f|���A�X�< mh�� [2�^�4���6�j�B����s��]߭x��a�,���m ����:	�U>��p� ��B�T�����{�ݹ���S'Kehn8�}zyB�c%�%��4&K�Ԟ�=���KS�oF��]�{��Qg���v��?Z:D��/d��꾗uw�<���]�Sz.�ꪸ:=��F�8��#�`Sm�W(?�2��G�$2�ht�L@��d�c&�^�ѩ�eZ�#��uT|@�xo	n�1�K$n%����޼i��X������W �W`�r��Yً�F��]�)M�{�{[I���=�).��_�}蘧��5�e��&g0�X�x�w���M�n"���+����Ahay���w�������j}�r���# e��;]�xk��߉�����k��Sz�_�����g�Q�e8������X���"���MV��>)CYI7��3�p�cH�
7��_���/G�\��Eĳo�G)�����R����rJ	��&�z�q��8��rÇ�U��g��AB\.n��t�O1dI1-�)�2HLO7��vYC��ǩB�_T�O��R߅�_� �筊~��
%��X&��m"]������n�_���#6�^� �}s�8��aE��
1Pj�y�gp�{Nh�S�R��z哚:gK��8��H���u���1N���������e�,+܏���w���hD����*�\Y����Y?��_�/qa/��nq�tr���	�`��fv������D8Y��\v�1!q���QDZ�Y:��WL����6%Y���A]h]/�}��(��������&)SQ���������` eE�T�?��bW�K��Y@������Ң�@Ѐ�>���2�Q�MRyCxSV�)�g;28��jL��)��}i(��ðסA�~��XeGa�v)mB8�9�?�ѭ�s�J�����������@��s@돵[��g�IQ�6|�3���cz�zب.[��Y�h��[d�l)R�ޫ<��`<��Xw�n�C�HW�9�Daڻ�T�ɍ���SC2�D_}^���k�pf�J)��$ �%آa�ҋ�L��dQY.
����>j�֜ʡ���U��f�z�����9��N���k�Hc�>4M�ݺ��k�쀎�zh��'�!�`�-��r�~�z����*4\biJ�$b2<�;�+��O�/"���(!Y�7��'墏:O��{7�^|���f�Ԅ�z&�x׻�j�%��!F8��aõ(Fx�^�kb��E��"�F�=������V�-�[� 6���޶$k���X%�|��^ �j��L�4�
��<4���$������V���q��(��4LW�K������-��Z�GɆ�8ӳ�Z[��V�ާ{�e�hjR�u~:(��7d/�i5`R�,�3�M��D?
��z�mI��N���:���߹dn�iK'y��G)PzY�EGn@�>Hh�מ x�A���yEVW<�����+�1.jЩ��t��B⊮��K��C��l�7#� �?� 9�
F�?�Ɇ=�<PxeB�Cm�?�
J�F-��jBH�9'`���O�]���l�o�ZW��z �������;l�Fp�欅^�1�3W�<V��[O�m��P��L��y$���[Gݲ~PO/��J���ת�"7�S|$O�Ft3���c�^9��9g��'���{K>���E�S�|<�J�>	�⊗����~ �6�8�����d��>�<�%}��^Y��� jt[��ޠ �(�������*�z�e���Ѣ������c���n�2b�!SIH�6�MO����9o^P:�S�p�e�P}�
����{��m/�@����D�N�2j9դ��0&�`߇�ssT�ս�"���V��Uؼ��|
	TW({���ʂ;�&�M���t����\l>Q�|����f�M�O'�zvE�	ֹ�&`�s�B�>r�W����`���0r�l�������	lc�sWl�R2�͚� �9��i���D�v�l�\��E� �Y��&�[��m��@]r����6��Ɠ��G��M����fu �M��ɖ��7z���	؏�P$��� �kܽx,�dw�/MԖ-����?Z�F�қ�/�Z��p�Z����Ǹ��PJ[�+���}u�p7[_H��uY����=�	�@�*��[�W�ϩ2�u��
O�R�T}wy��QQ�!/E|y�+~��y$��ЍR<͛�"�)� ��;��\�a�Q�=��X�TxO�ϫ%IJ�蚁��� ˯�=��R�lz�B��I�A���xi��%I?��pc��B������ 9lu
U�lKh���"4Ҩ��p�dLN`#f�R�P��&$Q��iɁW�B6ռCL�|�ۿ!��`<`�GK�Y��JV�%TG��tT�:�q7�]$)C���ڝFs���_ U�h�L�.@�w��QW;�V�S����͠@�ݟ^(�tS���i��������ub�����Qe�<�ݧW~����@D"C2o���<��$b�2�'c�I=6��*$��#��ͦI���$� ��^_Qs1Ȃ�7�HJe�r���L_!�i,���z�hv���{X��:���JD�G����+��<�	̣�ױS���Ƿ"l�P{\@A-��kl�w��-x��t�i�Eit\���>���IޗǇтy��!��Hq�*�g�
�1Rn�y���X�m�>H�'=�Ը	j�$-��-��
?ɒw�$���rݩX��=X��#5�$�:��� ��,�ZHT�#�����XM�LIT��nP�BB%�|ږ���5��{�nla��asp�WŔxטP����km�G��ۦ��J�ji��]&I�x)@[������"ۣ7�^��T�5Ed���l��^����/���>:Tp���E�L�J�7�Qծ  �2'M�5 P�#��|[�?��u�\��fԞ��<���{ڸ�((s���p��F- cɑB�����:2z��쨷�����9;�F ��G�,��{��_"��zHh�\)s�Q@V���?�'uJ*��#�芬{)��N����7����\���S�) +*��s�I�6�Ǖ���vq�hMAK���3f՚�Kݻ]Tn"��!�_�G*P:�z�-2VK�_�;�� �9tH�1�Ǟ}R��Zbg���,��-� Y�p��Ϸ����u�M��� _ࢯY,����JRn��b���4 �T����CKC�������ż�P���b��t^N�V�h����о[�������wh�{[>���ۊ�#���H����^�mJ[�82�B�d�sK>�).t�V�֘T��̷�*�M�t�+����W֐��Pa��S2?�)�uRud�F�����$�6�~�j�;���J�4�Ѩ��/ ����;	ss�Hfkd1��]9�^�ʥ���ْ���W�{��0���^��`�S�/'�s+}�~2��OWl�i���֑��aϣJ_�^�����5j�c7��O�����v���:�0T޹�̭���£���v.�U��|��zw��[T��4�;��X�z�KS��z�ep5D����Ӏ�e}3Y%I4�r�!���(Mw�:�ӝ�z�W.7� ���E�G���#*PLƝ�@[��r�����V��Gx�S��@���7�bL`��<!\�`�ORbo�qNd0�x�Ÿ�M��i�un׷R�d��ja�d�����,G� K�B��ဉ���:=ѡ�u5���HN�Y�O+�E�Zԋ��҈"|/v=Wȹ�?�M��<t��]�]B>�F�����K��/]hr��=��"*�ٺ�T����&�� ��pc��J����{�@,��^��+�Wo�`״I��F��D��RpH�Y:���U���U�"�'I�����Y�71�����7G��u�I<�I/5$�ݟ3�h�H:2�Í9����6~V=kÑL�[9���;�����D9Ea״�I�&��w핲��UKD�dL�p?U�+p���*���jn#�ΕH!�Z�<��BQ� �'I�&������ʐ�>j�a�*�p��ȧ�w�Eb�c�^�j��W0@�-��oġ�a�;����eJ�},��H8}�oD����YKQ�����*9kD��C��]��0He�?��k>~[]j͡�y�g z���t���5&<��#���!��p��x2��f�NyAqc�� u
�tE��xz���ä 7��<G"��d"�w�'"�ϿV�����y�<`M�x5z��B�va{���V���Y����6���C��OZ�=3?�A�/��c���qNS�z	F���]����Zo���]BO���A޳C͏|Q��K��Ĝ�2,'�fq�E��(����B KQ�)�ƒ�<6�(�|��bT8"/w_A��M�?ַ��Z\�� e��m�Ί�E�W�CsٚY�s��҈���NPu�n*6�^=<z��*�f1�Y�hnx����T)�B��ð��R�h��h�@s�b�O}��B�?��=�6���rg�]~��"���y��s�Nvs�0- �����cz����T�����{�ՐA��p���9��}+��ޥlf>mf>`���žX�2����~OG��?��䝇������\%��:�i��DA"��<�ẁ)X�;��[c��Gz�l̶�ˁ� �k\ߠ�/�ͮ�f���� t>�6^�]�����v���������p�:�]��F
�^V��Q6{*��y�z�Mb{0�������k�`�?G��? ��CUkܹ�w��9�F�P���h�/�qS�(W�OmH�ue�����[��G�Y�|�h�ୣ��8«3Gd�1�yk��	%K��P�ٔyG��\�r�y��*K^=f�bX��݊=	-͌��ؙ��Q�s�lE�H�h��a�Aΐ}BVB��������'��\����};�h���n:���S�����Nw�O\ȋ���n�9�WF��N�f���􎀫��6�Nc�Ъ��L�C�!3�!Ӊg�yG^�^�E���JAa��m�0(�Tˊ6�\<�Jj} ��@�HF�cs��R4�!���BA����x��OP��E/��+�`�7zr��^&�k�B���QV۰_�ֺ�q��͞uUe���Aԣ�g���h�bSMl@͑k�;%�9��_ac�<�צF���YUk���	�������F�+���k�^�8��댾�d���p��4-fY�l��eӝc���ry�s���eQ��+Nб{ �b*���mC�K��XjW��r⎨s(����Z��CJ�w�7�{Y,V��-�+l��9�,�P?m�a|�x�7a�o\��(Y�x:�U	�L�(����έ� 1�g;���\�Gq'+F �d�+�*/#�?�i�qIW,�
��/�إ��ѕ�֬0N�C���X�y����]z=��A0�F�
�n�CXw� �`�¦�t�z���Uk�6���|lR[��e�PZ|�ދ�N������R��l��k�C�]�c���YX˘���rs�������5^uOVS�gQu`��ƨ�?�fRf�rx(��k�;XJ���I�]��:���O>����y�����z��@�E.��&��$��2�r�V�5��v��(�'�,G�$GCp-���۹u���ڔ�����&��Ml-%D��{6F��Ԥ�_��M_�SȾу`�cd���S������k�t�Í��TZ�4  ��JU�%C���>K�Yw@��he�S�y���ǍU�X���1�S��EA�ӀF�V�'�r,h�i��Ou �%̣�4QW0��wG2[��h��<����XՋ�l������Mt#�"GJ�xmB��
����|��aV�(G�/�Q�bf��p��h/�K�tj�~�2�`;5e���6^7	B *�J�������>�}�[B���i���j9*T�78����cE���0-k��;��QÌ���"�CV?���Z8��)WY�u��V���6^E�f7�q���0A�ۯ|�9�k�ڑE�|8��|�:�+�O{ڌ�$�*�������f7�sO.&Cٺ�ޚ��,����	�	[��r���}�]�#J������ؘ�����t��@��K"�j�z'�E�IK��䕽\���Q�h�H!���F�,�D�g-b\?:�����!��n��.��r+$�β�B5_*��KI�o��3��(?��30jڇ�2O��ɫ��Ϭ c���j�Xo��o��U[Y��-5��\�� �Ee)U���o�H�u�eZ�ɦ�L�*8Yn�;�	�-'�gO��pt��a7��Eu�e��e�/��|Rsg�w�q�a7 fCBY�yŕ��H?�&/�g�*ao��y�F�h`���*��7����S��T�%GU���	Aت�P��8"5-�t�q(V���k?��lX�F/%�kO5���P	�W؞>�^w�ɘ�$rPd���N��q�q�B�\\�ªi�`�ya9��-bA��z�cebJB�7���ѕj{&*��;~��)���5n%y�5}Cǻ�n��8�じ%����l��c���0�)�ąc���T��f	A�$�:�,��p���c�8�~BxW���CY���к�����z��;d��d���o�e{�T:��O�JV�u���d[��na��Fi�A�\z����*�K[����\j�'����l�f����9nQ_r�/���<qRDّ~�n��>�l��kSLeq  �Rd�CuSC�p>��ޘȫ����G@"][�}���tg VW �$�<�zҊ"��44�}����,qƆh5���V�����r(���������&�'�[�w��3{�q8�y6h]e����[��(�@�����J3���cV���٫>d�Y�F�T�D����5ڱK�~���s?�6K�F�2P����:�vb�益r��*�Ô��*����O�������F�9�o�Tx7�UDSM�gt+wB��`5ñZ���r�~�A.ɂ���öWᡞ�Vۑ����<�J�������C�S�:���?`N�j�f��Z~r�gd�F�FZ�X���<�ƞL`W2�%'�!i;S����ˆ�	ܮ��Q��0̞��[�A{�M0^<������	�u�(�v�.�&��s��v�.ra�<_��ֽ����}�щ��j�L*!�~�����kE�E���6���p\��Wl(���s��A� �<>��$�j�ݻ�br8|i�n�z���"쬓��F� ���
A�4C'�ٖ�$�g5W3"� Q~�x1�
�	�#ǘ�3�����2�P�3E�-x��I��۠���Q!�e�э\$�Y���<�Ns��[\ P�<�C6��륽��kLv��8ƪx,�*���������z�IG-���(�����ay����UøN��+��3v��<��^�?���|���
ed>v0�x���r�7Uj�
 ����*I�sː��|�G��9_R�\G�JM%�?�GcCx��3��2h��l���3$I4*���G
��[�ײ	ϙϏ�#��V�z�����N���U�)u<��N����F��O�����tؒ�#U���x���<�C���d�AmX���s���6bђ��x@5�y��C0?։-/|&;<�	%��s�.W�N�P69qA���r�9�yP�KC)F��C_�P�ͦ��́C��t���}\�c�~�B�)�`͈��cF�!L���Gj�J�UY��jR`+������Ϫ[��;��{ƽV�'M�/J�wi���a_F����ߠfB��8L�'�}�������hZ-�f��� ���`��v�l�ف����;�|<idL6
���ք�+�G���~T��D-�F�yx��z�M�A'�Ul}�	f�o�؋�E��,:AL��Ԛ��q��F3H_,��5s���涞JF=���q4�Ǆ�d˱��K����Hn)�Oa�;<�B��Sޕ.g:œ�A�ؗ������#�Z���x^���V��5�ZAG�|�C?��*Y�����_^�t���/�'6�x�d�Bw;���~E�KصX*_�0��OB�g��=zq�ov�4���OX6�:�C�)�n>U�����i���?w|�7��9Ov�MmA|��DT���{���xo~�⽲F*#�PC��҆@��M��in���@x��#���QEJX )��O�2�E+8����n�C4�܋�ב��Ѫ�O�_lѬ=(@��c{i�"����&o�'[�}���-�i��%7��c���Sn:�a��ݨ�ɯ5.���bH�0i�K�A�뢩i#�h�k�i��d�.āAkNLF���OƋ�6؁ˑQ9.G�]kjƥ� {�'�b��Z���o�1p�ϳ:x0S:��)�tm�@!~,�X��"�G�'O�+w�G <W3�S�����a[Q�"��E%Q��o%x4(m��eF���}-��<?�	��4+�GH�:�;'�����a���2�>���׋J9�I�}#���o#F@q�=������ql�.��Q}�f��0��.;Z���2#2�!&y�J�Ko�^�>�C��k#9���;�&�����E;?#��-���Ҩ��ژ��4%�rN��Îo�F��$�"�cS���O���]�V�h���7&��t1�JӀ !�J�����W]�������0C]�J��s�i�b�7g8��{��B����g��GU�n1�kr��~�;���	@G00�b���Ԯ�Pijq*��p��d�o������Y��|V�è��YO��k�ϡ��0�L�|I[�����Lo����V���o�i{�;�J�\��
�L?Z��ag¿Z���ۃ"zs]Hrl���vbllJb���|�w����c�4���:����
t������H�f��CQC%]��"9�b��T}�����k�B߿���Hf�ծ�g�M�E�`��bJ��Y����?BG&�WDU噾˥�����I��=Uǥㆉ�j��ā��'���hT6�z{�K���> �9�}�(�c�	�}���~\=��^ MߧL�ч�}tq�cCkѻ��`(���}Y��.�Uw�b$Z�zӧ�H
>X{.R1���S��?��
�N��ӣLAٶ��˅�
P~e�!�m)|X��~�������������3�9g��s�.կ�P(�*��层��EؔGU-�������j�e��Ӧ��ސ�bEH��?$3��F)�C֐:��/C�d��/tų�ä�2k���Q��t3._�F�h�P���s2���4}u�*@Er�����B���6�1�|�����.]*,'g/$%x���Ѕ	��3Y"c>����K��q� ��r*B;)G�r�I�zg���[J�52��5���?��6sP/1�	Z|�Mg����f�)i������L�?��/��'�gzE�UA�� �͋�c���0D�l_Ѯ���-R�9e����-0OZ��1�5��l�J��!�o�풧ax�Y�s�"�`�A9VǊ_]�N�&b��L��2�,j?][OB��4�i��j#�8oN]mTm����� #V-fs�m*%/�zt�b` ��E"Y$�|��%�qsT�l�\VPۇo]^{l}X��q|J`o/4���o��|�52���*dҹ:@��Fh"?�ô��q0f�L]�'��ݛ_��~�vPo�24���,,�U4�n��V�r\����J*K�~��������"�k ��e�ܭ�1�SB�Gmi����1c������us� �͜�!e�VM�6EOO~��CF.��������<X�E�7of�l���;[�4�� ���"q�Ȝ4�	�Vާ��D�q���CtoFSi2�d�+��K�a����&f��rE	*)"	��3��LCiu��,�ow~?@��P4Im��>��hӏX��"���c��C��_¹��*l��sX���o�8i�j/�9�A���� �{��WqI�m�=G�~j�2�y��C��[bk%�ɍ�xt��9��0"!�����λ�[ɯ�1����t���~n.q8L�G�֓��X
ϴo�-�����|��՘��NRo9X��%�����I�˙$2����a\Yw�H��a -�&/��op���EU:G�y�F��� \���z�t7���-l���E[��1�9F�����H0K�f��G���J��czYj]$��h�5<�އ�z$�bYA�\���wM����a+f���F\W�_$�z�
[����K���/e99k�3{�Z�j����!��W3�wz��b^q�O���z��z�4�?SYX��Ez��w��m�3�;��	_f��'�M	0�$���`�0���Q��64�����n�W�b�!����V��
��,Xq��X��v��5�����ij�2��-�6��zs� ���{),(ӿ��J
��[���f}�{7t�RQ��L�/!�J��3=�F�ʊ�N]&\-�����we�7�΍#��������կ�0x;��h�ٽ�Fm�o��@(���kL������q̘�og��+��9�dz��Tp���`@�k{w�|o��Gt�jx��am��l۹��
H�8�E��Mo	������8�f@`�Iw��9D��z�=�:����ga��@ I�l6�c�u!��� )Ͼ�uQ�l!a��Ƣ����#�r�h�)�n���W�:���̸���xc�y1pɗ��}ϥ����$��0�O���v]3r�­o��m^J��%���fxZފ\�0�!�R�e���;{�5Ǵf��%���Ri�5la�j�dfI�f�cE��'���<CINL���� �����v�]	l��m�y�5i�g:���R�[�q� ���,�~��	|Q��SF�_B���ZYR���8�A)�6�B�Q�3�K JnK?��{�؈���FȀ%�d���WY�'iK�R��L酔ᰏ;�K�m�t�C+�İ��7�|�M�EXYdEN�h��2��n|�oU��y��/����5͓(C��H�<}I��殬ɼ?��A��0����	��Tɚ'{$y�xå(���Θ��mV��%�[�u�V��/6����I`�����T-L�-����i�mK{�pq�!ȼ&8�(���<��n�1�}[���x�^�+���u+��x�eH� ��1���%�<H�(B������);Pf�6P��'�7�sJ\oD=�pT��������<&L��Du�m�g�On����\���C���f,><���l�)�Ü�o��0gQ�ڃIU��q�o�Ā��v{�L��?7B�+{��������uJ8�Q���7�5h� ��OdE��!-�[[�����
�=�d{��f�ri����:���^O��nj��!����N2Ό8]�>�#�#�vC�9��k �Xb[p�#�F|�2Ԧ�a(*�:�Xi�m^0�͡��@�yF|�ɕۧBD��[�����HS��"�������R�4}�XDH=���^�ҽP)�;���>r�ng�8���ӁEm6�߇E����wτIt��'�:�id3�ͨ�^a��M�r)C ސc��$\�#�[,I6pH��#���hES��Z�0׍:������B;��|1��<8g3h�פ�=膌���X'��)���MId�����y�8�+�8�z`���p������S��C�v�2 ���V�b�-(�bV�F���y1�����q��2�o(�V�2Ȕ�u)"����	��2_��;g�/��B�݇��-�!�v]ˠ?�<)1{���e�D��"��)I~�G�AL5<�on�d�%{�5��>�<��(��a���'t�S���%�їCX�_�����t�wJ���G�����|hh+vK�sM�wp����ޠ����n߾��VδG9���N��l*3�K�LĶ����H�$#;�r����B
��-H����R}����3���
[l�ֳp#ʢ�����x�q��n1/�i�a�'�'���0!������5qq��S���LW��Bl�G�J���ͻ	�Ŷ?���B��)P@�ʏ.��`zL�W֣&k;B�[L����R���vŽ���>I��+��i��ӻ�d�KӴ��d�j}�ܬ�l�q�pV�\ɋ���{m��y���DI��ꦅ�}Χ�6�e5ϙU�5f�=S���cܶ1���`o�@v ��Z�݌66u9L$p�-��Zȩ������M.�E�uKTwaN�;�Y�?+���s��QP"֢Pyv����eƅ�!��w�}��5_���]�$�l�{G�x�'��q�cDز�IƆ�\��1����_�N��HK�&9��K9sG���1JS)�#?�O
V���q��xn��Ax��9Rgܹ��g�AG㢯KT�z`��B��1��d(P�_Q����{�TfyݚwH��m�恋g$V�e�V�XX6	���Lz������py�ܼ�7�d��w�H�:�m|"�����Y���[����$^4;�JH���
V�¡7tG��[�j��, ��[�-ͮx�����W�i�T�t��-�r�?���p�Q��I�K��}���8�l}���*E��u�c����P��,Of3� �W�|�Y�L�;�l<��6o��G��.��a�,�A#^;V'�W���lBF
D	�ջ�@��5�E7�u���i4�a��m�I��ѡ�;y
�W��cH��Z�I��)˦mi�_)%����q��gG۫0!,I%4ڡ.r�"�Ⱦ�5��l�]y
��@�1�ym�P���h+�@�wr7����ꜞ�<�U/uέ	��Ѯ���9f��y�G�v�$BB�~i�'�H��X�,��R:�"7>M�8h1Ļ�k�10A[�.���RE�������k�q�b�~�=�s�.|���|V����c�y6#���p��;�hWN��}��B�qC�������:��܅�)�S��g���$`�0�8�a��)t�(�%��o�U`�uHc��s���o�*r�1�*DM�0��\�T�t�j$;�y�`)�y��r|4�$a�9^N��4�����>6��x�Sh^��k�׍YU���:ЃO���T��:4l����rP�D!��ŋh���ׇ܉^nI`�9`�*��P�R�]�� �]�q%�[S�=�k�Uh(�P��L!�a.]aG� ��r�;�~�8��ъ�5��G�i8^?���lVw�A��rEϽ��-�Î7��a���y�(�p
ЗC����3t�,��dl!6�I3/�a�#
��r�����Q�h9�~:q�aM�A)ii�)ﻬ8������ՠcֶ̮0q�/<LF'X��5;چ�� �"��"��ȑ�f�G�M��.F�P>6����hq���,!X��ܡ�SqW#䌛f�`�Y7����}��&�� o]���`��>7v�$b���t�\��_޶�.+�� 42 �Hɿ^?��)��{�u�����4Z(̑��?���JOg8�2)}+�m���/�� �st���0��d!��M[ӭ�)��Q]߈>#)���&\�� �N���	��y/����*�tm/�|�\���<��
��HH7����z�X�T#Kp�nQ���+YP���f���lJ������.�b�F˫\1��_D����Z.�bT�w^�|���X�>�*o*�%8g�jܞ@',*@�������E���T�.����xo}V�ō!U�:�8H�5��ٍ�dqj������H�� ���;�D1�m�?��@����l9�*. 9�����r�[��c�i��	
�x".Ɉ�Jr�"́-�H�^'9OM�w�­�R��p���� ����?gJY�|�W��+B�+:�*,��	O�1y����\`&���a�t�X�y�T�K���WM،��+���7�=3���ͤ�jiu�Û�pӧo(�84ٮi]M�b���e��2������J�R�9�J�M��1��*fB�iJ%3� &�C��.��~��T�!���m	��+{)o~xO��$�7�c� ������H� ��e��:줞1N�s������j��A�/�8�H�N�!���$t�����#cI ��baƭ�Hّ�x�/1�r�|�q�M@����y{��h���d�i[4���dX���*�mg�V�P(��q"%��t%8]�ʭXZ}S$:�}��Nt�3ۤx#Ƴͯ��F��|��~����|v���`}��S ��?
U.c@��A��n-<��a���}�"����U�e����Z7�=3��j�EqUd� �T�L�lS���wڒ_}ɾu�)^�ǩ��,2*8y���܏����9����R���|E� �o�����0������B@4�$�HcC<���.��b����NG�lS�{A��e�H����z��#/B�rn�'�\��C��>�H�m�IZ����v��jn.�<�&�m ^��5g��G-n�a��(�W�k��sٮ�Y�vm.U�_�F���8��A)U�ČUUF�?|�[���ާ,��H����ݖp�Mo�����Q��%�v������Ŏl��IW�0��D�����#R���V�8T����b����2X���4���d2;-�ծ�r�h�|����tk��E'b�Y�#�Q�^��6өG �~��$!�����}U�[�wK������L0B�U���"b���'����M�q ��Di%��|t��WI�.�����~��)�v&�J��O?�mP��0/k:�:���}E
�w��t!?��Ot��:t�7���_�6��2#O(�_��8�1��_XQ��1*/3�8�P  G�kldB�g�K 2۟5U�dH�60�Z��c����'���#����%�^�t �d��XȒ�>W8�4��1���ln�3�=T�V��;�A�̘!�~�UU��Qp^�ה���8���>�׆��"�	�P9%)��P�ܳr����lB(��{�$�dOI5� ��=��z�L�H#�̀���C�L�u�!%Q&�X��*˨�$~!"�[;��{P��:���e�4g�pgon��]E2��Z�����}�Ɂ�H���/��UHE	-]��d��?��YR�'�z�j?a�[h�h��t�֞��e�DA������?y�L��D9��r�8-!�r�"�a���fr7��.¼x0��G��p,S����%�8����;����;JF���7{W�F��K�w{�2'��5�I#��f��q���cM����E-���-']g,_rB�[ŕ��p��5�SŜᘑP=�%!beA��%5[�)�z��ң��pi@�zʣp;�C�� f�O�o{�f�X�HD��R�?�2�oS�O�c����I�WEס��2N��TjQb�/�1�S���TP�,j��WR������M˻*�c���v�/��[�"�w�J��єz��/yּA����O��8X9Hϙe%�Ԃ� b�G׈�J�^ �3@o<$Ak���-IѬ���x{C�7���C����|���,dК/�@�� �'C�=�#��[�za��ԶUQu2>��V^_�����7�d��+َ��5��)*,�@^4<�Iǻ�LSDжo�*A���߼�[ J�`�n����:l���%0T��Oخu1�L��I^�%�:�#�xs�ޣ+��Mɨz�i��خQ���}Y2�>�1=ž@h�&�s���z?�l`Mj�{�	\�F��f?����^�4�V0c���oo�;5/C��g��h�z���۰���*T$�$�t	� &W�7��[��ՓS�ô����d��LB�\1�4�����K�����Hr�MQ1�4�G�F��p�:4���?�ϲ�"������T�}�G���Eb�:�;%��'T��Qh�ȯ�.L��]ĥ��д�9I�!�T'����1i�s���7 �r ��gI�Br�U�{�,t[�^�C��w��!D�@�;��vL&������'I0�
v���B}��N'I�o\�\�u���Jm�t�ki�R�&6ϣ7��Q�~�z
࠴�8��dtn��b�P�x9�#��Û�/��f>o���.���eN������6����9�=�QM�CT�u,�B�x/5y6�:dv薡E)RM����1�-�U�"�p�B�ڲk�ؖ�&z�ET��ЈFZ�,��5�6m؂�����@��0��3J����Q_&�d������q�������#oq�%���̓M��W{W��w �F��69�`�',�e-N��Z!��m�D���R��{B������h�˪�cL��h{���^�lo�8�6����ַ�`~?���BىX���v�l��|����-i����Z:��8duAFTI
yTu3���nʙ���L�����H迩!��ꝛY�{�D��������F�pq]穽��Yֶ��蒥�� ����5eq�"�=o���<�K?V�Q;��H�"��TE�y���{�){�N��NKő-��Ҿw���e�Ԇ�Fu�Þ)n���+��Mh����r>uh��膦>�FR��qM�{�>Y���d��TyJZ^I)!e�x=��\�䉑14�Y����M[Oqe*ͤ��]�eT�����{=�r�G���}5��B�����5��e!�^�t��	Cv�1FI���������+�g@�{5��#X���T��E��X�H�0l(D�^�d��'���,�86Fk���p�M�w~0�A.��Vq~`�eeQ]�5�E��o�'�J8�6���@&�X�j�*���'ڜ5�1��W��Пs�����=���"���4����Ut3g��A�|8����)8�|��<A��ۀJ��>������ׄ(���YV~Θ����5���y�`�R��E;,�������UX�x��Z����I2M��f��۫����t+����=���=�9���L�9��w���?1x��}݄8�\��$�{����ܐ����b[�h`g�(����q�;[� Kc_̿����j�,��PʕV����gtF��u��me K��I-j&�F�[^}�},���2t�&��+q��׵�<���pľ具�X�gͶA�)T� ����.��EbC����б��7�7��=�9���'Cm��G�!e������ҹ��bS�jІ�1%�}�򨎌0�{޹l��"�������z&A��9R�ń^!�	.�������1¦hH�&4�R�����%�7��y��NDp$	�I������ȌC ���%oYwq�_^م�[iMdE$�+�,�J�,Il��2X���[��Fu��c�b4n�A(�̊�$�M�m�������t:zO�I��<[��^r�6����޵�f���5���
�{N��u¥�t�qH��@g��v���͘�7O�e�����$��eLZ��1�+X���稇�8ų�ވ��o�#������R�,�	Y�4ۤ1v�X�ha"ʧ潰
����_����[D��xB&<��0��'��&�J���r�d񔰙ځ�:i<��ɜ��u��"X��-�T'�8�'�$}|`��n�\�"�Z�EH^X����;�jF�5����f���YE8�v�;����d-fT���I#�G�-*��m��LKBϐ�y=����X�0���y��)(�y�5��i�Ħ�K�Mn�/X'���#���������T��%o4����!�ɂ��D�x�$&�C�_i����yq��U�!��o�TMvx��h`�m"rϨ��=-�MR�����*#y;*�	�J9aH�I�ŏh<���|$�����!��(X��y�3�?J+b� �*½�4��(t���dt"65������(�)+c[[K6��k?�HDl����6U*�V �N�bmG�{�}��0DÂ�E���sq�H ��ƣb2����4�#��,���Y�������$�nr�w2[DV�uQ`b����pm���ve1J��h}/�
�y�̜V�,�l0�*�pvm+U��xQ��-϶��[���`��N����o��@N���v�#ն"�d���O�	�9�Yl�O�O��xa%�̈́I'�խ�I5(=k;v5�lK��C��i�����3Z�Ra�|�N'�
M8����������V��~&�RFA�@`�z٣u�;]=��(�]}yyi�v�6�8�	��A�Ӌ���#Smʍ���l��H�^l�9��#�����.�ۯ�,V^�DR�ƒ��HG�R�.<�ظf4��4�:!O�J��݆u�ʛ���8A�Q��٪��C7IS0ՠ�Y��d��@�Þ8�{�����KޡC��N��]�^�v!Br����5+)��x��Z�,M�
 �]"��	�
W�D��v<o�_#���[C�[�M8���qKH�S��x	Ie��ۖ?�w�ur
�柉�ユ�`7boY~�{����u��uz ~�l�T���$<��`HuiP��`�� ����5Z�Om�3�/��j����4�겘���4��G�A�D��PL��-�����9Z,N����#��b�3��ܺ�]U �tG�(ˠ���� �7�qW�lR�8 '��^����0�%11��G�'��1�vGGBcL�_|���ti�)���>���$VY�&o���5Τt���>��R}/G������[t��9wW�Q락.�.2}�X�Q1*�p�c��:���M+�_3��$�0��r˞�T��?6dgb��Z<o@��cy)���ҟ��b�����H������r�H��6ea���n��@���D_�������cv��>���N㡪r��p)��ڕTr0YF׌D9 {n�·��l��м+&Y�F�������� OꍔZh}�9?�Q{��O"@�K�,�b�3G����`tH�6rsū���n����<�;5N�z�����[�!���bͤr���B����hj���u+��'�@Q,�	o��"�<�y�b����bsPA6�I�:��ʯ���~��\o�-�칃��4�T�]��"�][�����uϛ����Eyj����).�E��[j��%�ߊ]oǁ�.�k�YR�Ew���p&�P���q�o0Z�� ɉ_���h$�mu���[k�މFB���+��i����L��r��f�ν�
�)l��lS�M4'���	f�.����@zѾ�'�	g��}�l2-?iA�mq�K޴qV1?ųզ�5:Dme�t?�<*�@w�t=9�( ݈ɦ���G�>�<�C:����Ք�P�JX�p%����q������&Qޙ � ��pģ~~Q��Z���3��X�ȔՍS/�;�2�!���';���"��%��@�_��][F%��uw�	�;�Cz'��:��L>�ypl� ��qm�2+�(S' ���g=s6��Wp=�4۔V�H6?��&�����QM��pϝȄ�Cd�;�]2N���I��u�Ź;HzYuW��y1ѓ�˲_����x�,'���6�Ҷ<`��F�S�$�V=�a�b�ل�s���憾h9�܏f�>����Q�^��E�c��(G�fx����8~��Ӗb���ʇ����eD|U��ho�H���N^ڷ�������r*�1х�B���N#C�$��c���H\R�"��'a2��K�M´u��z�Dp�_H&$���kd�C������.���[����������5oB*i�X$�E������(!*�-��܅�[M�'�w�����u�~}7�E��v3��'����5� �`H.�ޝ~Vg�A1IL�u��!�g�JV���/����wFTc���T�^���ҟE���),�w�����{1�l΄G��y�ؽ���45? M��@��}F�&��U�X���\�Q3.j��f�ؼ i'���"^��j-6#�U���Z�%��ìE��l(B�����Nn�)3�#�Pąz�yj���5J���5�m�g���a��H89�d���Q�xqwu�D����䐽�����8~�&;�OՀ̐3�c�@�2�!� �̤l&�Xڗ��7w��2��R��#2�
��������#bw��e�Ti�6
����G�����R���h����$�1�5j��jۜ�$j��\vf�r��"���>	�&!y��4�U��� )��-VjnUU�p���Ye��t;�4B�;�۾��v�����=zִ!���WlÍ��G^u��0�X�*�v��p�m7g�Λ�d:�L�Ar�+&E��6��:�����Mf�Y!|s�j+'�-��Mi,�̉1��k�Di���rV�cz��U���a��WQ���O1C,nD!hW4��3��Č�3$g�C�_�h���h�.��Gi��u�e��diSӥ U�ُw��(Z̟��{�By7�_^��yL���3&�)�5[�����i���g���Z3�o߾qk�XCIgY�L���O�*,'�!��6�������}כ}IG����W&�m��)8.�_�zs���i��js~��
7��a�����tiu�B^m7��j��rM!w��k��I������̌M�$��"<�!Pg9��%P���4��!��ҫ "Z�#AD�7���T�Ԛ���"Ȳ���Rk�%�$��b#N���� ��[��
X���y��I�t�C^���g��~l���zy0��d��p��ȯ�D���SB7ʛ������ң���N`��(��v�jjqG�n�������U��Ự����a�'.���<��L��Y|T���x�G/����v�Z}�TG<2%��a[�%�S�ݛH���,I>W��ߠ����|;X�z�s=�x��~��z��6@aE] ��Ϳ�t����#k������Y���SiG�FG�+�޼|�Be��K�
fc{��!)���'�a����.��X�-:������k*}�`3��MA8��
m�٧ހ�	�x䎃����k�+J�N���g#������j�s% ��[r�u��Zv�#Ų�|�e�p�29�:�Y�CR"$^%��\��"��>j�����*R��<Y��V%g�IY�$m:�lr�h�5���ya�h�㶌I�@����R�Y&L���v�I*�=�8]��w��)��\G����C׽��s5�k���?������5<�^|�7��`jW"f�S� 3����"@	�Ib��I���$`�.�������_t�~.��Kp,<'{����Eg�-.��Ӽ�G7H�]�U�&c��ߥ�T�>�h�kz&�qaN.}��+�f�t��Y�k�<� �8�%��a�(��I�c��%�Y�ʾ�=�^el�Y�گ�P9_�/nH�TdDG����vo����_;K�Tʵr�]�	�7r*v_��J���O� ��^YM �'�S�.��y��1m��G���`9e>	��VOb�S���	�+.��ތ���$�Е�/%���<�G���l�y�]�&h��*��I� �\�ԍf=m[Ӕ��-����zd�v�\��cB�C�E���i�i/(l ��|��.*����uVx�w�yg�6٠���Ud�e��oR{@7z|X�%����e�z[<W��)�Ҍ�9�h�dFC���L���ZYP)AF�	^�)�@e�:�U���r��T����;�s�A'�ǖ���ϼ���f�q%��
�r��x�����������[���֪�Х��vM�9T��$fe+Y��)ʮ�'�C�z,��Zv�DYM�9�MQ�p�Xa;��da+�~���P�fTqi���!J"Ƕ9e��}�whݼ���y�`��zU�8�Yˊ>�<(.�3N�C��K�UZP����J�uzmq�B�PE��=O��ԗ�|�k�xݼ������帏���͇�I�]��0�Lh�)�����[]�r@_�X��]�O���tnk�c��a4ʄA`�1U�����.�����E�`��y��ʼ���r����O��������-��4Q ���¼;�&:+�w]@x6�*���T�ȯ�ꛃ��`$u���H%�^�����-�`�$��d��7����Pb�,�~���av�Fd��>�����L��RXC�؉�|����S�M��P-��Q�@x%f�}�����C������?��ͤ�X�
��ˌs �h�[�kd��Y�#E��+�dR��� ��2	A���k[��Z�"`|���8U����j��M��b�9�_��+����D?Oѝ�Qz#�,��A.u�q���J�����k6�Js�*#r_9�	2�ųѮ�K�$t1�9����}��4�o(F��:����u|ÅP0r }]�)R��~ҲX����OO�G(wO	[��u,I#V;[ْ���&׀�>�D9�$��@/����e��S�s�����FK������J2b���Y��7,���bLf���e�4�/��U~M�]3���3�C%��<�^{{n�7��SzЅ����0{��_�{�ʬl\��m���WF�������3oD�*�w��WP�'���Utխ��E��%Gg�1�wjac.|����ֽZ,O��>���J��R�{�w�F�If/I��������U����aE��J���?�=v����b���k������X^i�5.v�x�(K�
�!��8�:'D���K(S%�p�=�J�:)[�ƌ��P#}��TY	�QYT��/�l���Tb$� ���|�ÖQ����d�&�.�9�[ܠި�,����h<�jA 0�dd�%��@�L�Қe!F�ޕ�q���	 �P�+k@.SH5�qy��"���&P��)9譥�$Y�(��#����& �"���h�*?02��,��\2X(	7ۭ�ށ}�T�[���E�RA���5���`@X��%�<˷t�|�U���3�o�~/;�-�t,������ƾ�j�=�u������*,�2�2��Ø�C�݅��PhQ�
y��5Axn92J�f&]�1��'��`�"h}[�V�ľ��w��bn��X�L`Y'�4W�$Z{Q���v�Ĭ��tͷ䛏m��;~J���k��B�80�PI �0@��54ʦ�\��t� ��G���+�,g�;��J�:����6!=$�`�;��@��]rEvv�b*�XxA���r�Щ�"+��$�8T�-�ɁX�"O/zu��\v�_��V�jEJZԠBO��m41W��s��%����bK[�!cF��j���» Q-??ke�}��\}���O�
�l�f�jm���w���B�L�#���KQ���;�57�ǉ�[�\`�o of��,�I�W�8�XT\��݄�%��o���J	�򮬑��$g�~����EƩ�3�[(iBQ��� ��}Ó�h�	�1y�+������W�v�)��Ҷ��Xe*���W�ك��ƙn&3�2x���O�>F@�P�L:B�I/�@��?a+�8�l�u>_N�((U��M'q5����<�	�Ӣ�f.�Nu��QV�ື���bx�KӠE�wB[��=������t&'0��>��@I0Ϡ�0�y��D8�sxv���J�����)���_�P�1��
���%��ײxW}?2�f����gQ�]ChM� %�Ւ-���:�|Ka�ڃ��`���ql�}/��Z�����5�ߛ:T�̓�"*�e�;���e���{�n������}���㷸j?���G���?H(�����6f��e�i>���7�|�:qY֥VG8oӗ�CS#��b_�sa ����Z@�މ��f��M\R��!P��X"�����N��������nO�\�k�O00W���HM��i1Y܆!���W�/��,m۠�aU�~9!�����n�$��@�?{i��o[�<1М8�l�"M�a�Z�����x]�A^l5�̸%
��$���>:���쳫fB8��:"���#j�cEu_�մE|��������b���;�*�Aa>�Z��BEiŰ��=���X���M����(�:���+�0B���|F��o:3���ob��"�p�,�=]?L��ف��q�pU\��B��o}��A���~����o6�ն[H$�5m��Z=�/�0��n�[u����Ώ��&�E�� �UU���qG7���K�oHЌ�p���u�s�*�����+2^ks�Q `�T���/ⱴ��1g978c�StP�0��x���-�.G=5�E�Q�����9�(ދ�1ꋬl騖qe)�&\63Z�:���2�Ɂd&12��O] �ػ����W�+6E�s��|9��b����ޢP�˦eLw��J�]�ס�`�p<����ҍ���&�*�>~����c�g���N�ô/�x	[�� TK;%�B�竒֯��'�R(p~,�9k�\\yY�,_y)��tr)'��
B�Q��wPn4/q�\}1��V�O�4l�L�A J�}n(܌��MN(� ����Mi��U�D�$;;3
h������b��1,R^Г��H뗹Y;g\I�l5�#��U�M5K԰�%��7��;�����5�~"T~JwDLr��g��V̡������`2�)�i�.�������Wp�#��\��N�_:=lcT� ka ����H���Xsӏ����d�}sh�����?K4�!;F�j� 9�KC�(��~z�]������Y1�M��1��L!Ck�L�$�IL
��"��@[�v[ʎ<������Ĥc:A��fҁ���J{e ���U�lЫ�qf����`u/��&0@3�|H��A��G�j�Ě�:D�<��$y�")�����}��_�o��n��C%K�Pt��/���6E����``�l2�#�GE�CCà���A�ls��&���PU��o
�~��(�,(R�[�\��aR��ID�U�˲�c��-. �:B��)�Jg*X�*P��z'e�	`=~A�~$�c�!�LL�Pl�\ #g1��`�*��Β�-�|�G�����ad��u��+�ر΢��=���O�K�,�̸��#􁽚�eo��M�MX[���nV��%n�d��t�m�ځS:�6
g}�"[��IgJ� ���o�Jv�N=	!
���T�Q��eĸOxґg��`_�U��ܵ�UD� Ika�V���`v̑�ߏ��}S$�E.�7'C�|�B�.|h6T��@���� P1�U� �d����'��;�[��3�	��`9f%t�sw>Ӻ1�~?�k��~�2��a�)[i@�"�)�m���&b��UHz~���p����Q�V��In14x=E�ľ�����Q	ޜ���+e2g����E���at�.����|����SK���cy�����G�l�9iέ.����E��,�R�/��0�"ZE⭉9�#[��(��>qJ�����g�tBL��M����;]�F�J�:-��2T�SY�De,a�`�f������jO�k�4Z���ns����~ zw�6�1�De��� j��Ji���i�CcΎ`�<���{G�`�;��B����l� ���7}*������}2��mS�k�i�CN�P:T4�&���|��~�*9"�D8v�gK���6É�F���]�3��`�R��S�(�b#�Ŕ��ZJ���y�(][��I.zR���b�\�e��z�eK��03k�M�pn@y��g��2I�Xe���G��b�q�: ޲0n}��mc ��~��D��%J�B���'��#���cc����I� )��#�VI	<zj���X�)j=}Iȶ�uK����lv�)ɩ!AR��kb9}���yʷLE_��Xê䜨j<���~�GD��L_��py�p�,�U��v'�enUFʏ%��1~���Y�@��*08X=��sw��}��3����1ÈtQ*����S�BfƏ��+�6ϔSjK���w�RP�c���YM��$�5� y��e��mi��άآg��Fm	�d�a��򬫓{��x��Q9h��.�X4j�x���/�kQÇ2�:P���1A��W�U�J�bs��@(*�\{γ�9#4"�Gi8�RX#���h��h8j�!£�s@L�F��<�����mj��(?㶊�5�����gO=y��Hӣgqy�v�f�˸@��p1#�j@Ҍ�`Eqn�Ғf���eB`%Zԩ���
^�p��/^�\������T,�uppm����2�l�^���ԉDY`b�%����o�X?O���u��H
ы�I+���0�/]9W�O6g�j�x�tĄ�_j@ϥ�}�߂X# �y�>x�o�;sQ�����	���N��%��A��Z[`X�;l�m�y��v8�V_ �\~��[�� �� �4ٶ6���Q�~G��?�<�JEKN3�3��V�a��\W���w(ؔY~]�Rh�m�#���L`S�����07 'uG������y;�s���X
�k&� v.L�I���jJ���
����ѫ#���XX�gqXK���rMϭ�A���D4��7���97{_�zv|�su>��o�#g?�]�"1,�G����vJ���� 9�T
o��i'=��#/hr��2a����ڱz������ãR������A*@�VD�����\7�|��Q;o�ZBĴ8[����o�ܨP�'�\��;�'��GT���I@���g�ad�����,��mۑ�hga��^�%����f����9��5#r�P/�M~~��w�`�e]�/ا,�����wu�oi�J�n�����Z�o���X�mYk�ՂR�tVښm�[#���^�qW3�s�����'�,��3%�"A��D�:�}�����a\vg��|(�!/>���KrI��֎�.z�vI���s?ϱs�*�
�_R���d�����%&��ˉ_�"^�ςEP~�g����O�o�y9zŧ��x��2Dp��T�J{տ���!Ƈ2�\(��I&���Md�q���w'�� a���{�AԫdoҢ���2��,��CK���<������a�#��4*����P�c͕�u�D�r<(zB����/7�w�+w�*ԛ���h�e�r�L���0H�گ��!�K��H�O�aq�+��`X�{~fθ:���	�c�?�3���^�G
&��~���1dVұ.�9���O=wj���.ob�s>�`���`��@�����ZXﱶ@�捓6"��`���E�0�0�t+�rN�ȿ/X��wǌ���`�{�]#�2���7�N�����{��ٳ�W�j�u��^Η���8���������|�=R(�|:�����>`A/<�~�n�d�z��k;�1�� �z��Pn�ė��ͫ�cǍ�)w�o�fil[�Hoh#ٯ*���Z9*�������/�>��q7�LS�Y�����.Q� R�QymO�>
��I2�tr��`#��"��8$���u�=��YrA��C��%|Wb�T'm�"��_:�i̳������\ױ*�J��`���id\8K��O)j�K���[�����#�,�w��!��Q�zև�M��8�0�:������XOCf.��a!���Vn�흹�_r�u'	�q:��*#^:z�n�ҋ�-`�BG&O���9|���{�� ���d������W�Q~x�ci�$�YPķ����$t�W���z�D��=gQh�y���U�����	&��e�V�¤!~kް�²t0^`�fsn��8&�rXyL�$8D�)�g�?x@+8)U2�s�:���+$�I��"����d�RICql�YT�w�ō-�@�F���0��ir3�G��og��d({��oP)���W�K� �u�j�{���7Q^BK���F�.r-꘹�.������i�2I�@[H{6��<��ޘ�Bh���R����Ё,1�c����0��8���W�y�JB�j����ɶڇk3qĩ���@��H;_|�a�|D�\�4ɏ�|L��Q��K��NQ�N�ԛ0�[��v
-��k�)ɗ~!+~[KBR�uҦrP� S	�*89����p������:�0�R������y����<t��8���;���D�/	�}"�:����ۂP~X'1��1[�*ǚ�p$���I
�jE�MJ
�ؼ�5�����2��|�R�Un
Slvu)��a1��ЖهvQ� �櫽���{n&DO�����#�w��Y=��93�Ƒ���	d7?	w�-�uL��x�jj��K*�jq�����np�$�����=;ձ�m��&:<�0Z\�=-4�nE hu�w�@�Nd���O_�h�����w�K�P(���)�!��Mb���yEg�g�����Ժbh�M���.V����)�>�"�[:H�M��eT�Y��/�)h��Y�vf���e?M�oB��E�ēw�^}����[[p+�a>5���~�9�bD�e���b�C��;���a[=�m���S�"W(��s_<$Y"��;Ð	uT߀!Y�/�R�z#}m�t(�q\��<���Z���^�17Ql�`	�+�5I�s�7���M�Udd��J}56�o��J��1�3\��G��
���'e5 ¥�n��t�^ʖ���2i��U��y��rP��޻���s�C�8�#�灧���5ࠨp�|�y��/��^���~�$�y���������W�S�o|v�O- !�5�� C`j}�2�>����6T󖽙P�p,/6�-��@��w�YX��zdٸ��6a1X�E���y�/���*T0'ʈ��ӭG��^��;���J�*��A�&�s����
{�����{c?#�.}�:���
�2&�^��74���ض��9h�������	i�L_�-r�}D̎sq]L4��ō0@�JgJ}�>p\/@�6� ��G7݇�-;V�
�T�u�ˀ�h�ELY4���C�����
�@�,F�{��B��ًŁ����S��
x͛�2��N���d��d�4�:���X xkFo|���7+���a���Ѿ;���^���IF7�p��}��E]Lv�	&��qX���z{�i�Mif�.�M1|�?޽%�x���'&فG��{�j�0~|��F�Y���E��7۱ �?�sf)̎����R4O��µ���3E;�*���]�Od���9ч�oh)��R�.��[М���P-��J��Q�Iz4f���O��v�"(st�^�T�d�M
�OR�����5-N)��"C�k���uKtgW�����W��gU<䈇.*S�;^�s2�G�����5�=<���{C��i��ȟ7EڵS�/P�#�c��ր�>G!@E�-�C���{@kEp��1}�I	�r����-�0���a�E�5�!oa*W����z��mF�*D�3�\��T�����h0YJ�|	4�!+��֘��
w�-��w�_��"����-���d5.R�W�ǫ��>=]ph�_�i�b�K<_�
7��ڂĨb����+-Di���if /q�b7M�D���@�.�����%fD͡���v�N3&|�t �ʨ�]��Q59"A:�@���FI7��F�A����G�1�=d��K͖����KQ�����{���3�j�聬XF 
����'�R�W,���"�>�*qҴ�(b��ϦT�s�"Ze#zѤ��|#�$�v1{��b!�����*Yޗ��1@Ƭj�C�8/�/�����ʊ��S�����"��3xv���ݾVR���ޫ1�w�)���>)�FFoh7��o#X#fOc8��0�:&��������eƀ+��0�ru�0��U0|"U"��ۯ�������@�+TS���~ ; ��[���BMs�r��:�a�mǱ��%��ёo��l${��(�gK-���@oj"~Rt�����;�?�Z�]ȗ�U�9�*��L�ՈUW�O�̃9��+��e�>�\p������(*�K4LQ��.X�=guh#l6�	�}V�X�ٸq<
F�+��2;k�"8<H�{�嗴ނ��U�D������jNq�p����G�"f$/�0V�;��P�����b�!O�'��F�p�
����3���&}x�,�sG:
K	O�/}^2�;�+{�Lbcu����a2�1����p�� �ʺ�����ǭ�S�b�J^L���[��l�8�M(&>�Ď�b-wu|�0�h�h��=K:���
�B�П�
��izh�rD�e����s�tu�#��X@J@�v���6X�X�#�:Pyt���̈́4Q"::n����hȩ-���Ѷ|��R� 1�wؓ�m��?�n6�[	��:�^���* �F�o�*U�=�8)�;�,���:���b��kAu�8[[?E�۸i�c�Fw��z��4�O���z��NdC����C����w?=ꅝ�B�x������?'���	��`ï:M8�ʛ��M�����b�d�:B��w�w�l�;2�2d���"E�fđZ��ѝ��)ѿ[ ����,�_ς���q���=Wd�/ce#<�S	����Zc<�7��y�ӋpN�f"J����K���x�}����8q�*+�`�#�P!IF)�_�!A���ߚ�Z�j�l^a���&����Q����D���w3��±�lMсj�=�Ԧ���ʆ]d�IT���xZ�fL�=����%��Ǎ�n���Q���Z�E(������$l���$�m�����<�'֨r9w=[֤ЅςRW�b�R���@������T3��γ�7Hv�@[�;�NJ=}�6�H]Y���G�*���a/�)Ti',�)����&���-g�e����tK���c-����r�a���eT������B��J�heA�L��H%SƁ+q��yWH�6�I�ay)$�-Ha�4�yv�$���|���y��S�&i0U����md#u?^N�y�^���	�G�B����x�v20-��U�F�)�7/��<A�C��A�ȸO ���\���,ȇ�C:��B���~S�@q�}�PηM�!��	�Ĥ�E��-ש���6�W\P�����%�Jo�FH��´M�s9�i΍�x��ʜ}z>7���q�����zۤ�׏D7@��0%�O�쵤(��Չ������a�}��{�A�����̿�b*�.�E?��u��Z�'Kώ��=������`�{k����K��=�m����X���bm³2�z�X,�V��}6�b��ƞ���J.�6}��vP)����X��/z.���?�^�4n����g�h� �Sy���e`}!�+�JQ:-E������ {����/�."6�eƳu��uO�]�3HT�kJ!��TS�xN�,Y3�b]�e��C������zٙ �k����h\����y/<D��v"��N��v��y,P�����%@.�l�R��~��5��`������ 哈1��u�'{Nb�2kA0�jq�e����M��P��Iq"���zD������[���ū��	ē��٥,I/u�X䳰Zl�Z�p�8qG{��4Ek�AM�d�r'�J`{W�-oҝ��e^�}���%a��y�Q��޳e�#5tpQ�toj��v�_`pX�������>?�/����~�u�l�=��::')
��g�E���|[��#��^�Klx��HW���T}�������o�E�l6c��۰@?S~��K�9y֟5�{3��38{8si4#9v������'���`p� ����!*�.5�#�o{�X�����gh=w]itE/��H�}�sm2�����,����"  p��0�x�&�Y��?��I�=NP��W�ư�s��p��%]�m���/UJ �ׅ�T2�\s2�����"9W�*�P��H�0�u�~'|^ħ�=�����]>�(����`i��(H+3sG��X�M�(*
�|�ݪ%Vj�l�n犎�n@4TGK0vF�6�[Y$jax*b^�?n��D��`�2��>-���)����ĽJH�w�%e�co�z���(�$?LO�5Ѐ�d鹃:Lhu���e��z`延��x �:%�G��3Q���NA˒H@�3Z�|�9�$��K��bx_E/[���-�O�5�}�]�V������;Z�5B����'l����i����a ې����ò����I݄�/d`��=��z����&�R���~ {�X>���Qղ���[�cy`'/Z�,����#}��a���
'4}f����*�Ȓ��-mH���k}2a�;�t[d�����f�6n-��闥�Fo��!�4&��~t����s���*5�d
��������Y]���� �@�;�:D�ݫe��O��eu��3��5�@�i���!��F-��iV��ƈ5�o=�����oAwp>
���[��Ũ�P�ԉ9�����v&��Gxо1���*XQ0��`���A�;2 eُ�,y�����s���`+�@v�z�Z����7��2����OW#�9�^7�
٨	��ȥ9�hb._��MU�oUa+U!���U�n�$l-���E�x��=rXZ��M�y93����r���'̉��8^9ҳ{��3��޳�FV^�]��潫�<�l��N��xҬ2�pʢ�s��� �b����X��؎���Pf�-�LQ�5�;���&�T��jꥦƫ_�O�6
�\�'0�K�Y���2��z@�/
��	�M��v��r�w8��."�d�O���°�4= ��$���v����z�e.$%�K\�����<�	�
�O\'|�h(@�
�$	��ײ��^ĕ����HutEeȯ����� }k�&����U
YB���w�I�h���[03JxV�C�&<���s#��� ��r� 1���с�!��/���'�����E�~T/�R����L6Տ���\x�T����I�I�	����p��D#��H`�x������.N�E��,ͣ�;ֵ��]� >�y����.D���j]HH۱j�5H�!�t	5� �y2d�M��@�{q��Dbh�v�sTd��v�E
(0�#ڭ�����t�	�� �dG]����
���r�3�1�m_���'�l��0b ��w���[���ЃB"�����B�OZ���*ZkZ�XJ��j�{5Wg����0� �ɴ�ٺᠴ�ԧe��iCz(>���K�_�.b��'X��BlC����{��#�Rd�[�ަ�J�0��+��9ed�Z}Z��IAϹ�nm��Mą��р:������0�j+^r�i |D��3�$��i{��N<�a^mƼ����T5���')�qDF�ts�FW=�5wӸT>q�t.�Ҍ���@ �@�2����XQo����{��c�b�@�2��&op�e@��3,��^{��us��UUA\G��(>~J�#���6BH�b,�}谷WC�z�D
�=}ͭ]W$��_S��I�4?:D�4Ɗ�Zm��fkh,�ol
�\x�}�s�Ei�߈=1Ar=$ �h�mގ�Y���b>��.P�k��i�Q��II���N�f�����.)4bW?�J�`�,�ߙ����tF4 ��ڻ�v'?������gV��+3�-F#{�f��8���b��G�v�_	�>��B���@0��P]F��o�v2�W���nZő��M<ު���8Ǽ�!Y)̷V z{�Zd��*�i����mom|��IN5�C,�K8�U��*�We�'�d-,�����Tp��f�F7իbB����s����õn���<=��/�3��i��r�1���85�&�s;\F|�ԇ	>-�NO�rq�zdI��{�/���L#���j�P|����7�ш��Y���2d���-鷄��s[K�� �N���Mt7Y�*�7��CX�0��C��,��
��<E1�^��ofT�N���w����4��j���F 1'3Pʡi�����J�gT]&�/�e<~r�ؤ�%�.M��bT̡ �QMf�M��O�Ӥ�ʃَ^���Й3��V.��T�������1
�+ʕ��u�Ƅ���q+�e� ��?��]�b�����TE�_<H%
UK�������{��C������Ȉ�؈�^� C\#:o�8%W�IK��u�E�va����WXn4�[M�Q'�J��dD�@n2T,n߄�O@X$����GӉ�i��������)J���~C�BwL�;k���&�����w�`=�L���q�蒖yp�Ɍ֛~�m��'�:4�J�䗎%�R� 1��'����*��Xa��D�-�T8ܭM���uQwo�������3�[�z>�������ҝ��4��[݇�j�=�2<��j��'��S�R֏���W�ȫ����w'9�	�M��F��o<��VS����p�j�2��m�m~�i�9"���N��)C⯚`3�4��w/�^�0=�C�a�qM䴚Z��3��z+�������l�g|L��z�]�mTsK䱙ԓSb���
pwdNN�Jg��O0�oU��٨��"Go�	vC&���6��ø���R��A�o�BŢ��UG�=W����!(!�x�wg?<.ʩk(�L�~_?��ڰ~	;Ӥ�ϏѴ3�fY�f�9O���NB+�Cu���NoB��P\]����ӓCqN@k�g��9�z�ᬻ�ɵ����<��?�-��{SK�'pPs����$2s@�b�0�~��<�;��L�1�ׁ��?n -��08P�_-�hɈ�8��������s>|"m��C�\ ���Jm�I��WsG���^.u�`�r�ᇣ�c2�_���%�	�NHZm�L^Gٹn����c�����0zy��2ׯ�@0w�Ў>�n�ُ�ɢʤ_������ݢ&I�Q(P�/�;O	m�Q�hz���rvL��߲���O�`[��jT��V�2��Vt���Tؘ9ROMiʚm(K�����Ƴo^���|i�N��z��%�,��Y=g�Jb����0�#.���E�Y\�u;�D��zQ�A{��k�Dz�7�+��&1GN�-F�_��W��B�G�Z��b]S��-.�D��6��[E{@O�#�뾞�/_⟱�]���O[�#�C�m�(�� A.��+;��A��k��mq���ֻ�� �t�c�5�Rl��MbqCK"��p>�ioEN�D�]|2/?ġA��q�������H��#M�/U�
0���l�� ���Z�
O��h��R��&�:Y�Kq&I�~����L�mW�`�L�b��K�����;����%���ަ�I�� \R{=�KX��o�8X�+�u�m4z>��=n)P��M�]\�S'PU��I�`���x��I��o�[�.7��]�@Q���kA�h�:_!����R�M�Id��hc�yJ�U �{�,6=�`%�������<�� �õ��PY�>�#�����;�V��/�@+�a[�/o7t�,�#WBDd���}����2�i[bn�� ��#�,����%R��\�;�x������\�p��@
�.F|n�'��x��>ׇA����K�.@�Cj?a8 5���HZ�4Xx�.r�hՋ�9�1��M�B�߷�j�0 ����/���ZҠߞg��-��������=���Ѵ4$W����䳽�1{��%�"�J���9�Q�^�%4�舤��hI��5q�r�DO5	y��K�O����a��N{��/�mCv"���lBciN����w�~ʱt#r������RġF{yTUAeC����ε�� ���ɰ��#}g�w!��x�ϩY����g.�[�����-r��-#�D�c�1<@��� �0�|Q��J����?�;]B���j�}�p ��m���:"}�.:���6�/�@�VĂY���v���ip�<�����g �x2�Ѫ��>�a	�ho�ϴ��B�}�E3�*A���w�:�^x"@�����y6R�;@[���m�I��$~I��ߩ�a(���v��JN����.��eI�vp
37ٕ�84oގ�Bh���|8{g���B_�$��"��W�[J���ʶ&��-��#�vKZ�hg���`m,����1%!E���^�	,՚7#��֣x�C����vǜU[��J�G�{��H)-%�ʞt��l����rv�Q�}�T��(���8�V�	�Sum���|����$y�-$�Slp�FY8H�́���1�>�P�yKr5pHx�>�����H~:�q�o(	*4!3
nbyi|x�9x]~�J$�7�~�UF1�����W(e�d���8���w�����ȱF2�2HJ�kּ������G������l����X�������Ԉ�!�JC�?P����f�XYu�~z�pC�t'nr�8ƪz�<��B��n���|�yyl�g�'��N�^�����&dt����� 
���1>-����(+46*�������	m����Z��n~����+Z.9��i�	Of���r�+���f��|�;qd�7iKC�^ ����m���lK�ܸ�Ҹ�@
k�7p1����0L4k�R�Sw�TW�.l���a��?��VU�px��V��Cb��J�A椀,]�aHM�?��K=-cC̣3�Z�wV��ۏ*��3��IFP�C.jV�玟Ol�#X$~��.ϭt�>����n}�"m$U���<���Η*���+""�:����F��.\�Nפ*�G\D����h��a���c��4&?��	�� ���M/�p6��������G��2� n��c[�����4z�����-?Ǟ�1���מX�a�bI�H��S藍v�&<��@)��|�\�<jh�o�Ux�̸�.w\�Ա�h���=q����h�g��Wxk�ξ~EݶB(�������+��F=�y	�eы?r�����ӎս]��� ����S�"��^�SL[aD^��("d��?ZL)"�ȂӢ���b�|RK_Y�S�)Ij���gG�ynA��#���Mad",Ѣ�o��]�Q�[��r��@� ��Ѫ�/���	pk�yW�[_B�H�p9��C�f����,���I�櫱v���]�&쓶�?dtϬ�J���0����MȤᰝ�1�]P�ti� �P���`
,`�>Q��&J���ￃ���bL�9^���N4�H�k��b�Dp��"���:3�(p�`Cyo1��*�ɝn���4B#�����mDE��L>��+ei�P{j+?{���,!=4~�^k,w��>�d������$�<��@P+{9�: .�Da���L�/��^1C���a\M��Iv5?S����M�P��l����{�_Z�n��]��������}[,r�4���2�\[X�]޶��W�2֍��2�M>��u�#*H�m'���jM�<b��oM1� Su��g�kZk�{��q;Qz���6x�25!����s}��>��[[sDJ
���(4�H(R^ F�j*N]�`a�l��7C)hchMq����̭��N�a�A��kup��ԙʨK2"�Aa:w���rY�ܓH%;'���PZ��c���/���k6�v	�fdz���<��7��:x��p�1�m�+�sbR�T\�È-�^�d6+P�)O\V�$��.vm1
����Zk��1� E���8	)�S��<��N�U|�>d[���n[�޴�y��^���V3�<D�(@�/yP�L�n���h8�������_��{Vq�|�fDRS$ n�=I��z� ��5��!N���3��PH�\�ލ\j�n�6�|�E|����b'����S"�ϩ�r$��d��^y�p�JB��)h���T4�d<F��	�R3،G�^�~]��4�?��,-��5[f�l��dV5��s�l�[����Z[@����6�0N�~4�9N�{.����c܋<W����.�WI`�&�����2C�F.m�R��i�7��tr5�l�8^,	���Q��l\��Y�˭I=~���C_$��J��d�Ŏ�{
o�*Zw����bD �6��i����cw�+gv���ѹ�zَ.>�vtM�&ō��`<r$��UQK����*�m���J���y��[a:e{;������c���b��Q�~�:�a���RQ1�����y�A۩�f.f,�W��0����^)�w�Ì��8��J��S�u��@8��}�&
XŀV�&,�'f~��7h>�C��<��F��|V4z�� r5�t�cF�7zIɮ�%�$}X�$h�5�`d�������/�$p�0J\��0}��r� G�C�-�%VShF�g������C������)W��oK��N&]G���d�O;A���+=���]�R�&�	h<@�J�4+�� f���Ctz�$zE��#aL}�t|&Y�sh}���<�����ֹ�����S��m���Q��SU�9������5�,N��z��C���1JĢ����1��z�#�����_�|�?<n�^ʞ+B�E���}��I�Ƴ�D@��Q����p�J;64[*E��l5�ੂ�= W<��ցa��K׭�7��m�ud|�,���DF�-&�u)���Q�ku��V�wz{Ib�P���y�v���h��)��"k��^&JV-O���;�h�Zy��|p�
bq[03qau��3ン�/pQP�ֵ�>z4�Ԑ�laV��с�H�d�5L;`9V���)דpgʼ��"��)��u�i����E� �#�4}{��3�1�A�?�c֎�A��pb~ds=T$�/g��GE������;��x��}���t��V��Z��"�cy�p����ʂ��%*�D&"�p4�l�QI�.��pG+��d��(=ho�[���F�M,�b�~^LF�d,@Ʃٿ��q�my�JR��#\}��a�f�r+�iu���XG����M��BKC���qO�~�jDta�Yz���jWj U'B`шi�'�؁c�B�<WB�'�#�@U�'��P��aHv�"��Ăk���v�b@s��;2m�0qd;�%Jā65���sh��u�M-�fai=Ub {��જuyC������J���� &��*�*��/����#&3`y:�q�7�� M;Q���@{ eo���r�9�p������b:]RbbS�c���Tj|���Bf�jq�#r�O9GZ8w��~���*¡i�6�$y`�:���T3��"���;Ճ���Q�jUh,S�f
ӎr8]V�.��ѱ�![�Pv����7�>��N��߉LЖ� ?׮>�jVV�>Ck�`U���Uw|����J��䚹%7q=����G�aJ~��H�!��B/_�����Rz��T~�����3��}h�h[�YWc��F�J�L<m��q�#%=���MS,8zx��I�^[a �����A#-C��e���W�Ӭp�������L{�ty!!�%�F��<킴�Ŵ�4�����)���%yAm�rc���姊X�W���"
� ><��,��S�$(h��"N�NuPA֗��?y�>�Q��͌�O�8f��O�%�~��o����lb�͡�F8È?�߿��.=T���S�ډ9��J33�Z���itq��dʥ�R	���A�*����v����Z���.�Ƞq�v�Zo��&��\�C���_&b\����@�H�p���yc�roR�,��Y�&���OH%ս�8�Jw�=*4�;�y2�eC���jP
����n0:����r+�Pv���,�f1<������P4LA��E ���ͭ�\���@LH_
�A�e>k����>Q���ˮ!�7A�&�����i7܇yp|�ZZ&� 6PA�%��w��W��B�Ay_�5�3�R4�k��w%� V��/���̛�9`qx�CA�Wq�,
%��/�� �GՅ��Q�	Qv��c񲿟u�,gM�F�C�U�����O3t��Z�2������L���`j?F����*��c�	�$�O�@E�yVm�Y�]�I�?A�G��� Ǧ��`1��k�/N���6@����
�n��獛0ݞr͕#��N��g�����C$TR.T�q�+OW�����<ס#q�JO�3;Vr�Ot&
^���6�#���s���)mGN��<�#l�K��6%j��M91k��d	,�+��<k��\�f�Y����Ιv�V,sg��L�e����S�Ȍ�^�F�.�����,�$U���� K��0x?dI]���%���׌
�_�9���ӟ�<Iv�U�C{!�����6Y�CtA��A�����p�%��a`�J���qB���	ć����qVoafg���3�4����WI��>�7�� >�VF��ԹeP]Yup�IVgf�ZЊ��wOAux�iYM�[7yzB��f�(v��;W����T(��4����/	�SW���:�ީ�s�BkD��iH�rMÂ�a�蝷��n�Y2T�z�:��lV�I�;������x������i��q�1.J������RX�[�_�H��f�^��G��"�`
���[�YUc&h�={��y�����6M��?��M?�r>]b+V5�<���=�܀R6�Y�q��)U�"�o��ԧ��*J�Έ�>"�΁�2-�x���������wN�ȫ�~K�i"�8�Ņ���R=�F�Zfd�����`X\�����&����u�7eR������.l����c"<�rǻ��!��������ET�|�k�|�D��w|k3*���f�Y"l���9�-%�f�$�C�y�5Es����@�Kfiӹd��+eZ{����pg�r����P�ږ
Q;��M�C�Ƀ{�;����*���R)
{!��'����3 �![�W���#�G�V�ۃ�n@�38�@fp�Ɓ�f�������j��/�rq��*� E�vv��ǔ���p�Ir�ʛ�_��M�9�2�HJ���|&���)Y�q��#2HE�����ᑋ�Q��?xM�ށ.dǤ���cu�v���.΄eW�vΔ�m�=x�E��M�E�~(�d)�M�D���G
m�C!a�	O���d�W� �4�ڨϛ^�e�����9y��x��슌��/K.Ϸ���\.8T�������)�>};�-!U��1l����淳�	��X�5�Ex������p��Z��}:�N���*x��{�ͭ�\�f�j#��\I3Z}g�(�/Vrh�.&u�݄�E��E:J*��kP"\]�����D�Ű��X*�g=A_Tc(���#���i������ou�E�D�h3g5�2��l��w��{��$��Z�tG���s�"��P����{�	�eED�Z�{�ϗ��xCϧ4C<Ocm �%I66ؔ�9]GM�-�K΢���8�-�ɝ����l�*��m�T��Q1�Z�Y��ą�I��ls����Äpǈ�_li���9���+�P>�d%j��{�(�h��x�}�rH'�r4o�Y(4��qV�V�[�,��5�E�eG�/� u4
R����T�����y�+s��~/H�8*��.�y �� 8v��k@h�u"�aIՂK"sg�
놰`s|N�Dk{�r|M%�g�]� ���������M�NT�B���f��"�r㚻�I�ۆ��g�B�#�]ҜE�
�7�U�I�Plq�g6W�6�G�	���ii�=����4�WK�HŚ��V!�Z\,�6�8%a�~��0��+�y`ȝ����w���JW�Pr��y�n�p�kQ"�ݲQ���C?���0�;���-�,({�r0k�����D�����[V��dl�buN|��Ϙ`ك-� ��O$i�0:���]�A���4� �|�^X��P����0��y=�{g�T����mg���}S��u5�E�T��wX��~�^Ak�*/θ�{򚳎V�؄�vsZΰs��$r�7ޠ��h���'M�K��ך�T��v��?O�
F�}��*�8��]�4��.�jҘ�VA{�_.�mQ�X�:Ҕ.sNnn������}�� @��v��\@O�@�$(�#VB�sG����()o&�|Z����/��<\�Iz��/��(Xv;�1^�ײ���P�f���V�_v����HRw�(1{�3%2�BLW@B��yD9��������_x<���R����GΤ���r�,z�a�ȅ6�iݵA8{��r��(?��t�H��Y��N�Pdv��f0~���|<5)N�e���Ö߄}8�������e����ʚ����u(�c�č'�@i�G

�ZHQ��w�@���fp�Bqh��RC��&l�w�i"���� ��A�}�t�����h���Ɠ
r3O6�S�Cx�n��R������`)I�������r.]G�&ω����g�6�`+��3n��Nw��H��j�T����}�z�����{a�AY�B��>S?�z��a���k}�P2���OQ�S�I��{�U)OL>N�Z���9�ֵJ�Xu�qc�3k�t��ɯ(�z���b�7��Y���y�ɶK�	JE.fl�*)?���2�����"^�r��k�|����(k��܇;����̓uE�y����Fl,YCl3=�����A��j���ܕ�i���v�%�eѰ��o��.bHL����ok���Q�o����.h�\�C%֨̆E�0R��;�A����9=��gOG8ߒ@�9:�[��z�T3m�F�/��#�ud�+�;:o<2TO�=>����]�װ1z���jr���N~Nr_<O�gڴK�cPu�ϘeŁ���?�i�vωrD��&g	�w���Dy�P���3��a��uZG�9�&��pM��߽�����9A�ӘCXT;��,j�]>׍������3ܝ�*���0�Gݩ\_���������6��Ț 'R�q: 6�dO���"1��5�=��8�)E�Z�DV�7CH��9L����0#�n�/�ꅟ���H3a�[ޠ�"�GbU:��+�����5m��h�
E:!�k���?΢��ֵ�9�&����]|��ۘ��d}�2m��=y�)ٖd�2#�b�{�N����;
��"�������3�1�k��^�Mܓ\��4�@������m S�����:mg��Jh���[W>�z�:�h�J��+I��4�Ѹ��N��)��2�T�@������#*�H/�Cvv�L�K��:Qz����M��L�B(��#��Lm�֭(�t���l�#����@�F���p�-DE���J�Uf�m�9>כκ����aq���Y��mZ���;���.�m��w��SAZ�4]�u.I]��pϱy�;A���y���}���&�8H<�7�D��xOR��;�=%��\�����q+o�n�����pʥ!�2V�^���tq����,(�_�͇�*��zі��4��|Kb�G��v`w�j���}�o�m
2Y�MUהM��^��8��Qfv�[5a��aAX�����l��Lo�\�a�������P��jP��D��~Fe�J�*����l˵?̳9a��Fvl�uJ��i��f�W;��>�'$�)�N\�� ¼#v��UnC�1����d�N���)�_L�Z#�ڕZI���<*N�3��0L˱ݰ�[7�?K	ˊ�%U��d����Gty�s�V����e�=�ꔬ����}�e��]uμ�9R)F4?�>�8�<Ɲ�(��¸�VO� �~Y���v�BX���C�E�Wh�������l�	�n�`ch"4JlL�u�c��J��H�����Wsá:�����T��=]"�A�>�օ��5�lM����b[�B�<��h��f�O]��w��J��������X�ް<ꃔ����5>Q�qz��>���{O�7j���HɄ���,B�wzw\�%���l�J�wI��:!�6_��$�UX�'N�c+�S���#57����';�T��&2�j�^�5{"����q��4p����&UE,=���h�rj)�8�Ԙx۾��Ca�a�	�2��}���jH����xѸݔC/�Yñy*�ƫj���,g� ��0V.�ƯVi4X���Z�cϏ�9���7�`��m֞M��=�l����C�8�P����S�8�V���C��09,+sT#�;�+�sS��U�Ŕ�����R1∎�u�A�ɛC3�P��?\�U=��8P�"-̑�v���;��WR67��N�%�U0�Ƭ�5+��;�rVKgA\X�u��%-�s3z�4�"����a�0���-�����T7z�PfZ�3�%D��cjPK7����N����5�n�A�����-��#���L�l2�]!l�T��-��� �����E�X��&B\�[�Cqjj�-�b��`�����n�j5����:t����"���hD���FkԶ��<*p�\0�Uri�O�ۃ�����P��Vmɠ]��b�MC�:��?�<��Ev���p�2(LB.��IJ.�v���O$7�C��������o�k�uv<�?�y;�P/��;���~��͍Wֺ ��B�B��A[W� *��^7�+^�VX�P�bb���;>&����6SO̝c�j]���4bze9����se\�u�|���	L�${�´������E�䛖����մ�HK���V�w�veѫ��
���ρy������#g3��Sy��j]<����|��L�B��\�(
���(�I��)��E"�㨉5��X��˾t���pjo&���^
1�P�G��iw6w��־Nϝ-UN}�d�2F�����qle�5Cus1�bY2�E�Rm�l ���.��[f��a�$�bھ�i�w�,�o72!7#�p���BՊ�B��x5S�D]v2p}ُ�{�(}xt� �WbxɦА9B�pǚ�_����Z,�:����5L��n>���I�C%��Ĕ�����y[rB"�N~	ؼ,q�z〸{����_K�m��0FQ�\����kږ�Z@���"���?�LM�m��!�z��K�$[q����t��!�D�hԍ7��]"�FգV�?��@��d{��HCk��	��8k�s�T����:��xđϪrsa~��5ǈ�cu��M��}* nody9��m�� ��N����;ݚh\<�`�bU�7O�l��8v|K�����V���mp�;��k���}L%�ky�xN� &6w����P6��&<,řDP[�rߋ����p���Z�2�[�@fsI�/H�q�.��P>�h4�?��0�G-�k��Y '�3�b�-����z���9ѓ���KE�xJ�jH�V�ofN�V������זM��6E����b�8�EjrgTh�lI���^��a,z/6
�'���5�W%jЉ�q��wh�y �qp�^.�4�i�hs�;�Vv,$��c�.*=�y*�5h��d �i$�1��!\��0l�M�����zk�tO �P��tu �2k���G������A3%�S�`�6�/�OY�U]ˎ��fG�?��ě���d�\��M*au���/�;L=S})e�[w�J�Ll���y'`nр���"C��զ2~�Z.FLf�uB%��ه���&ĭ�/�Q�a���ܩNe4���S5,5�^<)p�&ɋ`�Y�@6)�Q_�YV>7�%ղ�7�cH��f�/9�"5��e�h�jX2��$��1&󱽀0�bX� ��F�����)ֽg	�h�$R�*�=�8��벱x)�#�ਤ�x�
��<������ ,�=e�5�X�lF��'8���<���UP����d�f�^S\����	#�@�?dQ�Pd��M�\Z��� .�v.�wi>�J&  isv����B�����C��j��1�7�=ve/����ӝO��u*�C��> �����[oi�Ϡ�E?��;��l��8�gh��2Q@�V6©~j@�.(f��׉�y��$S�0,J�>���(\���.���(ԟ�;��K��w\�cV:��0Ƶ|�\��O�Kc�Nw`��;�x�Ea8��&�����&۵6��*x�KS���УCe2%��)(�F�XVy�7|��l��<���mn���x]D��ʢ6�1��47�7 �Қ�@q*W�=�{^�~�١�r�Yd>&���L��78�SO�ؽՙ�t"-�DUr�<; R���?_�	�g��EI�8<�DAw��z�RJ� Ȫ�R�X*qv~�oi?�ߠ�҅����oJ�u�pI����@]��G�9s%��b^�l;Ѝ�ɝ|`�^ݹA��?%��f�޲�ޝE��+�&ٗ�O?�q����j�H<��U �?8�_��A�dm!w��c�~����c��/�-�S�Dǉ�d�-׌��v��!j�nڣz�^��*����#7,mH(ꤲr���f�NF���������(4�f��#��>�@M�&� D(�"�syê���p8���Q��Fݖ9�ϫ�e`$��{8Mg�J�=��+�&�A��<�7��6 `����?'U��b%�@��@�u������[d�{L�sA�#'<�������;�%��a�?�A�v�J�Ԃ��QM=ݶ��z�Y[��7�?5:m�Mј���H*7P�G��$��ܔ��{3F����*L����k��42i��R�%�ejq`t6�I��*y��?��A_լ���f[����]�I�=��/Ì�,�8I��f!b�a����tv��2x{/c/�;�G��*ܞ�Y�Ô����ƕ�����鼻�*�k�_�n9 1�OK��m%
s����?+�w��|�x��ke��]�$\�@~'�r�c��&�ڊNm�E��
�X`l���rX�������|Vo��#~�68�
4��6J2y���ܐ��SeH�0$8D�dt9�x��+�
D��X]�}��f�q0������?�,A��{���#i=5�M�8�L׆ʭ׾�tt���˒ۉ��q�W��ٱa�T'�Ⲏ,Ѩ�YP� -<�/�\�V�2��Bf/�Y�x;@��}���H��䦦�ʝ�mb�b�g��7+��~�Ç�c#��vR����(�͟��$n0zD�֍~q�dÍ\2�-��g9�U`��f��0�����7���.{VH����a���:8<ԭQ�Eo�W��z䠙jpu��9DD�]���c�������J��e�@dY���T�}�����?.2����o`]�j���)C;���emO-`ٺ�ԺP�#�R������P���l�$� �:%de���ʁӿј�z�/�"�]�d���&��
��5�3�b��/c�o��,e�#r�T��u�������]�j��c�̧�t����p��e�pr��S���YD��yBmU���LJ"�ǌ�#$j�et�/��2�"0�����x~���Y�H���D����ʄӓ�u'r#�9�v����R�-	�Ҁ�}������јpgj{��F�b��B��~%�t۳��_Xi/�%h&�ڡ���KόJ�ʠ�W�a��n��٣A ��E�O'�b��cs�ܞYչ~�0��&�p��a3/~-*;�C9(��V[B%���e�C��g�.��ro&�?�5����˓����0����r/Y[�Ҕ+	*^��|��[���8\H��`�Xg��@w���I���A�+��#���MG�va͹�hR?
i�Z�f��pWd���1 �[�)8~�a+>�s�i��:��d?HP�0<�VZ�O�Y23����+�����یtS&{L�t�1�!uś^�#$)���f벂��U$�Xu�W�����X>��e��~X�_p� �oр�㰏�}�;yE6����^��ԃ�W�N��� �� Бʙ�jF�Du��a��Ũz�*`�q�d�>��b�*%�b�i�4�v-�c�m  �R�u9=#�Pk���ܒG��4w?|�F#fl����HFT"�|2$ ���~���������Ĕ�P�'�*M��J�xlV�;֟!�l�ٴ����D��1��G _��-�oĬ�T�=#����@P)P�q��O�+6.6�zI�>\i���ڀ�PP���UK��=�1��p^�Jw��ԗ���!u,�~��-$��l�,/�?[�JĞ����_�h{���_q������8	�޳R�Ѣ)Z��:�l�H	�6���:
w�]��.�ȡ1+�.O��Z1Eƻ�TzG�$�����8`7u���\@Y��\|A$���T��;����R�.��^޳��Խ��s�"��&)���a��ia�����˝�m��/�^0v#��@��/9s�9I]��>�F��%��K���m-��5֩p���G���A�g�?�"2$/*��b.�J�gHi<��)�ދcʙ�˖�W��{���#�W�(�q�l�\��+)�T�
�t�i��=G�7B7��.��7M�����[9�#rt��p���>�=2Ts�i�9Y�J�ރ�*�wP�\��u�̧�T�ai�v���/������A����)2��L -�a�Z0���KC�xg�ӆ�$�l6��� ����꨷��8���� >�|����$�k�`�I��0u
�@@�(y��'┽�q�u#���<�V��U��E�	�D4@X�����*䈶�m�]塕z~u��F~�����B��+����׉P⵩���̲?�Vh��N_�vO_w�s�ُ��J<eJvM��\����I��
�F�(��������&5�^vF�2dXu����Fw8=��-B�u�����n�8/Q�k	\9�(�V�!��Gs���%f4����9ɡ��P��WO���'�	��6�)�-0�h9����<��Q$��!�gf���Ӧ ��j/EVa����2�SIS�A�ٕ<��&�eE�����.i�-��	{ 'Wv (z�_tM�E���$��X��	a�].x��`�Y�yK<�xIF�w�!�� ��{ʕ�O"�(�$�y�A��Ȫ��j�Q֌�X[u�A�(1��5|��Z��1]r\b�9IM䷥��&G) ���x=���:t��w�r���uC!�o�����+�y��ްBs�'�<�#O(�2Xq8��?1�6��ϳ��Ͱ�P6W���8���n���w�`[��S?�����Պ8��;I-C��#�H����H����K���Q�=�7ܩf:�Z��*�q�<*e!,:�n�feSc��A�Q��:v�,�+r{�}ކ#*h|0���V9���Ɵ�W'���4�Ԕ��:Lv���DqT�Q?�֟���a�;#�E��@��g�Ʒ��ç#"y�i���^�0���k�_1D��dS�C��/��l�������o*�k:LZP�b���>`�X<�k�nm&��K!��,��u��I��<�JP���d׃�����ъ��«(���B9���n������+�c�>eΘi�48��?G��eI���������^(�=����	8%r�W(��̣����:E"�e[�q�lAq9y�Xq��.�~���1b�V�Vk���%w��c����'����^��	&�� �	��b�O�NٹGe}<�M��������'���2Bޢ��꿟%Hs�����J�ҕo1�L>�2��9j"2�O��C~5s@��]fvԠ� �]h����7�����k<����L6����@�H�O `J��Wl��6��Ѳ��N#>�*�S�	E�#*j)�}�{��jS��f�F�ϲՍ���A�����ƕ�Ȼ���P$ʡVp��]�� ���V��'p�Ĉ�,����^�B_ j~��IczP:N҄N�^���S�'�p��9�FM��b�p>����y)�U��M�����P�uF;;��$w�K��]���8x�|K��j��a�4.q�3��E���$��3m5s�[I�(¼WS�R�+S��LD?}�码A����"��%���_�6�v2���l^��z;���F�i��G�*��3R��_o�� �GdޚO<�&'�Ve�G��WH�vV@	�����Q������ÁD�����\��r�\��rG�oW��E*E�!��-w���@�U
�h�!�ymK܆.�E��]a�	=	'�7Z��-�� �%�g����'��6�Z@l���A&�(~i$o�rxd�7��MG��|������Bߔ�2����=�%"�K���2�b_���������5x
y�Y�&�JuĶ�� ������RկVz��9�~ͪ�C$�28����㍦ �����> �2�{������J����pd��Z�)sF��dD��J%���3�a��H��Xͽ����ϯC�x���F<eןܡ�{������T�
Z��
�P�x%_�R@ѩ���E.篋�����Y�$�AG���{�|�@+����$���c�nW�P�w�\<9���߇�e*� j0��{����� �V�J��}W� �I8Q`I|�]�+� I,%�*��9��g��c޹�+h�"g-O��C�d�֔&��񫏐g�U߽�]g�p�s˂�D�
���l����x�2L�Xq��c�׉-]�-�uh��z(d h�I^ �}e��eњ�	I�p���*sC�G�r��?NT�5a��R�i��3|���FD#�3��|q�O��=(IwL���s���R0��ȟcِ�B֙"Y��ܢ�J�w�(6l{�yfG�m�*(��a���o���k-� �So��O>����L	s19�M��d	`�����!>�ſ�nz���6ӷ^� 8X�K��7����CKlmyc�y�9�4qRQ�˵~��389�rS�B���h	�!v�1҆���gu�i��2B\+$��`H��Ӕ_�r戹l(q�Mc���Z�g���ŇC½c�_E+��X���3l�[7)ܴ��	S��n��C]Wց'N9�d�R�unX�O�E��H�|J�A�n����[б_"щ���m�ϲaV&+�?HZ=^+�q�I��������.���`uE��'��M��Ν������7���ە���8���������d��BF]�ѽ�:�xGu
oc}�F'>�3�āY��1~�HX��!/"m��M' �oasB���V��+��1�"�F�T�9r�T��,+.3�d�+����`
���t]��g�wG�~b0��0�u�Q�ʘ�5��Sf�	Z�N�Tŷ�C�9�����X���~���܈L-�ݲ�kPy</g���g7�MRɕ��#�>0��	A��iM��v��b'��e��bGm���w��_�k���o���a}�]�,�yG�D���9��6�2]���3I0���(=�l�r9����ң�� /��#����[�
�7�
�E�=~�PJ�y��܂� )n�vNv�n�z9ʹ-����U� ��h���Lcu�};Y����K�����O7�`�����J�h�d�H�7�J\�+�u��i���:��=G8j��So���4��'r�B�R���z��Z-KN��it�ˢm�c�i�i���wɦ@�������@���B�p�	p
�Z��.$�:a���-$���g�@6���s�-�"�mZ�M[R�Cئt�W�{��ΐ�Y�}aN@/��pM��x��e���p���*,��M�L{��YuE��D�ƥAo!�8'���R=��/�iqD ��;Ӎ 옭��D�r�oM����no��W�T�9~�V[�*��.Z��"�']u�j�O���'��q��e:pI2����|���	^zq�ʫ���9�q��\l@�[�~]��I�,E���]Q���ƴ�ͲN����h������/�0>��m���^g͵�P֦�}�	��������QJ�ja�/V7i�S��v���锃R���H�n�-��u�&t��1�� ���<B��ߙ�!�f�Ӧ~�)��o����*r���Ϣ����-n/�K���=����~׹;A{*n.%����:���A�5J�Q}�#��q?l�͚��T�W��Ч�B�xo5�q�Z����-�>��ZГ{�i{���.�NK�rI��?PG�����l��������פW��Qjj��_R����+��&���pKg�7��)!���`z�q��+���Ј�a-�>�)��Z�2�n��N�ݾ�+j��:��$-8��W�����!�j�1��V�{�V��kS�R-7�4�r���og3�`�O�s�N7�𓼟�e���� By9���6@5�.��x\}�3(MAD��utz���D%�O�9���?����=�q�%�Zx�ا�����Ix���S�ت�]�;j��,�O���[�h�P��P���N#lBpN�ɇ�_o@SS�a���(_��VX� `��
#Zs�ɏ�$�����G��0��.:�CM�d�5Q�8lK���8B�޿�=Yn�y�;g>-}�4·_/I���M��w'�ciS]��5�_E�D���kC.woX���Y�bb�џ:v_�5g�Ժi� ���l#�h�����xٟe	z�Q3)?�Ln0!�h�h~��38Co�w���,�#�%N�P�U{(5χ7UR5�g��$"��Mל_��g��%;�}Ծ�ʒ�)�4/W	;��eg]Nm�UO%R,5�"�s*{�sK��y�G� ]ၻ�v6#}�Bfk^���h�'p�:D�S/p)s鯡;9c;��V��TO�A��hˠ�x5�3<��OV
n^�̣�RDw ?��G^Y�������T;u��.��QL�HYu� %eu��_<]�t��wIs~�;���f}��W����;��x���:c~�SnGW 0�(��FRh1�Bͽ��4��)�x�5�c�c�]�����캌m�O������4�y����D�G��2��XY��lĳޞ��|(J{��.����J
�uሠIF	U����ЉA��[����db�кlP���?��0���/B[\�ߡ�hK�`�xHIQ�t�������Ф���:�_����W�UF�uW�F��R*��|���]��E����uܓ��f��*�w����RZRI�d�����Y��)�H�6�qТ�6Fξ�ag�n_��ԑ~�h�u�$��p,m�0���+a�L��ܽ��*���8�m��$jbv㨸��Ǐ��3�nC�u��ֽ���tK|P�9��Ψ� l,�S_G���i���o!�RDՇ5�D��␵#T�bÀY�x�d�
G��md�x�%,�FUE�����]��}�g��}�X<�2i�&!������JJ��z�2 .�c���>�Q�:���F}�}Có&N��n�N�1t����+9�t|�!��p^�^u���PWflMz�P��r=wHs�
�A�;k���:��γcy���G3��{�m~4h��p�p���p�'4��jh���4�7�nn=���:6�ߊ8)(P�LEcQ*`t�	�a����S4�<\F�_��9uӐ-|@}Wb%�1�b�!kHCG]�e�d��~����܀��?EM~�`���p{g��у�@�k���<��-�d�m��@�m�8����(�Fp�S'�Wv������s� �5��a�d�9Ц��	��Y�%~���W?�JK�	��j<R��I���}�Sj/�P�Xp���� ��3x���'��y5��vaY:Jo�¿,�s���s`�&Xo�,`K�r\�7#�
)(&��Yh�,أ"yi�4���
��PėO�C�o׸ߓ��o���\.�~D.���KE��G4ϛ/p��]���ie�˷h.����h��p��ų9��3��[1,]׿��|B��o�j �|{��-�N��H?�v�_�-vh�| ��v8�jNPjUDg��,�0��f?3��]�:�fSw�^-� 1VсF�ZEFY�.���RK�b�ǐZ�ծB�
b��{��k!9M���q�$���H��@gcK���E���$�H��p�c��D<³���;���=��%�ՅhE,��4�a�-�����2y���ݷW~�����[b˹�  N����W��Xꢽ��b�i�^�N����s���Vv�M��	7ލ�M+g̼Y(*R��{��,����ܳOzZ�H����	̋P���a	��r���Em�i�[A�syd�����R����Vծ�?�sV�%1�K��A���Z����u�.��3,f=g^�68�y���ђ�hvq�L2�ҙ(;�]��Ǡ���g�2�WqoYɰ��8�y,í�خ�Qh��Q�P�з�\
��3��~��kY��$p  7���a�]�> �������."Ӧ�]��f��+G)	��i��4*�vrN��T1�>��Y��)`��%a���0��k�0�Y��tC�%�k[~����i<�L#Cͻ�epۼ��Kay.́~�	�(6�H����a����X�]}otzϼm�hQ�X��[�^�/g{PCc�<�,�w��6S�0���������ζ�ݣ��{<~Y4M!��b�����F�wb(�XG�V��ȁ��8�ݟ|0W���[:�M�c�jq�N��}�YR�����= ��{�tj3�J�L2�C#�JT�]����}��c�7n�N����-�����s��J琖����A���10�$6G��©2��P5O/��D�yŎ{ل0��M����ae�)��]C���a��9�q�ޑ!p=V�e��V�n�NI�)C�v���b�Hf����:j�(�E$h�[f��R�����B~��,��Q��}4�:ee.������	�ܠG�x2����$�Z�ؙ�0�	NӅ�Qhސ8B�j��{��0�V���:X�w@�	C~���[%B=g�M:l��=.��hi�Hb�N�d]�D�(|>�=��w_�
 RK���ɃW���?��k=�n;���'j �~#��c���
}����������)艥aM��e{b����Fx��X��Mb���~7�Y��O�F�Ko���a�W�/4�ǝ��0�Z`h���m��I�峑�±����5s�a#l�75�a���lc䵕P���$5���'��9����&��4�g~�/mi����W���2D%�U���sы�L��)�P��4#]VC=���=�ǆ.��hSp����]a1��C[%d���m�+��k��J{����o��{�����j�!^�9=D5���_�ʯ�(�I�= �Z��VsX����w.bU�H�k3��'b�P/�9�yڧR���E�ܖ֊ �'6�^�?�h>!��4H$}0�h��q�G�&5����6gJ�x������==�uS;�>��&�L�@O�{�E���A���5E�)?���@�yJ�(��%��ۋ��;���a���C�cԍC Q�	ݸ�h.��k[�/rb�iq8���D��� �{Ĭy�����s�]�	�SۙL��Jz�g� �]*u�b��V����(��=-L��z���.b��\�R�f�fz^�b�L�t�Adk
��C��TG�!����	�lr�J1�ۙ�=���N6���
p�^�05����)ۇX��U\0ޚ
�D ��dM�@����d�Ŗ7Z�Ȃʓ�c4���"G*j�y����5
�2 u��`xK�ߡ����酅���c��<p��k� ��M7N�g)u�Z�S������@�@����� ��U�Q���Q]��k��X���X��y�S<N��.#s �� c��,�%���h�
�
T�����5Nw�'���xB��<�tUF��q����	&���ч��?<�I��Dr����޺Y���gODҖ	��� ��d���j���%���Hp׌B��.#z�|<��xA̤J���`�=JI����Tk�;�r��m�2d�>}G�������~��:6�T���6��)�9��.-(2Wf
T ����'Lu0WYϦGO9򴾏��O�x��Ng�Uj�r��'R��6�!��j�A�K������0��@D������s*��!٧������XE�����t��G=.l�,�&@�����UxjL1E��"�\�ܵ�%�d0��D啘1C�C����P{`�1�>)1ѺZye��xfv��BҦX��N�]��8 ��.�lASg��q�'���iy!�����e���� ��k�4ɐIq�4�{�卭��r�ߧj~�bC��}\H�l;n% 'N�2�j��̧T[Y�Y�]�7�1*�(��I�Ⳑ֑�\yf��&��a4w�����SU�4���z]p��7�X 1�h�!�����!���w�S- �d#�)?��bRA�f_�N�*� n}���IX1������,0��}I��o$��h�݈z�'�����_��^���k}O���0=�1�i�B�ٗ6�9o��o݀���{p�K0{�ꜾZ�$���\�Bz���g2�r�̮�CΑ�F(B��R����=(����w�͏|ȁü)35.����;8�nK��~��q�Yr��]�Ga�}��L�mN<=Cb��V0�_ˌ��AIї>]m�}�֛B�'���U��틣���:�)�D�EIL��bŖ^C}�ZC��oo�'��A��3�_k�s����	FU�\=�Z��w�Möӯi����C�e��/.�YL��8�R��i3s�H�V0*%�a_��V�j��"�� �r]���@	��$~jm��w��r~�q32��/;PY>{4H$��l?����З��QA��%��2�nPÓݫ�T
����Zr�����($�lv,�u�3L�r�P_�I�F����w�A�[����=��hK=�7|�&7��i�]�~�P��S_)�����P�� �n,����]I������ǰ�%k�k��`��Y`�.����:��U�S�`wxO��Au��;���V�(�j�Qҷ-�݈�$�>)��L��C��cCm�O����D�Pt���Jez{Y�>�Wy�7x��<,���2W�ϿF�c�F�!���b ����v���@�n9�~���{D���E��12a�}�l�	��鼹� Ig� ��r0h��]O،2��i��C޾���)!�[l[]���p�#�b*��:��5HsD⏳Ok�'�(�,�F�3���1�2���=���b���9h��x��I"�x�Ob�IA�
�X��N����VgV��?��w���$������yeʧ��C�#]lW1��>�� ȹ�-GvK��Xb%�����d�0��L;�9.��(����~�ɩ�Pn6���_oz�t�p��
jU�L�Z�|s���q�{5��9�f�L�:Fo(D���L�1a�����j3<��"_��m�#.�v|�C�lAX�����y���Ł�~�Z�@@z:����ЛJ�n�=�p���~�GuJ�i��l`���)_js�h1���8ĉch6	CL3�t��	M��gPìy���Ǒ&���o��ݪy�_�d1Ag��A��� a+�A��lf{�'�~f���į3;B6܊k�O�P�3����=�%�(V�o1�&���:����]{ä�`�w�O�^�˩|`�K��4%�X�[��ӰZ��C{z���{i�!^N�on5P�\ �5~U�Bm�	@I����U��k����֭�90�N*�	��I����Ij³�)�h��8�����Cu1vlN��p�-�䊆{>�'���D�G垣�P;bϦ�RZ]��}��F/� ��$����HJ��b���8��C�� ���"'#��B~�N���l������R�C��?��4bNv�8سj���PA�q�xj�і�z����_�����g�� ����<SB���;ӻ 8���~^��Y�
x��0��=�>�*�PHsh��x)t�P�7y�l7���߬�G�Jkm����n�.���a5g��9h�;J,��.uT�4\2�ܞ���]0�pO�K�
PU���{��8�o��o�{_�K9�:/_j �0�}$���=ɓ�\�C��T�}����&�Jqn;��;m ѕ`�������~
cY�yωt���ŕW;�0򁸲�2�� O!̻�@Ŗ��[���a��x�3G��ِ�g����˩B^K���P�jͲ�1�H�̜�es��s�?"!�QLB�d��Bk/:� �w���V�3{�M��Tu���2V��!~fg=��1I�$l_P5h���}�8W Rhω�R��Ŗ�sk��J�ۨ��$�JC�j�7K��s���Ǚ��z�e���HQV�f��|����h���m��Y4J����lIAN4#�g�N߳�۽�~�s
�8�{�'a%X�T�ļ�5��6w�*&���=�V���|���a��'u��l���xR�г�,�*�Jr"�Xa�d�_I��.���b�����r��z%0�.N���"��2��h��7��Hz��
P��Vĭ��C�+���'�9��Y6j �ڲ��[.�h	����L�@�(�q�g�m4�	P�)9��nF��5Dwp���:�K��cIUu�0|�[�(GW����ɚ�-<�0-}ֵ෴�{���tr��͜6��,���`��������3�Ѷ���4��2�����#z&�Дtf��+���R�PW��d�O8c������b���k��wzw%"�������Xߑ�w�4$�s� }���A��̅��өH�f�R�HA6�\��k�L{B-l�;_�p$BB��X�� _�D�hwD��%�f$3-<��J1�DM�'�����������L4�=���~|���%��:q�����Ӷ ��Ռd�%��8�V��b����.�(�X��p�:�Gr�MZԷ��m'�V�Æo��dsI{��#\
G���X�BٮO�#k�ɓi����5X�:ú������8w��1;�������Ɨ%�q��"�辞r��>�����jaـ���`�'b�"��cK0!^���*H�������B�xS��!���d#�3x	W�e̲�vq��p���-���D�`|/¾�p>h$���ߤ�G)���3>B��̲[i�*։� ��m��}v,7p��m;��XY�"lF�|��Z"�b��j(����Y8����=/e�>2"?�[4�����4!����۾�;l`��$Y��#ͅ�a�N�6�t;=� ��J0��?������L�ط�Ƭ�����z�Aˋ�<
C��9V�O[���Y7Q4�Z�iZ��}'2�u��[�h~Tu�
5v��o�;�G?�f@�J��?U�y�ߧ������|��"_���b'�=�B[ R��b<*1��96�BV1����M�[ٟ�r���Mr�'ف`��a���sR^	�(��X�� \;|(,�V*9c�0�yZ�[�m��O�{��� a��3��	]97_أB��������~ff�C��Lڍ�7'�h@,�)��)��v���EX�SN��)�}CkjL��w@M��/���������J�ڽK
]Pq��6���Wb�'V{�6����N�YG|h�= ��&�jc�/�V6������9�>N5�1���|;�Q��_I��.�)�[4���}{�
nT�%7#�o�3�s�D�|�N�Ln��hk��vU�G~4�Kbq��eTN�ҵ�/�Ŗ>^���g�t|F��~x[�g�#3���^��J��\�,�J7M6��c(|�a�\���q=�9w,:�qZZ�	�2zV�it�����,�U���P�h�I�����*����{�U����Ô�LEU>U�H������k賙��.'�hfE�%"��얾��U�Z(>9��G��1v��d𔄥=�Lһ+�N:�$�#*�4��OhCIz�27�S���N�?��D=�m���O���������hȈh?�?Y�Q�1�J�
D"�3��������u� b�#�>��m�W�c:KeA�	N[a?���< !�B`5h� d���ǰ�L����ӤAe�]�d��`I��c1gC���>w@'�'u�����=TPi�L��_wb��ŘB����k����w��Z��d��ܼӡ5pq�X����>�J��90�k9Ʃ��\�w��r��uM�[hU�u�)�&��!>%*�ۣ�L��"n�:s�?T|:P���[l2v����|f����\S
�J�p_����k�p�w�j�fFVP鉂���Pi�?nH%
h�;�J*O5�n�������{`�J�1�:�L����J������ΫBd�Ʉ7�  �ʞ?�B��ȋ��%[�iA{��f#i��T},����:���g�K����$I$�� m՝ԧ,(N��0N���|�;��a\����N�WR�(i��S4�Bߖ��xR������%��ѕ����h�)]���F΅d���BaO�Kϴ�`��Or�'p��x'�&"ig~>B�7��ګ�����I)�9"�~6��Zc��a*��eׇ�q������{y|�r��eݢ�k�I��>�,�����Tj�Ah��B�n-I�3A_�|����xBKB��;���4��@(�3�y1�y��s{�{x��b�S���ޒ�`h�I��ۯ�*ٵ���)���W��<��..E���T�����j"�nJ���*'r &�&@��TI�H�n�=p8_�g%I�0ݹB�WJ��Qj��p��K�-&�`�-��0À�6���MR��1iK���[q!z)�>�e}�b���X�fC��ơ��|�P��Ȝ(�<�B F��2�̹�bX���bZ�	��va|Q���ĵ�={�<А��M�����5��U��S�����7ʴ�Cy&QVPL�\�omi�zIJ�묭s�`?���7}��X��,yK~��,���,m��9�Uak�|{n����!t��0I�;��׳��>oѾ����VD���р�c�b������RKW�7PK��H�Cr���kxMmV�k�aO��2�y�dz@�2�Y>9W��Y��_NPV�	����P6�V�hb��Yԗ�y6_J���P���l�|G�k_��X��Dpm������>{�*��tn���#�m��P�1���8"/���B�؀�Qv`c[罡�r!ĹT�q���Btk�=������C�I�'��޿p���\#mp���M�.�%/���Z{ux�\Q4�4�o?�P@wvMc�|������p��d�|��' �m�WIv���ء�h0�96ζ��VBb��u���au��T��͆%��޷4���,� |�q����a`�7���x�a���ko<ӟ���4v�=�I���7���wB2|���kC �n�t�H��uF �H��[?@M��ʍ#�vF�i+�DE&晱���f% j,���?�W���(���7�bEh]:}��~.Of�5"�v;2�n��卼�Dgw�#���ƽ��I�C���8�28Y��{N^�D��F��ZA�	%�C<^Cni�M��ų���S�-�#���$-��.(R�o����[#G��ڱ@����.��>�u�#�
m��G/iPc"�	y�5�!z���$�.8+\n�(���vٔ�^O@�5O5��3��j�P0d�F||�Iw�g��q�zxt��t�d�bD��s�h�ɴ?��3�[X�f$��.2��9���vW'{����mp�:���&ZY�rm�N\��3>�=}E�Ņ��ح�D�@ų�/��Q졢{�MF���lGÈG��4����pS'�q�ϰڡUF�e�8nl.��%\0��x��g�	d����D1�ʌ�R����q��4Vq����)l�+����"y��?���'gc���:j���W����2��H�Ͼ3�����:Jрф;��ٌטn�jI��/O����FÍ6%��b��z�¥)�ܹ�ұ<�1`IY��=�6�pU�/Վ�!�9��g1 ����+��\Z�S�O�4yE��l�&>%�T aT�d�������#i�so�[mۚbb%k'w���Tc<����rݗi#w��� D����F�N>� Ho<A�@A����������n�[
t�mǘ�����bG��.Pnb� ����7m��EP�2[�y��C�&_u�G"��.�y��Sc��5%S�ѫ=����u"��8�6���vƟ���Z�B�,��ۡxB䋣t�G3������2���U5��N˳�c�ꂎZJM��!��wV��7'ϙ"q@#2(��"0.�襤ΉU�N&�;\�"�<�f!A�Yck]HA���Oe�gI�L�A�X�c�`��O���>%S�O�|fR��䐴4(P��";�v�$�wP�.�����!�������oJ��5�
��>��)�$cU�m�E�Ϣ-��\Y�T9/�`��<cS��\���6���8�2$D��M�i�l�)±t���e5�$^����/�'Wxq���$!w@�rⱙeq�(˴F�<��a�����w������5�>��d��e�$���w���̌��5|�cR���&p��P���V�O�������b���ɪb��1� M����d^ei�.|ƀBb�����<��nh����)��рC%��ŧ����&��.�(C�Д�,�AGU:�=l�n���+k�������<7���`~vSh�C��dʯ�~ʃ�����D��w�4��)$�4�L��x:m�ܵ_H���*�'&l8M����9c��s����gF�Il�7PL#�-e�a��B]i�bƾ�=4B�ɂ�h	1\Ǳ;�X[��OH�r9/rCAV��Z23d��g��s���yϱ5�J�"���
 q
����<p�+�4Rfu\z�z��Q����v'K��|�T�'L-�f�Ԅ���/nm-ᩉ�a�g5�����X �< �>K�Zt���5)K�_�����A�+��{}O�?��iei��\6#�V�����>��+�,�ɼ�kk��@2v9s��Z��'g��:�OU��
���x�Y#/lIa�1'��M�x{��q˪m)�vk�hUM�
��l��9h�����#��7���z>8�)�vi��翍���F�4�[����R^<���/�j�X�y���O�f5Ly{ꈏ�K��q��E��*_޳��B���<��ʌ�'eLfV����dc	( ӣ7u$u�C��[D[�:��0�Dݿ���)h��i�Jz�,�� �l�<�ꢶRf�nNx��3�� Sܩ�b��~�Jْ�<���Υ�$�i^/tz�"� �+�C��T=�
����/ĩ�
s�RQ�{-�R�	>��*@��0ef_\� ���f��8���z�)�Q��-[�<4y6^{Z��5�I��Ã6��K���ԟ*U����|T$�Υ
8�U�+S4ɢ�8�jg�Q6xPqym����1^B�*�p�2����\��b_���7P懷m�"t��\z�'��.\݀@:?$��p b�����Q1���>��ב�/	�'�[+ӊW�Y�b����Bv�b=0ɠ��u��r����I��pg7�\�˪��{nn��b.)�3��y�6��E�l-��'��re3�4#�ä|yaT�Α8I�d�����S��W�ր<_E��z���Ja��=��?k��Ey �u��]��p>-�)�4���1���df�#R���޶�N6������M�M���y �hH�CL����'jՖ�9��HQei��=M�R���k�{$�١͓���N�2����}a�4����E�X�H���Oa������ͥyl��J����7��H|
�1z�k�bK�8��r��z����|���~~��M����3�E�z�;i��"��!B}$AW�kކZf6���p2��ƒN�%X�!d��>׿;BGY����'׊wdK	H�����k���o��N�,D����x#2����a�������%^��Ο*�غ�
,�t<8\"�`��T�e���G���k�¼ЗK�6���Va*�Ff4̿�)���3	��96�c���m�t���;���`Ӎ��tK��+�� �g�0#�>����?g�w�h�\^����G��	��@�&W��KIU�,2��=�ST���a�Aa�+�&o���Hϋ����.G�����2p`J�5p>;����s�Ҩ�GkU��2�r���co$P
�7������l�TvAK�¤�{�_'QH�x.;B�dtW�Q�vͪ|���4_F �3���	��:82�Q��Voތe��B>��@�����@���(�BI��3�'V��b����5�Sr�(��ݿ۩�\?oRnF��nmL'O�r�0�vohГz*�)W��-s��7Y��ÊȽ�����H�E;��\�Z��ᕅ�l�&���
�,6�x*��6�B�KpC�I���=,�����0�O�1��3�|?�l�O&�Ϲ�_܉���f
5�ߔ�*�^���3?|3^�&�ӳ��_�٩�4{į�ŔNʨ��mV/�<>��?s�i2�h��ʥA�={��l�F��˰�	��Odܑ� &,�Q*�:�3E8��	)�'��U��}����
���-|���}R���%B��H3J�X嘇�B?����F�ؠ��6��b�$Dǡׯ98���)�)����x��P�fH̏u��Z,�ry>43br�+��xG�gj��3�l������Y�5�s}ɩ��b�R[��떬��ؘ��d[ǗX��ª���ِ<��v �T`��%s3cb��|�2nf�Q*g5v�u~�X���	C"��m�s-Gc�����Wm�P	�a
�0����6�%��x'?ͩ�ۯd
��lFE�gI'Q���z���8K�L�]{�T���9�꩏�V"�?Wn)��z���LU�YC�4�Ю[�Z9��<�G�oF�[y�/Q��&�+<�d>�E�r\x�3[�����#�k]^�E�FyΪ����P��Z�a���"�彿�Y��� -^..�=�����=(t�%�F]˩H7��X�9%��*
be];���y��OI"��`��5d��+��t�NZZ�뵫v|&���ǰ��`��B�[c�Gp���:�t$(�t~�R�����Y�>�]'���cL�{Zл`|�%Ns&�P ��h�D(zS��/r��޻�0����k�'Qϧok�,��Q���8^I
��v%���K��T@L!�7ed�\^�ǭ-�,{/���g�~���2�i;|�X�^�7��ć�Ʊ2� ���~oB��9R�S�9����RfX�%A��0��	��T�"�1�m�:��U"ă8Zz�c�G�����^#%M�ey_l���K��-�d�v�O�����Ϻ��݀���(�{@����g�����_�t�����o��.��1617�9,�Ƅo�X �|o�΃=�`�X��Y�Vb�S��'J*�"W�N�s߰�^�&��m1�/&�����^s�T�uo�� �:<{�x��3*2��,a5�w�EӼG�%�z���H��%N:
h�}\Ō�~����;���<��r�����r}�5#�'�[x�S��N� �qt6�������
ڛ��b2�.
���=��Lj�s��^�������zW��(@���ŀ��V;Tͮ�8���=U���D�P޻���̖��}v����q8�[�SM=Sx�@A{�����1'G�S;0��5�I�go���k�t0�D�76Q?Y8��0����ච�r[Tb�B�8`��9�RQ����C�1#a��wtqU!�/]�XXi�t`t��4I;���\q8�@_��A�`�^�&B��= C��xwШ�|<�M�Y4����(,�>h2�2��S<�{��4Ps�w�I%̧*F�g��!�mV��"R��6X�c>	"��"0���&�ǍqS���Yjn�&���19�t8����k�02��x�=7��fA�&O
����v$�{t�ad��oWJ���j��W�;��T��]��O��j53�rNk}r��f�C��
[�YP�0�)H���ů�ȝۊ;h*�\2����b^�F7!���غQ��&W?(�?�B��.�=���Y��&�@�e?a��7�S0�ĉh�#�r��+�a!DT��6�|��ͽ?��;�����'���9�q�m��W�CHZ?�J6 �G����EӢ��%բ?������+� �X�Et�W%66Lh|黑�]��A}��c�|�a՝\��gV��3�iwRO4x`���gQ�(L,�PjLJ����Hir>�ܮ`��_
3@�8o�u�j0�����t�1��T�����iJ쨌����m~Hf8� o��(�V�����q��@lR����L�E�#������EQ��F^�m���\����bj4
u�z����Q��~��(~�a�k&C���a98+���z͹c)U��Q�!��5ӡ��^oS��j�s5;��y���<X/�Ǉ� �6�T�J�õ~.M��E�6��.�i�{&ԳF9��s��O��#�Uvb�󶓒�Ѡ�h�N����=�GrA�&�,&�N��^�~&Ϊ��d9�pd�L��י�,�*%u9�m`��>[�R5'�*qb|�gq$	�0ԹvBBvk<�CH�b��2eFd�'�~h9�i�p�	���ϒ��L~�.b�V8ǟB��t�4���	U��T#��ϲ�d<��,�Չ�1�<�E2�p J��:s�^A���_���=�v���\-�g���!�U�y��D�~KИ�h�A_���y�JgȆXP������������CLׅ�&��n'�\Q"0��K ^��Ϲ������^$B[�2�����E��T�sg7Yݹ� 
-Ǖ�z�]��C�}d��Y�P��p��"�q[ �c(�͂Q�<O�-�tǠo~*ɻ�Ϯ;�@�|�M�*Sܺ�-Һ�;b�Ә|�&u�]ؽ鱷5�j���jZY��· v�N��%�7��R�ZG���*Y(��t�C�+���+@agf���L���Dbe�VV[6_�dg���r�Pm�!��o5�GAwg�D��w&����y9mCV�%�B~,r��A���ı8#��:�>�^w���h�B
�Ì���r��T抟���y���|�<���#Ӝ�$����W�Nu7⼯,?� *sv��?p�wj[M+b���8�d7&�t�戈��ɠ���Jt��α�q�?��>Ug&q�A�Wd��ܔj3p=dxۍ0��q�+%����r����C� �M���#��d֌�$G����_����w���+��=����T sF�	�;++~k,E���N�(����QE2u$�)C]%�9���@����n��L�5�Y��f���1G}����u䋻ߓm^�(��l�-�ş�����]h�<�!��$^�+6eE��O�}�eC��ٗx\?X��O쭱~�M9 �}����uIT/��o1<&���%3mjc���[�רm�E�u7�r(�N<�`����� ��\o���&�������C"	`�e��yC�?�WC��Y���n��ٟ)��˦��8�xY�"�r[A#�@��ퟸx[f��B(t�JCO�dh;�_ ��(2��ͥh������ ̰����c�yK���)�ߜ��x�uc��Y:XYQ0.�[����|�Xr����	�����`��c�)����,.��P/�Z�̼�b��(g����As��
N�$�+l��	��1�ŵ�Gcc���f��+Ơ/M
��ӾQ]�S�>k\_��rm�E�.A��g�㫨�J3���8EЍ�hʩ�����=}��SN���57e�k�ံ�T��(O��%s���vG}�#��	�@�/ �/̄W)x9��Z�Fr�!Qo�@��S����PC�2�����e0(�"�_�&���;;������@��
 .�� Aipo$�9�d�ʌ�+R�RZ�e�G�7�e)�~���2}�ۖ7��e�|-p���(̜���f�V������gD��P'|
'm�9[�]%@��۪b>��hK�MW+y@�LV�"L&���l/?�IU�ܮ��L����9���X^IQ�,���.�L1��{���kmf?�XJ���:�_e.�o2��f;s����,u���哊�d�7u d���2l�*��;⹂�gC�N�݃j0P~�����J���\��ȩq���SKUu��z�/��Į?���	��%z�E�՗S�%���Ѝ~���/-d�R�a���ېG"�&xzާ�p��ؿ����U�f3�9����n{\�꽘��B`?�761l�>�Iڽ���G�YB����/keY!IE>����⭞�c�ƅ/VWk|��˥Y�o�dB����3�u������MP��36��B�~�<����쾵���H06�w^���,�VW����fhYߪxH� �>V��5%�)���|�"a��\�aݖ2� F���m�߂pM�r?؉1���h{����>�5;�y��Ⱥ'9l8E�"ژ,�L�v��и#�>Ub(�����<�� hh��~Ϝ+2��|+���2� Nv#��[�=h����x�~'3�_<ZƱ���GsQ�҃����z�Bۮ�����(g��QcTt'}(�:~!4l��5O�$߳�n���DH��W�TS��k:Z���`��wTƆ��"%f$ddY�.4�D����=+Ub�
c���K����@!\�H->� ��GK&ϔ]�WD��.�d�4W�����OL�Խv�(WT;iX 4��E��s�lv潛���<�ngpxDlC�".U��/���@�sN͔m��w�Zt:�W �I80�W�CD�ǳiH#����`o�N���"���3`�g������x]�y�:Al@G����,�ݡ��m
��h�Nb�X?_'�Dx������=��jC�~gSłdn��tp���U��8� C�b�GE��V�Zi4|��X"a�anRUh���8ˉD@0�v���#�بBXAny���"�����)o3�ez�:�Pz/�r/H�6�Qf���X�� /(���O`aY~uX8&��h�M����[�����iq��)�_S��\��輘�����G1�����Q��t��[�<kMN�� m%@z �?�)6[��M���F\7pMG���Lobxj��|�N�
�^~`��v�p{���Y�֊JY;y�T�c��mxy^C4�Fw�Wt�a��RȪ��;�eV���x|��t]��H�ٹm��9�.�ı�M:��o�|�m����3���n�b�CtV r>�Ӻ
�$~m���[���q9��g�g�nK�m�5h-�|V!g{r�C��k�cIx���S��{D��6�{��j��֞3�����ϙy�Pb0Ҝ҆�Z���y&�����;,���|ޫ��.X�M���xw�*�->7-k��=�,翴X���iZ5ӹQ�YT�����ǟ����10%�,X߽`��R�n$�C��>}Q�p��6�����J^޺�:��p���4�<�=��)3,�P���u�§�P�������*���]��:5�{���B��w{�� �G���-���	�7�������� �s'2f2�(u�+o,k��ɼ����p�ɳ��<���<��&��>8h)O��R���d��想�ZC �ZqЁ^7݅5�צ�dߏ%�[J�=���p�i�sR�e��k���Z+���0ooK��/)�y� �d�|'���-�E��,@��Kj��=k�� �_ �}QC������QX�g�����R�$��<�u��K�� �HBf 	-�d��e���y��9c��]2�h4$$Y�eێ'��¥�%���#b�%�C/�沈���s���=��dK�:��i�w�L8˿�31]��|�h��a��)�eM���0�u�!��!�޵��j��x��}p�ƣ����ag�A��ؤ�U������/ʥ0�,5.�9��,J��?f���b���'d0(A F�]��d�AY&�TPʔ6i��;�ݣ6?�W!��%A���/	�U)�Ј���᣶'���!.���cK�5��Y����ի�������ͨ?��v#����Ҟy�Un�+?28~I�NۓR,̠x������bx�l�㱸��������α�H�����$] AE�\�|>���>�N����I�S o�z�|���HCKW����h�V��h�&�,��������:���;݁�2�+��aG�ܕm���]Ie%��'Lp���;[�T��{�(߇�"�S��ET�C�S%l�b���g'S���JKR�>�=dFz��%B���2u�}V7���B2�]h::P4��'��?@��L����G2��ta���*1ͯǺL锻q	N��k�6A�!�o��vVZC���E2�gn>�Hwr��~:�ն��1�t)��F?`C�vl��v��{ �0Uqz}��@ٕ7檓�e�m�n�s�p�&�u��^f�@����i2y:�EBj)��6�\�5�����a�g��sI<����!pց�U�s^	%7�]NWʥ�z���Q�������2È�3�	������e��j�M|���x@s#�`:�7P%����ض��*��������2>_	��k��-�ܽ,&"����r�i�X���y�!�I�J����HՓ����W1]�&j���n��6ⷔd�/�>��p�p�����!�/�8��X���mD�t���w��<!�w/"����
�i�`%Vwz�����o�����Wx�����2��~�/!���A2�/E�O����>���p ��&^K�đ�>J	�h��fh?��!�71=h�ڥ�:Ɨ��#@���1��
vU�P��)ۂ�0$l��QK�J3J@(|�*9["�$��"��?@�( �_���O{3�N~p�3	���W�;܂������˥��O�zXU���̸6����n13������}j�ʚt�o�-
Vۚ�c�:�ϝ����WW3
1Hx���Qoz���Y"LEň�%��+�|=D���w��	�o�J1B_smM���t�)�U՜��)U^Э."��X��R��lV�<�qw7�#����_����{�m�m��mvMr�b�՗��K�����m�b��ɧ�F/RHF���<��������ى&:}���^W���q��� ���/H��ա!I���-$�u�W�mF��R)�7���%�d�mR	�O��@��xĸkݮ$3UNg+��s늷�6o�ѝ��]���Xh�"��e��g�tů(ۧܡ����_�X�Ѱ;�fN�~@��'��⡰�jN��W�&wT�+!�d�od<�˼�E<m��ڀ�y34����"��Q�'Ȼ|�����P#+f�x#è΂�g`i�6|P�	EW��ƞ͆���j��S.b�^X�r|Y���Y�A��U�UXT�\0���nVڨ�Γ���s�FE��F�,��Q��c<C�h�qӱ	�Aݞ���p/��1>A����j�Gb�����_�*���O���]�!E��.y�@���"�j	9FWb��PE���e���j:��@K�L`oJk@���=���QLp�����b?t��*���^�$-�{��_VP���;O��k�z�T�ܦ���Т����٢�N��}�a��4��NX^<�؞�/�mb����̮��s�����#	 ��=v1H���˼Q�0
�!�>SZ���(��̼ �6E�H���lZM\u��#��\�3,���N��s��i�v��9`v?6P�����uQ�%Y�����2��p�
|�Y)�����K�o;X��iі%�&�1vL~ұ(��uZj�H��F$U��b*�Z﫢j^Z�EƷ{?�Glш�SAQ翃���8�(g��Z��q4�%��"Hl��V) 1a:"я��(����H��Q*̄`(�/h��<%B��#�L�s��n�@��@A-�nwmV�߽i����{�=a"W5*\���eM!7_�D6$<�ɶ�C�+��׿�΅��94l�%h$������_z��S��86M����q|�B�	��[���/����Q&4*���jK�i_���(U<����ߩ���֔nW8��Z��s�VF�������W�<�����3ŦQ�;P�Hy�F?��.�P=U̶A]v��C�f������������DB'&,p/m�mϹ����}:��+��
tCXP�Y|��~dH���������C��{�4���9���&�x�EN"Au�*������(�A&���G<��{[ݙx}a�5'���"+���u ���V$�7� ��ߥ/qZ�M3 ��~��E��!;�J6s�w���� � b����͢"�}�N:ӑG-o�L���v���[������IWC&�v:�0մ��߱&�� ��H�VR�߻�+��c�p9�� h���H!8���>��0e��k��Jt���G���F�Xt�C+�� ����D��p"�wq�)=�ҩ�}����L7�s���/��ՍT*�־Xa�JA#�y�wAm[�n��v�ժ[ �t���sT�N݈��)��5$��\��{8)d轝��zJ��ڵ=�&N�a�%4��96���n0ޜ~W1[L �������yH`Mյ]e�����Iq��v�������G?M�]�$�슺Pƍq��lT����,�s�B�ᓄ�Q�הف������-�v?^'�󋷶��jy�h���4Z~ȜPk�b��}�PzJ/k�ZvN�k���h#[�J���|CUL�@�h9f^�7*����F���ԙ#\[��zYjNT=n�1��i���z�����Ɠ^a�2�#E�V����3|4�xZ��Jb�0A*��=[��Bй���+�Yz�'�cCj�A֍ok�����>�`A��"6���K�$��/���hb�+����i��ܱI>�ıV���2^��$
�=]bEj9����w��NlEˋ��� ay�E
_�5@ìE�P|r��8O{���{��H��
x���RsR.��T�����	�K�k�ؗ�$�j̓@�����2�լ>���x�V2������hJ�B-��<#Q`��>|���X��(��l1I�Z�@f����!)���笉��ނ���.m�u*S�6(����git��j�l�r�2����b��9��=0m�+델v0�����<�y@�\smcw?+�J����J=t
d��h1+�e�C���K��e���qɖ�0�b�=?��՞�<�>�A-����h������&*!#Q�ԥ����ٝj4��1@���gs��H��[�����a��[f�/�*���$��'��~�+4��q�#�ҁ�,Ԣ� c�{'`j��io�b��PbS��'xH�W>���дX��\��+S�"(���=���MR�C�kB(�����uɨ`�c���e�+<�L"k )a�Ψ���[{	�0��S;�<�D+��L�������>Ỽ]R�;��H3�S*W>��TI�]�Bؕ��~�:oaW���.(q_W�= ��]깞rA��\9(k,\�6�u��azy	!f! ��Д��FB	���צ�j�E�Rz�
����`��>g�/8>«�s��~!��{��
52p�|��f��q ;�4�ߎ����Ҟ>�c�=�aO�@�|�����Psx�Y���Dٔ���U�n�E�Hc}y���M����'*�w���M��i#�{x�������t^\���N."�~-����a��ӻ�q��DR���^�AB;�^�J��泍��!��(a���y�||����,�,�������#��[�O@��^e�˙�}���cj�[�[��PJ�gfj�@i���YM4����]���aޏ��tőy�����ʹ�\�u�����a'��x�L��&U	��'`�X��Z~-���uc���nI�3U�	��7ݹO-͌��(��p8F	��G.�M"���4;���1��4�Nc� �:T�-���uH��01Q����G�g����7;'��P+��.b/��ze������.�?��O
�W4��K�-�Ι0�̺_���%�3�l~��o�y�Y��3�&���b�%$��\�(�F	7�Wv+�
OpMc�L[� 7 ��2�<f������O�l��ە�C<)k:ـ�Uɣ��\C�T� m�s2~z�Mqϓ��,�^ st��E������*h>�`��U}���P~�*�}���^�*��[�z��V�`�F�$�B�7�ʫV�2y�ȑ�,{��*�&T�lW �z
Q?���������gU�~��Q9�NE���Y��~�k/���d�"��Ҟ
�a4���o�_yjp���K{ ���(ܭf~V���4�����Z��[�8����m'��-@�g6E�j�<�~$|# 7nP������U���I?˹�|j>5܅��Ȟ��ɮ0?���Z�N��lfb���������Ȱ�^���BG�ؖ�F��;����E���|	/�8������Jr��ْ��ɽTi	�CԖ�:`P0��˸��U1ŞvWM�!v�����x��48��G��箨�)hn^�e%�1�E���E�Ǝc�f^��(��� �����ԅb]��M�?� �U7vj���b�MP�1򿲑��­����w��h^>{~C�g�Q_l�@o��u��[��f*�j�M�F�yvƜ�L�:D�g��h�O(��|�æZJ�АX���&ܩ��^pw��=�'��������Nb�c�D�k�b�⩂aj|-=��6S�Ġ�[���H�@�vu�C�����K�J��k(M^v,���-�<b{WYB����V������'8 ���)�*�[<x��H�/��b��^My:�\���Q�I���TD�,x"�1�ڠ���ʎ7��2����C��H��Jn�!Փ/m�X�����:;wz�\���W�ѫj�Ҹ8N�O�k	��.���Jyͯ.�������&�b������"�F�w��j�	O�`66��:�P�㻲��.o	�J�G��~��*�L�9U]X�I``8�[��)��~a�s�=i�t�����\h5��E���z!aJ�+N������T0,|�|��������1�L�)�	I����Ř��K���A3刳��������͆�a���׈N�f��@�[�t�R��w�A��zC�L�R�(��'By:�r��"�%{/�n�����5�g6fV���p���0���Ɲl��˿��bV�q#�l�%*�vϼ4\�U�'����h��:���W%�}�9����|�2	�m�w-B��g Hς1��:%˚5 �n����3��(�S�Yjb���gs0��j�2Y��j�F��fe�\�~~�FE��B���-jH	ҵ�!�:Sޥ��� VrB�:X�q�ƥ� $�#t�?�U��8��O5Q��|�%W<k���ZQwN;	���t@=�T�η�GǷ'�#�Q�]-���c�y�s�;V�!7��X~e�[ H2��z���VU��<�eJ��dw/�����Y[�a�Ȃ�j��on��u�j�G�I��$���@S�âB�>����U4�٧��rn��tԒ��?ۯ2S����]]�r`/w�ܠ2�j�^H℆���~|>���~=M�r o/�����^��/�:}.�������GR9:��M�3����) `��� �CJ��!�ܤ�^3� klU�m�����[�dx�^1a��������?2���[��@��Il�V5�Z�7�>���b�	�w��ľu�|�p涬倏�� >~\�-�(�M��M����9�ƈ�/���sI�9�j_���L��?Cr����/98���[�p�@t@��\:=�ԏ+���k��v �0���w�kea�.��Ek�9ӟT�q"�HQȥ`k9w ���Q��l�J�{@��)]{��M�r��E�o��5�nl#8�' ˡbR�{����˭��}���=���#��l�ݹ�9��REI-�\�q�`�P<�jˠƆ$�
�?�>X�
�2���2��?6Cǹ[�}���@AG�L1���z��)����I5��@_�L�L&]�,��O|�ht�%�-C��-�'=�~���s-d���Ȯ�.�s�4�S�A�P3s,��mրe�a9
���s�7�ɺ��Y	��<IE�c1ӓ��� ��Y�_��{:O�., UU��h�	����m0���u�rw9�>·�j���d��:>H+��K<��aW����C~����a,B��e����W�m �j	t��A���Ǻk=U�7��s�Ke\��Y���:�\�b2�B�[�R�����%{��˄�pU�7췉=��R�4L�gULEV�$�wA�x�z��u�q�]<Lp�񣳷��4�j��5����%���4�A:������6GW�03"C����p}AF����yS�R�~A�Ul\�F`g�#�v��^��D���Xm���w�.[��3J�I?��z�RR����}�?@�������.�]�D2�f��Z6���w�~��1��w1Rm�Y�oD���_Mt�)>b�����3��j�x��9�UX�e�h��%9�3�N��j��.�
��#^�o$3F5���:׈��x������"��}Pv3֜��3sP���G,��#�������&c�K��Q�,S;k�9���@��S뾳���>1�сՊ��B>ħ�&�1��ƅ��d;8r���0����+�>sVm|��%�_N��eg�Y���,"�̬��n������DB��F�e�P�����y��X�.y���L��:L�甛i��u���Dt�7�ґV�Ǉ2�_��-�A��ւ�F����TiiN>��zղ�U$I�\���u8C�і�+����[�v&_�ž_@��/�b���d�K	�-r%9�}.��C��[�f��MS��ԒZ�:�-0�����!������nS�.|�Q5���om��S�a�}��&8�&��9B�F]�D2��,IF=24�×�4��x?J0#QxS|]%��ߨg�B,i:�W�u��n�)��9�
�<��b�q�����/����[X�i��q�[��dK���%3u�� ���T
��g�wl��0葺��`�n��� K���= FB6<��>��D�֕Z �5v$[3�U�z2��r��=������C�A���4T�=������
��*�fz;���6�Ҙ�5��@V�1���֤�'��͜7J��2���Q:+amY���{,�'V̍�X��o��V�7}ľ�Z��2IQ������8�J��=}2}����E���@z�b���R�I�!�5����"���G���M�~���������ꇸ���h�i*�A�/�j�a_�/#4y�z)�l�#Gre���Z�dϯ��g��g�=k�8�Z�O9W�q�JR�Q�RNE\�BwÙ�y����]Εd�8�M}a���SZy�>�X���Vt 9٦���Yi�AĊ�l�n߷�{�ݤH��¤$��<�Z�Pe�|�l/����S�0�7o����yP&O}IN�9�!.f����)jseۗ� �b�
�C�m�1�L߁�(<���i2t���XW��&�ˌJn2c&�����s�Id��w�٩
Ԗd�e�ؗ\�y�I�e���ZV�`y�] "�J�r="�:�M�V��e�i����� �Y2�4V�E_W�O�'�����b}�/`����_�fJ���@��\�n��o����7����Ϛ�q_��`^, �ň�1O������f,g�|�T��H��d+��z��mxM�<G9$م�$v̮�v~-c����_�wĹ=Х��[ ]��J��)%�)���
������n�oG�pn�3Rv.��M��C��9� $^>z*j9���w&P�wEP٦J=� �z�;U}PAmD�7@�#%"����N$E�����I����c�ZY6�!y�����3
�=�#�����-�޹�Pbн��1�����r����<���]�r���kϘNM3���$~d%M��6�O2-E tL�	f�r�!��63�H�U2�\�qJ;��.��l���QՆ��b@�{7���i�d!��_z��dVS���W��AYt�X�	@�P'������3-�V�>2
�7��Dh���Ҙ)��Dn�X����ْ���ָ ]��˗���f X��˭X���n�G��iG�'��5�NG���;���&M��8�Z�s��?��/ɽ����� �M�������5r�O�>g����Q�E�Xa��z5I|�[�E�?~�����R@!�Hb}�����A�-��x,�K���rKGJ�K�u��=��LT�I��L�D	��LOc^f:(71�e��SAb�f�I/]��;^w� 5�U�U��>+�p������2�(��iyR�:�΁=��֑�"��R�<�n��Lr�؄u<(��:+b�L�>�Uf9�1��`��Jd�y�Y�z;^3�wX�6^��xwA|:vqG�����,w����K��<#m3l��m�ɄP/����������
�{�����߳C���,ߙ�;��:3_6�@%4��D������o	��[���Sȩ�U�X�IԇS�?i�&�!�z�����v���cjP�si�'X�h�Gz��S�d�����H�#�E>X����{��~�˹B�ov�ĩ��W�9kL����0�ڻ��ө+�I��J��g�M���2����x�G�N�����rG�8ֈ(�j���;���E�~.�Z��X�*D��~9���%�� Z9�����D ل���<�c����
(yg���́v��?g�9��W�g�Il;����]����%Ԧ���\�F�jV���bn!~��#���e��$��qc�6��(���� �WM	�"��Gـ�����F�>�������^�H�Ϊ�C{�q��\�c<�#x�>r�_���x���H29�p���7�΂��a{~���J�
���U�� -<�"�Ϯ��e͎הb����Մͩ�m�;-���?�L�\9�y�bfcT�f1:s���3jX	�1�����2�^��S����X#C��^Q��'����f
���)���~��;(=&��~?���ʦ�#}=ᙢ-�YOx����Ep�B��F�#y>�Зo��Qߠ���|�]q��O�ͽ㭝ɕNTzyJ����>=�Gȏ��+�8c��rv7
A���3����.#:���,�4����Ⰵ��A��*�!!����:�q���B�4��o����&��:lSW�y�!Y���Z]g�
��˼�3��C�	��L"*���U%\���o$���.��+1+��x��bd����D�8)6.�i�À���*/�[4�ä�Ds�0����J5�G����)��q���%�/J��If�ә�#Omf�(������vɃ�,�g{_��H�O��=��yH�q�R���bZOt�׌
4�����MR��v�?4[6�!aX�H����G�3��e˰"�f����{�ɞ���a��rQ:N����r��a.��|9���0��%-�U��5�($���]8��-
w#\��������A�A���Y���F߇TM�h�^[Y��b�62����ҟ'��|�I�H�UO �]�����o�EX:�9CqI�⃽��������އ��M�2%$�e9h!�;.���O�����j��p�'d�I-d�)$>���_�)?f��q�(����C_�ȡ�	i�1#�a  ��(!�$���k5���~���̃;��؊
��jh%D�����w?e1���PG��X#'�P�ψDI����/M�R�&U3b&��E���M'M���p3�ǋ��b���{����|jD+b�pp��q�K�|�ZX{��3���I^�}�n��1[��si��&I8_@��+0�-��g�:
�?�� ��А��6� �#[�`,Qщ^*3��;�3�kaV��x<�q��	��*j�p/�v+5{�m�������D�c��$91s�3�p}#q����P��7z�K��L�J��1䃹�Y�H��U�#]3��e�]��Ra�
ď�ώ�y�;&�`y���~o�\�+�Œ�bI���J�H�վ�5�Y���V��V�9t��r+�$��Q;�y�����" p�%�i�/�!����'ٺ����~�^W	{��V��\*c���u�L��K� ��sij��x�2'��CE��4���y�8Ҏ[�)��*�c\Mg���׫��䏿N�!(ie� �ۉd��y9�L�.����f.��2Om�6X��H_����A6,Z1���>�s�'Ũ������GޔgЄ�J"��ud]�	��M_D��͐�ɻ�ڲ,��q���P�C�.MN%;$C���D$��$t1j��l���2w�9|U6��'mHk
�s�4{��"fNI.�:�W*��G��р��î�E&�����酘�T)Ϻ�tV�Zʆ%� ��U&��A�<�wl��/�0�P�&?NǏ�Re�V�%�õ�0=hGG�M�\bҽ��%��5ݭOY��'��:m�aH���ݖ)vā��#7O����dU�qg�g�jj"5�kڡZe��.�m��.��8���mj!w�X�Q��`�O$��CǦ�c=u��gL])ਲ਼�:d2�F˛P������qˑ��'KZ~���] :����-�Hha*�J�m���J;Y�i&V��<�D��>-���;�i��� �x>@&��3A���Q�/�缮޽� ӂW�%���ɒ��]���) �tT�f��������$��j��MZ"�̢� L�k��]���m;';4!���M��I5�h"oj��ܯ��.���'�N�V��uT^@��!�P���٪z�Mw�W��3-�l��VO���=�Q/�g��TH�/
c�R�F�I�2�j�P���Cٳ�k�P��V�].a����B�~
�%�jP7�B_82�����_"�MSn)��S8��+�?V�*�V_G���y3�o��+�wx����;�J�q�d��^R��%��b�����M��y-�^�-Ɵ
��M����Z��V���n����e�@_��n�����b��[��Ԫ[2W eMЦ}Y%�=__�-�}�W|�=0�?���=�U�8w�ފsmH���LӦ���q }׌��Q��.R��	��L�q޵�0R-��Zlm�ӊ������CW�[�"��"��%��ĭ9����l��?bU�����Ec���RE��z�4�������ޣ�1�O�6&���d&3�6�7r �rgy�m�Ý���񴪟s�?��pwrf��ᄥ�O��kj�o�����gp��stzkc���9�~���ަ��	�,d�GgM㓉j����3����d�(4��������lZ� D��ٍ��W��6yc�uE�'W�{���@6���pe�!���8 ���s�A 0K���x�H���/���h�v�/�����J�"���l9�]� �̏�'%�݅���������{Ҩ�w�)�3���uv�6bV�!��%�$���E17K�xXb�+�s���k\���4nQ �9n�ɴb�'J�A�a���]B�	��?p�r@�ی�,�	~���������fE(΁�����Ƽ����Kq��U���Z0���9t
-
�@*?����R�,��4�'�b��F)��,�'{fE����Pz�ѳ�dcN�%����M1$��sϱ���뗈AW�w;�0[���|~�>�G���":ʀ�F�T{�����)!�0�<�6�GnQ���IV�m%TX|��8P���h��n�w� ���� �Q%$��/�p�j�1��y֤U�:opمY�𱶹d�p �|m�ZT�
�U���+�[�жZ���d�s���:�9b^��uS����gɟe<�ʫ%�<����d(�͕#V��T���P�Se�֝�{����]�:2�<�떻�!,�
��ge�*���r�ܒ��؉z������㩠*��x�!�9�7���wd]O�:_7��䯒��	6�d
a�gg�7�e�b%��4�����WS�>+9�2Ԗ�v+F�$`�p�Ɠ�D�-�� ��,9�`m�YF�8�bS��2��L��I������h�n��w{� �L�d	�X�Վ/�*<�zS�SXr�w����X4q��YG��z�C�ʃF�{��7+�Q��[���N/B9=��V'�wbF^��dV�'8T�4M�L&�U���Ց�	��=r��H���(#xD��ʚ��x����cĽ��I��9f���nW�e���:���D傈x�s
fn9ϐpL�Ȍ���}�����?K5� �ڣxD\C��w���j1�Va�0�Z�ޣ�I���K^r��<:���'��;'�s����3¾nZ�Wc\7��m���F`��'?����w���Ak{}�����*%��\� ����ʀuD�|]�j�څ���֝��'}�7���^�<M��#s��)!51���yɇsh2��>�E��$3Hܯ1�mw�F%�N�g��ߙFG2h;�<������$���a�����<6����Z	7_���	�GE�U�u]�F�+��)��s�����Y.G�`�ߜ ���uM������T-J�D\����ꠓ�}�V�D���!����QX��I��	�|���N���V��A�$�~��9���i	 9hF���sO�G��<��@�6h3�ŗ̼�ΖJ0�^eb����Z��kk`��^)2��^#8�#�M��R5s�j,�Jz9��ZZ�߫������ڵ5�D���;�	=m����֏UYys_��L)�j�m艞6��m�i ����W���p�֧�0қ�1۾�iw�8+4Ef�7(���CRR�����02�Q&Tt��LMe��� *&:9;mӟ��Je}�7���F�@~�7���P5�wX�]��ee����#إW���axs���0<u_��2w��B;�����O��w_����Sj���|"8�����Q?�Xw��,��~�׽�Z�Wg��^�6�`_�̠[�����T o`J����F�a)�h�����vN�-�!�^��g�N>��i�e���e��m���
^�v��Ho:I��6�KT񵍧�����|�R�� |<���w�8��p����qf�&�����e
��Y�{(�xvƃ1Ϣ��+�˔f�J����=a�\0�orHIM[Eh�X(L���Y�n��]�W+�F�h�B�M���r��$Uݟ�g�1/�C��U�9�A��X�@.��=���I{�A�[A��f�pNϸ�(����t�[�����/-:�U���o�)�M�^p������JO�qV� HJ�|����A�����"��%?��$X�ǯL�*3Y�w�ذ���4�8����~{z:<�;�8�;��V�"
�JKӸPjm]Z�nqm��D�u2����r���>=�D�˩�G� ��(z�e�l�aX�w�d^�� $Ԣ�('��0l��'a���p;�#��]��6.QP����n۩su���!�O�g{P�?٤�}G<���[�`y8\�L���?����'�m>��)�k9.���i�i��Y%����K ���:� ߮r�N9� ��_��a�L_����h��{=C��;�A�|�z��P3�i5+����<d�9��78�ƃcq��'���dMD��xB;����I�+�=/Z��M��2��vt<y����R� 9�0�