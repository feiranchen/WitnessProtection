��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[����%��B�P�O� ʁtA�B(f,�yk�0�l��ؙ��'�|�я��vsZw�%���9wU �����9��v!;>i�������,��PY�C�j��\�w� �
_��]w{����ӻ����0�9�CH'7����K�\��zӰE[�$�_t>�_�����T��]=ƍ��+�E�g�������[�ket���k(}Cm����G��Ǘ�}B�~E�)-OQ`� �i� ��Bצ������H��2�I�IL�ᇺI��JU�����(�Pk}4��v����ذk��@�=�	F�v.屌�Z1��$�X��\�W�П���3A*�텈o�zg����� 
��T1���fh]��������:o�zT�ښ��D12�Su9���T~.Y<f��(�-/-}\;�j'����c�/?9�9�#�b���'���B��y��6#@�>�mkk;m�F�׈DD�mF��z6U�)����^��x �����Ԭ�V;=��u5�>^�=YsS��o[>5B���y���LMީ�s�[� ���trȿ��r@� ��0{	P�W ��^jj���g@�fF�X��B:�'Q�q��(��KU<�[K�/T���1����β]�)�bom�@���`n2*�����)&��<��&�1�@�5]���9�ucVx����d��^�R��)�}��߾�~%z���G�b��)���}��4�MQ�yi"j&;��n`�h��K�Q�K�A�Ư���q���q�Ht�e�F��f.i�U�����\�6�8��ala6�Ծ�V.	&�琀_3Z��y^~ɕ�
]癘�[��!V�lf\�Aj~My,�^v�u�� LH�r��ꠎ_�_��f�*���nu�� �Cq`['(ƻ�(a����B��k;���f��`�%I�>\�a��xM���{1��2���*PRC��<7`;�{_�����r�4Z�nI��[����y�X��I��:�F�
�_&J�|p]�c�`<F�oOϔV��Ν��B�t��l�����7}-����&��Q�X[b��/�y6�S�Dc@�������6a�H����$H��Lf��	�1�]� }�����u{��kɅ�bTǑA�Q�j���8�d�]H��L�U!�ތ��m�(}��Qwy)�O�x���ynY�|+�.E?B�2�M8�s���ؐ�<�c��z��e�H�@;�{�㤟�v��ܧ�a��2<�N���⟊���'�L8e��	�υ\υ8��I��#�KJ�1Ϡ/�r6w�p�������Y�A����Vu�~k^�?!�Y���g��h��j��;@Y� �����R^�dJ�+l���ר��/	�p~�Ͷ�}n߽3�a��ap �%>��&|�8���c�݆�φ�.�E&#H�?*OS�� s�}_Y�t��x"�������̗���CRr�Xq��7S��7�2�b��d�e,BƖ�/�k�D������?�������n���Ju���ޓ�Na�Y���;����n�ۇI����x�L��|��W��V��jn���.��{���<p��K�n=�5j���rH[�gѮ�"����-2'Nj�(-�,0��&lY$�!	jI�y�i�B����9�MuE��o�P8�ʭ�0�(,�Y�э�*Λ�D1��΃Qb�x߳a���D�BF�Z~���"I
�s�Xs�%�����y���G |��{�<�����Ȕ�s�mo�d�z�A s�c���cm�Yτ��ӹKn���*`���������;KB�r��l��~�S�D��x͝�G�S`B�!��g��e�	�����]/~U�4C_����Y���-��/ɜ� 'v���3�^LLp�� G���C���e(�Zw����	������?�2����;P���n@7���$�F�I�}v'�<{ͣ5��-�e! �\
n/,W�ϧ�V!�p:s*g��g����)������b�f���z���+��< +�>����2�z��-�@���j	@���F���(�Yl�����םQ־��}-�O�Qq��l��~K#Hoʘ�����4����seVF� &;�������C��t�:]���92��%�N8����3�d�=G+�
s}�����/�d��e':	R6=��}2Z�H#sv���T{D�8���є�g�$3{��2ƴ{ݮ).,� �"P�jj�#e�aiƟ:�1��<2��IwM'����~sy�J$M�I>�/*�ϼ�\��D|������ع�A�@Xُ�$/5���FVA�[� �x$=��a�'W�?_v]�@����5��A��}d.с!�k��3���y� B�����PZ�W�	,p��J���ԣQ�u���gd�s�;�1��]Z�ґ���:�|-���`���mS�_`��E-�ċ�ZD���J���1D%̛9l���*�;�2�l�JLk���@�J�>�|ɪ���k�)7_��Ⱍ���D�]+ȏ�'����F�>���� �0X�O�k��u��p!^^���]�N����d��cg>��0�8��F������-�D��¬����p.�]�
,����l�#Tz�l�W:��ݦ篠*����U�{̇�N��L&���di������5܈�f�ȕ���.u�:|��4ꦄ�kǔfx|>���w&��N��U�"K�͚�<��26%b�̂�F���R��8�~[��!'U\�P"�Mo��n�11��G1? ��u�>2��R?$�<��~��/���gz}�23�{�){���q�@N=rp���݌-�&� ���p?fj��9�N��Gq��r�=)�����;�K @5b-P��"�Jv{�-��;���,��ٲb���IB6#>�+$�I �X�ۜg]��v҄:DUC?��#�st�>�>�0�v����Hh��[3s�X�	��)���K�/��E9�Y�B��Ⱥ�-��<@�r/Fmᥭb�xpv��Ww+_�+ǍXr��=��B��xZ��Epj���o*[=��)�J:B�w [���s��~�Z��U�W{E7'	�]��}��[Gh�x�g�?�H��(�0#Vۧ��z�3O�p@O��L�Ά�)f��[�O�BF��v�����'��g�Mh�H������6��eҷc�Dn��8c��຺��"׎e�eea�0�B����[`f����f*87U�K���2) �I���������B ��!O��+�z�?%Tԏ�5��*O�x��j�F׶�PW�ž�.E3��Xh�>[.��d��7Y�B�Z����V�6�����Fm�[J� @�;�۸�/"�9(��k���/�X(��\o�<v�t�OyTJ�T��5�0L\�%���BҔ�y��D=��H�c�9o!�t�������d@L0�M��D&�z����z}�}}��~�f�96�	H}�o�h��a��%�`�@t94508�JS�!F4�3_�%���B�i�[¼�8;h,>o���|`�mW�Yu^J4V�p���]���蕺������4���j��)�q#���,�,�0�7�>�����pAK�A��F�^�P�}�� 3�� j�.�т��/�d�m��nI���?F��dj�Dǐ���*,�s�f�U4���y֍r5���l��R���8|� ?)O�씮k�:�~���b��.�(���I��5lw-93��
	6y���a�	*P����3�X��c��g`ye$"���WP2Rv��T���Fʓ!��@.>Ƚ��s�m��n����>��j�t��J�=/]?��2M���6�6������Q�U�F�w�DT��;}�ӓmQ�!�.-l.��&�gv��'3��46��`УF%���D��7�zRѓ�I�TTI�lh�-����"�(b�$��Yt�vR�̲>s��)I�}^c\y|`�e���;L2�*Q�$3s���sbД^oHGx@ݺ]�ԙ��g��. KM��(S��nw�ɋ����Cm��4�fۛ��'J�{�
�D�!�l!����úCm���4�!����? �	�v�Ӿ����[�bJj�8⃶��XRp�6���K}�Q��<�"�܀^�Z �N��u��V"Zs�������Τ�td�}	_����s蜷���K��=IE<d�4�ls��B��2�r0���E�d��]�3�ms��������u�����*}�(0-��
�>�=�o6chcu�n��Q�	���ܜb^�9�#���!���lP�a��6w/Z�P��A�v�b�<�H�9WW��	�AH�Ap��r��f��ޮ�y���άA�ݚT �bԞ�R[���Z��]�Xn8����[��熎����Vr���nT�ві?BuB�svg:�E�=�"m)"�!��u�7��M$P8���1�HU<h�ڭ:�$<�v�L�4%t�D5E��sȜ@���y���
��`8�sJr�Z���J�w �Bhb��ۅG���%�K��.:.�p��i�v/��a����"c�IsH�H��u5��B��޳`��7;R�r����=�:1s���EVa؉�/��4(hRVZβ
\�������'�Ɨ�˵K#�p�Z'�^��+����EZ|�ڎ���9]�@M)2ҟ��;W3�cF�*s�T���y;�p�9�&��Fv�@k��2f2��'M�ae���{�+ғ��ek޴�}�6���r����?-��_
��V*��v�ZL��"|���HG�~�X�G_�͡���+�K5;���8$I���x�ui�冁�ݛ���G���6��֑����YU7>���}V1\V%,�̕x���������K��?~y��2!��~i��Q�r����PP�d6��J���'���9f�u�ʺa�z�#Y��d({�=�ƣb�����{]�_�����/�c�L(p�?��d6���a��jK�3��O��]�?''-k^�7H:�q�4�r�v4m��:�zp�]h�#l�ÐY[��ek��^����^,L��T܂GI5f��l��v�0�S���h��=���+�L5V�'H�.X<t�m���dJ�7>/��,�%]�.W�fcϯ[:�D��vT�����@���8V�=����u��Q��]1��8�����I��]Ǐ"�#_���k��� ����^A���|n�n�Ⱦ��N8�<Y#�@�������"8AkC�*ȉ����BA�� 6������1�1�p_꯷Cd�e�' <�*��[�yჲ�صp�w�9��DZ���-:lo�V��0d���8��[���1����2ͅ���ł�]Go��я{ڮ$[����M�����&�D�����K�Q�R� ���o�;v(a���,�����u�pI34U9ْ@����JP�����U�������v-Z9������1{+�%���W�FJ�������I�Bo5a��4SH�V���z�B�7���&�Wu�U�j"�f��˯n��9��	���t%1~C6�7u �(a�>�:��u��V���V��̱�~-����:�cj�e󜬐K�-�Wʲ��8�]���d�A2BW���=	�a&ǉ�H�Y}.�1G������V��������Ф��(s,<���%AL�ynQ8I�/��Q�%��+|D(�Ge7p���gqA�R��J�~��e:{f������B!Du��;��^1C�ќ�_�+���Q�h��b��y-�IJԻ�"���5��ffq�����%}n�o��?w��pI�.����0�l����m4�ׯ�������a�%�ʂ�
�*C�R��`�N�"|yd3�*d����5j�
��9Q���AV% �{��&Fc���L�r;˅�!�6���'��t!��LN�'�U��e�E�y���`p���UO&;��3L~N�t�'v�S�V໳�����IĢ6��Ѱv�~�~\j̣n:�� ��!�t�Dm���a�B�Ҟc�۸Ż%�Efej�1�����7�x
��4eF�߱_l�����(�	:�-q0�Z�Զ�qY�-�[�/ǻE����u=�[��a�t��+�R�Ou)Վ8�<�޶���#▊"=�my\������I�#if���r�Y��q<���-m���(��L��ߺ�W7����<�DsAݔ�
I�і�r�"/�5 .���[��I��=m�D��[��
띟�ΏR= +�/���7�ҒP���uф�9T<le�}�zڴk�F�pk�g�3��Ij��� �%�����8"mu*'nv���ȗc\x�,3��1�s���|�H���f_���E�<WXNݮ]<�4�in�$�y)1��?eI�t�pݒЏJ��"U4�[�i�6ݘ���-��4
��[�h5 c�4����{�jq��+[y�c�4͛mU�X՚x�Φ��t� ��iI� ���T�D;��=�?ݮ�>��1��,!<h���/�lWwX9G�\M��r�f	�2��\>'s'-pY���ě�1��[�-��X�����yǐr׬�=�K�~���}]#cI�1��`���'Ѣ](��
��4)>����൳��V-,���Z��Ç?�S���6� �����l>�	;E�T�S�X�{����9ɏ:SΈ��D��it.�L��G����d���*!���WP����#����Ov~�2����U���K�;^� 7'-f�~�G_�q�m�ٰK��f�i�:�"����� �1�C���Yًn:亀�c��2�NhI;=� B+Đ@���Y�oN.LS�f�W���.߰�����d�L$d���uϑ���y�/r��F��A�Z[�!���JF2q��~1U�'CQ�����I|����?bmꅠ��h@�k��/�ְ	qђY��u{%�Ɓ|���t�mB�'����"��1�2_ۛlU��D#C`�֩�f��M�8p)��{칦��!�ʋ�����Ӵ�����Mu���3�3���a����b��~�}��Ӥ�Q��1��6�.�8�;C7�$�4���\j5t8foɠ�G�c]�ws���O�k��4��I�P!(���0K1�G:�� �����nk@�<$0'_/�x,m��/��/ �(�����>:P��=TzfH�o��!�ǲA�!�`�q����[05sh�c/	���)��9Aa�Ӭ�5kw�hZ��/���׹��S^U?�R��:r�1�q��_��UF�cE���ז"QY'i�rEu�YDFo��#?����ԕ�b���'vf��7oY�7@����0�h���&0��w#m17���Y��M�
j�����5���a�<B���Eh9[4�v�['�A<TҴ�q����.4��ō��!6K�'u�}$��a(�NĐ��K��v�����o`�'`b��3�ˠ��p�B`�����*J~�	�̀e#�~܃��9�k�ԑ���]l���aţ��04�'
`+\r����Jv��?�*ͮ�Q���;��=7��:%�Ŭ�@a �nfu>��MAuT����U�_�1�S�xc� �Ջ7�VrX��4:I�'���YC>��W�$��4�&u?��ڹg�]�]���9�x�c�͡�`�b��W�Ng�מ3���8�c���TM�����H�a���J��a��H���3�"+��Lt�}��nSƤ��5��P���VA.&���A���]�X��(5z:�d~rLnHؕS$�M�o��&�(�By�f�)GQ�'X���r��TB?�P�G7��t����w)z�#�i���C�O�]�侷��uۜk���, �b��P��X���=�0'��Zi���t5�3:;O]���B�)Ď�-���܃��K8?_BY��������)ԋ�>�d��L̇�����s>ǧ�4�Z��d5��`��Փ���4x�=�.%�ڋglZ���0p w����xA�����	畝}�LYjK�9
�EI�5:�F,F�&Q�4o��x{�Q#	��ԏg ����G��l��MU�D7�N���=2��K�zOW��V��[T��&�U �)�[bYg4mT��|�Kޥ]������^hEC���nR�Ͻ�孒m@��S@��YJ�Y��z	!���U�r���#�m��2'L��CA�u�t�9������w�ww�j�	u��J��] �E�z�X^G��Y
$��h>� 0JL*�vm@��E�-s��04��CK��>(G��S��}X�KoH����,u)�Q�{��ψe�@��k��T��~�
{/�:rW��Dܒ�gwj��h�>;�K��kv����(�ڶ`��8��`�]V>$���V���s���J3��G��t�ɏ�4��a��w���}a���$�8�4v5�Z߮���/���D��&� JCi�o!e,�c������Xu!*8a��(��B��u���:��#�S�!q�?�N��#��ءE魂����A2`;v�Cd����e��1���	8K>Z:�:I���	�a!���(!2Μ�1#�5���{�G�}�xcĳf��p�j�uURU.F��k���i��������E��i{r"n��"t+1�.��w���s�qZ�Z\!��&"�R��|��?�dC�}0�o/4����k@�+q��9�����)��P�I�I�'fe�3����*Ї5����1�ݲjF8L�X����o����&''��ض�C-*���؋�A�|�A��&�D.�U���� 7^�/K�b�.E�mL��g �꺁:�Mu� �Lu$=� Q8N6bPi�aז^Y���󶟽�yqLk�Y����չ���锿>tU_,�ZjB�@S2�Z�SPLu�ݦ�؁�elǾ�;�8�J���n���s���T�<W�DmAxC\�e3_-QA��7���5�wI�1åw�Ӹ�'!릦t(3Q��zR^�d!��C�q����J1]kJ�K�VV͟mi��^z9���dY�/<ڇ@�~˃���R�ţ&z�����t~ﳗ�l���p2�x����A�`�L+�1>tU�&�gx�����Z��"�Z��5�y�BA�;����C���ӧ���>u�������A?��9��%���Qٹ膈�U�ܬ3�R��?XH�ӊBj��A�	���\�ʩZ��봢���Ŵ3���HF�b�ջ�h}��ҥ�Q�������M~~u��A�7x-�����)��0��ͬ�hD.�\�쩳6��A7X��W;���P��N��fXۓ�w�'��Oy�6����ݽԀk��8�������� �]|���J�׳|1�DT�z�����/�|HgT,k���(4hx���6��!Md�Y�O�&���zp�]��0j<K�&z��}��(��jG�K8�H^�}��lc�9c�Jx��%K��i�^�5T El���ʼ�����\zp!�3��kȥ'd��e���4�`�XIb�0G�`��Ќ����/����><�jIv�N��an�B���p�Kޓ� �B*刃��yєH'2��>o�
s�"l��Q���G���H��	O��:cT�	�#m���0tA��c$�20E z؂N�R"u9��&^C��O�垐�����	byO�+��@ɝ������%H��؄1���ɷY4�Ù�|��֮�C�O:�{}�eEo�
k��M�O�u[dM�Z���Q�k��O'KxO��+
I����D8�ɿ��eTd��1�O8�z��8���M� ��W�G��Z��Ga�{�5�;�m������A���D�&��].:�e�a��wRC%o��a�F��[q�������+�R�l.&;�f Hct�z�%1����R6���7��`��']��W�'#҈�����f�e��")���<M�����Fn�V�.�Ny5M	�x��VV��З�2!�^2�ɭ<�`@L�6��^x�}B���H$,JX��k;�ҿy,cc�X�Qhɴ�1���K_n�D�r�q_B)b���;_ڇ+��z�|K�L�����I�]��1Ǽvɇ���5��VNUFH�1񿅦�y���oX�p����  �8�1����t( ��)ZR��r+zk�%�דr�=��l�n&���	��o���0(C.����JLS��O�6��GǏ����(�C8ब(}�;6ͻ'�C(���G?Ii'���b��u�	�tᖺ�[�V�I�IeN�jE�3�i)�l�Jl_��q�d���A�8��+Ji�@2�c*'0��0�ҿ���AQh�k��N�;B�D5���|�q<A�M���ǘҋw�n�4S�l�&"�Vm7��.L��!#/���������5�}����G�m&w�#p���~�(6`���c�Z�� X	XOQ�}�Р�1����"�������M"�#(�T�� ��c��y I��΄�R��NW�Q�x�U�x�E�}��y��v\0�2=5��6ŧ�h;*R�g$��+(�_}�n�_��6m�m���en���A\�7�(դO�ﮥ(˷����@��T���m���$�4�L�:��}$�/\�*�) �z���:n���X����|5��|�ꄍ �V��5�ʥ{Y9%+�H�N�඿�x�s�y'��R�_y6}N��	})�	
�g	�A�zZ����ĉ� 뾹,׋\��%9����o
I�q�j��<�yJA�z6�qs��K�b��0��+pDa2�R6YAї���C��j�Y��d���(yt�5 ~���{������d��	Lp�öLg�WE,�6.JM<P�g��V*=D����0���W�G(�X���ӳ&I-�A�V&����e�w��ɑs�/?�h��#���I<5�Y�y�DlB�Q6QY�RZcpc�iN,�
 ݾ�pU��UkY'�ʊ�W����
�	�F�,T�2�T*��%B�
����pA�i3���1	c?R�5G;H)�XԤ/z�������6s?McL�O7�zZǐo�bEӴ�>`.�-�u�TU�,��p�%]mk��+k�j�XFyy��Hw���3]Y�٘����b�VG�Wu!d�
}��1��8�fT\S�V* �;a�g�:
H)/fY�����Ф��gX9�]=+Ɠiم�j@�� ����7$�ďv�N�Fw,34��\��ⶉ�CM��e���s�H�m/9K{�����bҎ�n�� �[��m�%�,�N�
�I4�l�ae8�H��H�E�]q��p6��e�z��$�_��o�rx�@v�?&=hM���-r��
H]��F]N��}L��o/��r��*������	z�0h���P�� @��F���
՚�t�F&��fɶi��Y��۟O�0��=|�dh6t(m��(�_�)Y�����"�"��, ��&�-��ʓјw�uU_
ȵ=��ݣ_F<��hh�~T(�CN��/�<_h`�# ���J���������NG��a�c��V���I���7�����>$�i�,~ih�|䫅���4�N��<�V�6���u!QT�f� ���F:C�T�&S9n���6n�٩�_~�x6ࢢ�]Vou�%�܁8����KQ�=���"�rb�uHƸF�w2�'I���i��m(>N$�$Y*D�Hk���@-S�A����2�_+���W�Kx�!��x*�c3��"����kQo.�t��Ea���{n���Cp�#{��ݛ�L��`V\(��B����:��\�����]��g�]�E�<��%=�j�}�z�����n��Y�b��3J`�(�̔�H�c�:�/U����#����d����3j��Ta�&�m�n� ���C�an���z���_��MGV�K~��Sc.��_�+L]p���=&��,0���5���C;�Q!�̋9�����'���`�y��`>l��!���$��h~�݅bf����ɰ�?��W�e�nm��rm�[�!%MJ�b]&#�s�7���VEJ�x�% ��m|$:��J���c��aV�ʫ��Nn ��F[f��F`VA���eV��7�0�1.�:��
�4�_��K����q���2N��h�d�es� ���U�. �n�"'XC�������\6�Ϸ|^@�N�)%�H�����.��tZ�2�s���$���K�h|�h�B��/^D�Oڱ�1.X�����`����2$��hy��9��#Iϭ�]�����8�2���9H���A���3��VL@���B���'��U�9��z�ka.�d�A8�������w0|&zĹo�(�X��}�n
��.�����~X��n#+M������(�H8z�UܢP7	ą\{"2�No�>ň=��d������������`�I�W�j}����Vd.� �m���7�w�ٶс�&JY�XϨ��~��¾��w:Ӳ�YT}�[��r1EEZ���.�g�%�������v�@Eo���{(�)�S��8q�sR(2ͮ�?[��.�%N�D�_���BwЊE����9	�F��;��Aq\���~x� ����|J�H���d�=5��ƃ?o˔�����:*�o�<0[=��4�O�3�,1����x�Vz��"P�o���곍Y�\n�
)��S�G�y_[xT�	,��l�Զ�m+-�*^%�@���F
�;�e��BpM�` ��� C?�����m �׌N�]q�oS}�d:J�L�#m,�L�C�IY6��WE�M~�5�3k��>aƘi�)s5�Ԭ��:�O�.<�x�9�k�D������&6:�x<�d��'N�fh�/�4\�g.�󇽗�_(�Xޱ��� {��A���3����;���q�sԈ��x
ZSc��v�����Wpܒl�����Ȩ&}���^��}(v�'`B���ex���~c�����;I���q�":����$�ܒnNt���(*{f��8êB�V�Y��k�u>�K߲G�N��v��:Z���@�C*K7+���}�.��؃j/�m��˄��ˢ��t�L��ϐ��D6�j�~���7q�L�]�H�l��n�]|��f?���7j-�o��Um�C�,β�����?3����v��Z9�˩8�4��`�q�!��@}��{U�R-����.rN�&��2�xQ�.of�������N���6R7ZP,f�R���-�]�Ӌ�fY�e+����Hbz��f��+P���ja ��Hg��u���b�*�	kkVP����7�7 �}�P��o�T����R:>]��C� �ݫ����ꭱ��ob��wk����5;�(@L[�O+���V�Rs���̦���&�>���8Y��`��q֫g6Z�2-��T�FR����宻��sټ0�s��ѕ�J2�U�)�����sjм�/AD�Ed�$Qm�E����q���:����{ c~|o����FM�:�����vo��q��:ߨ�u�JIm�Qe����l�Q��J�22���}�����}1'���4�S�-���m�J�P�Ƭ��s-�
H��&\�Ԫ@��HLk��Q��ľH3�jg1y/~�F.�D�fV���Q����K�Q�9��V�pF�S�� F
�9�����E�?D��(���q%���W�e<�kgWZ���S+:���CǦ���+��ڬ޷T.Y�Q���zp�k�����BVe�Đ�������b���o���=!����Ռż�uDY�"�8�.j���̷Uw�m,��x���@2��>+j��geC@X�%{B ��dM���3t��tj����ѣ�Q�<߰j�X��+1#����=ۈ�J��$�nA�8��_w�x�@T@U��k��ΰ;H�/v���������@���񧕼���L���U�Q����9>���X��[]�!H��)h¥!� �QHn�i���>/I3��� ?%�$Ot�D�gP-�ki:�  �NG�N"�" �@��0lhLb�eDMG�a�
��责�-�l��6-�&���)�>��v	�&�t����U6�^�3Ͷ��"3����,jC�����g����u����@ǁU����Zh�
 �u�t�ߣ�_,���Ѳ=+��eQ=>� ��h��u����X�Α�Ս<�8M���@o��7]vTy�X�f_��ĕ�d�nUj�r.l����zap8�n�7�5��?p��L�FE��}�[cB-������K�][�̅��=�
xT�/��k�S(�����G�@�	Q��0q�T��I�Wҷ�}Y�$��00{��'�˫^��e�(I%�:@���3bq�^�=�D���@��~��5��Z�˂J�P�<Ɲ�Su��f���:�~����5��U��Y���[�������Y��o���OAYJ��s~�_����3}J��C�#�\Q��#��6��Qe�cqc�o7"#r��$���S�<��ν>�˖�#6CbB�Y*4՗�\L��5B���4_Q�0._���ǉ#��d�W���ei��+��K����ך��0��7�c=iD�J)So{F��D���Y?[6�4z�A�0���������]˲���!D6\փ9>Y���٬�)jnp�=�c�oAiwBd2��v�M�\W�/���`� ������!�4�G�V��$$��.l�҅XX�L�%���Ǘ�L��Ez�C�#ؠ��}��9��Ԥ>fm~S�����* i&>2��UѦ%��s+m��x�0ȥ���Æ���7�x�5�]�/UT�I����FЗ\UC6�w2�+����\K�X���Bc�5�Y�5 kꍐ�'�ȅ���1��{���w�ЦN������P=��k䊭}-�C�����g�F,��p'^d}z���PMk��oD�F+�q��I�E�9�A�h���ժz(Ai�o��}V�y``iu'��e;�%�޲�hj�B���~}�Z_�:��҇%QaL�ͥ��[:���;�8��_m���.��e�μ�c�`%�&��2�k�-�<U�� ŕ��ժuߥx�1~�n����(��l?��P.�C*�T�h����yl�ļ�ʟ�O��r	k��X��R�DOi���*�F�`iQ.1Hԟ��vj�w�/�� �������'�xj�R���q���9�&K0����C��|��u4���t������o�Z�i#�n�:	;�jO/�ٵ�[��F�u�4e�@x����5"��e�p�ǅC2��<���i�U��Y
���@�`�zT/�܍���^uay`�H�u�f�QBA|�R!��KL2�c8�m���
��g`R��x�H,��������:�q���1E5��An�0�M}�vQ����߷7�וPr�U�1�c�Q�]��#�)�!Sdj�����آpׂ�'ĝK��$x��'��/��B=��U��\����+�9���=��H�SHZ�؉ƻ|��F�?ш��w��U-'J�Mz�u�DG6��=�gJSx<��!�dz���r(P���v/�[����(7Q�aϺ���y>6X ƗoóM^�������U���$*ib ����qt��L��x�/3��\�|�*AeV����1�g��{�,^�3.<��z����PͲ��Q,^F�z0�qZ��8�2AR����j��}Ә> .)�� "�3���7j{�W&lP�̲KR饕7;;�ovl�8�ΥO�w�p�m(��g_��zS�o��p��Ⱦɖ�V#B��}o��<���9��"}Kԡ�DN�˔w_q���c�p��Jx��w�~�$��wg����Ovk�w5�.�Bҧ�Y�vxiuB����#]�n(�`<�~�BA��]nާ��ܜu����_����JI1�տ ��
�P+�4�{ǁ-}���0���F.J��R�)���ģV��K,�z������&FM��a��$l�j������S�>� 1��x������� �Ǯ#��w��gL����N��l��Y��ћ���͹�"9�x�\�j)㌔-��N��-�rv�=�&�uk��^�G�<���JU��5ި�y�e�Qo�~I
�m�H(�ae��������O��U����_*?5�zF%��է��=��qoރR���N���Ji�S�m�-�C�{��N%���Y�"��=��� W�~FS�H�]����|O�?�MBq��+�c��hiH3P�핊����Jno��.�fv(�7!�]n&b:����a�J�UOy�� �)4+�ij�H��s2іc����a'Hܛ��4��,���z�]=.����GI���Y�2�V`����_wcˇ�Α�q��y0��x)�I�����K>�6�k,Y�}��er~޾�X8c�Pٍ:���Cq�n�H�>6?p��(�,���Ё_�'��z��~��St�.i/5K }��3�4�z�0��Rƚt5��@�N,�P��:~v�~��5�l��!0�h�ӎ��Z�43��U�����޾@!C���òU]�n�^ܣ��6���f�Q2��������9��w���>�gL��]TY��`� m.2�[F'��b��T�RX���:�����r?�<&O솣�~��������gy�jZq�kI3��y��.�x�聃
Ul��wu��;�(ǘ?�� eRL�/TI�Ϸ�٠##�}b{@���vHU�)����R:W�C�_�������i$ބ��=NJ�.)�O�	�&��ٲ��e�z�͸���������4��D��-�*+�3�}�E����W��pgC�Q�#���lv^N�7��ÌJ�G���p����M�1�<�*���0�Z��I���,���ݍ��a��P	�g���Lj@����@�z9g�{�� �5IC���� 6ࠕ�3��$��
���Me0����B(v ��NQ��H��?G�J���!))W�L�W �iG�����!FM
Df/-J�ae���%����R�A^��Y<�Ա8<�k�Gv�2AA.���A���^�T�M�G�\�z�pmjַp�� 5��cCA�.7mI�o�1�E�4��B��H��N��I	TO�;L}Z�E�KzF�őzm(�c��=��<�]����MmR�{��n�YOP�eI����Vw�	(��K߸s��oG>0��_:7\�w���hl��k����a�ac�Yn3a����c_�Q����[��G2��\�����q7�j�ti��G�轻�?���������[3���E$@�!C��n������L����y"�v��N�[_XdD�K��6�eB��cw��cn��ΐ�%݄�d�S�s����H�,]9d5��UG�_�}:
�LěD�=B!S
)��,�q��64�nB%<��+���-�Xx�Z}�넓!�����c=�B�DA��`l��K3�s<	~�Ma�X�`؊1���%��ApF��٭<��s�4�^�hX�<�i3��Ek�`GUYp��(|������tO��
-�Ư���~tc�O?S��s��%k9���c �,��@*|+���P�������u�]��wI(B��)�"	�:��?�O�6������kW�*'M�|�*)q����?K�������]f��4��6�iI��X]�f�4���\�]Z7Zм��1G�9b������.�X�2��D;�0��%����s܂�)����f� �e�D�* `���M��<;��S��)����?��`���L)��Ank���.l ̍]��e�d���1a(�O��P]����!GI�/�O��i�qN�3�;���fr�Ie�+ ��(�P���2k���N?C���㉢/���ME�6ɢc,;�]\��9�~����ُa�yw�H��q���g1J![��ٻ�ۖ�#���
M����	��H��֖��<a��������̬Qo�+>=D��{��^z������QUb��-|U���W�c�
2&��K�nc��n`{�+z{�J�&�E�r=3{��=1޿L�~8��l/崴Y~*�ћ�kt�Y����E`X�f���V�/o����H�U�8������lD�L�%�����
��̏�D$����+[�&j`�z,�A�k���j�O��Ќ�^�i�^���0h�^�Ċ�V�3�'b�V��x�(�OWڃ =�4p�t\h�ڗ�(� j5S� �Ozp���*Z�7�3�3�RWX������m�����H1V�_�S��3G;:ψ�1���|�CR7m��G���8���"�$�G.p�$�Q�.�y�#�M�h��L�C�f��w�<����ݰ~�	ci���Hxlh)4���Ea�zmu��S��2��7?�+߃t؊�
���lV�Z�d۪��jl�����)Ow�$�{=&���l
�+�YY`(�5l`\����]z�����n6�(�t	��#�Eq׵̆��ג�O����Ԯg�(1huY�_��B>|R�2�X�"�6h��e�8�=����dB�H��O%0����Š�87��{�eT���p���z����}`r�Ŗ�k���k\�d�֌��uj���v�K÷.,�$Zd��G�$�H�-���1��К�G����D�˴-��D�������z���`(��J�n��q�\7�GRiCtc�)����U8c�.���ҙ��Օ����[%�Q}�u���a���G�w��(�ш��H��$0���S�|J��7f=~8*.u� ������F�A�Q����G蕓��TEn��V6�<6fK�JX)٨fӠ�ԓ�h���u�xS�C5��)r�Jbrʪ�gv81Y�ș�Ͷ��o���i���g?D.m(�O�k�B�Ȣ���f�ަ���;�^'Z�ޘah��G�cZ�3�М�B�W�r�����m�|���e:�[�x���:&��}�� ��� �x�Df��s��3��~(r����⨰���W�+x�,�Ҽ�ag8ub��ali���USs+!C��s\����w�e|	�]/�@�6f2���ϧ��Y&��L�AY.�e]/�l�Х�{�a:�(���gٚ���*��	,ݟ����ÞhP���JŔ(}w��[O��&;ݸ�e�fo�̋~���s�D��L��׊�Fm��˨�dX���oʠ�6�O����D\�&
�_�K7>K��P��5󂪮�ԅ����L���u(w�w$�&F���{]�BT+�����d��7�( I^~@�!^����P����W��>�(�uű��厵J%GD�.�
)]�V��/!ܥ(�ȿ{]�
r;�Cl�TRJ�$g2k-�����u~�7NQ�O7�4��K�.f���5p<�|���fd;l�ae�yv�$
H���2�"	�dj�J������������cȥ�X�\�#0yT��b�S����U�("@y��G���p�R��<�5���(�~pS���&5 �zl`!���=v,�6�  �S�7���{����E)7���O��'`<+������4p��_���A��ԗ6�*m)+�Q����7ܛ8�67}ۙ�H,7�YcZ��mtٕ��w��,���e�ݸ�J��b�N�U�F4G"�����|�D��]i�H;��5MG�x~bm3"?�B�"��w�V�h,�8�}d�l�K�?N���J%r���x�;]l
&E@�0����m#��+e;��O�k��\"ԒTq��ahf�}cba��&���E��^\B����:O�9J&Em��|KF��cۖ��Ɓ���鉏��C� /={2��}�Gg�S0�M����8oʓ����9�˲/�>�*�?Z!��/�'vY)�!П�/BT��r����&tR�?X��\ OΙCz)[�%P�/�cT��sř��kx
 ִcn���8�5D�Q6���$j�e^,�;-J��F7U7b��_�q����;z:g����̼s�G�͂B5�+[m��y���V����Ժ��A1�h3�kF��͹��>�&�t-�]ul��az��sފ�K���3\���!�<Jrd��]�Ea����Off�/�I3����L��qɵ�&�#Y�ªd���?[O⒉֙Nע��e���c����ѷ�3M>�������~I�Ki��Cx�(�O>6dfDc��.}jL������@����X�A��F�-�bX��ru=G@��C?RV�v��9p(���X.�+�)mm�BD��*w�'��}c�|�7���R?w�Η�1�5.� ������MS��N�4�@�RT��R��Y'�o��X��
��o�D�z��O�]sM_u�L�f�����0� ɺ?�Bx/�Jj��;.��q�B�R��*
���,GY�W�T=�]�)�sz�A�����[�9?����[�~���:����s"1c*+Sy&h��|sR��$C����]W��,$��z�A�w{\Jw>�Q:b��t���w5{�+�/e��f8uK}o��'���5���V����Y36�UޜDc:i��8Z����Y?���P�˲H̉�X�?<����i�E�Fi �m"��sҥ��O�.�k�� �p��]E�vr����|ޝT>�-���!��M�S2�/�	l(0��y���>pe�Pw֯���`�@	h�r��ǿ�������l-}O���1��&b
:@���GAK�}���(������z0UjR�c��D�G���f�&3a�� }�<�e����+Ӛ_'M4V.�o�Q��!q���Z��v�p\b�w=�g�Cg�m�>���fŃ��Ͽ �q�2&b��mD�&�C��{��Z��/�C�AR��.+����z��6R%F����0&t����Η�8�)�m��;���|n��w�4�уO � ��,��#��V�3��4��Ko�<ġ��e�"Ҳ[$��x�G���HX�l!
UX�#���������z&���b��?t�W�.m����k��^4,�z5B������1�5�3pTRT;�4�zm$�7Y۬��X�{A<iQQx�vJ�y��``���誈1W�f��Ԏ<z#�m�sN�o��c�;�!c�����g�	-�B���_P/ѩ��*�O��.�9B\
���R-�����~�6�8���m�e����iZ&��C\!�#r�Ş��&�(��%y��xa�9K�K\;x>!����f�W�K���m�/�5��O[�&S�s�H99K�����T��e�5�|��Pn*��Y�E?\��iƍ54C��~@
�o�E+��}%��x	�*!3�Qr�5�'(�$�#wJl�R��M�2�v p6z8:,�I!�:��K�~b��#�v�@%�(�]�Ю����=�Y��G��]�o4�]�Ϟ�_ew}q��P��3I*��(R����Iԙ���e�.��%o���P��C�zBKL��ﷆWv��w((cdb�|��맊w�~M�0��3�i��_�=.��} ��W�=�y����ح{c�ur�Lf���uw����ߌ�GG<��E�;�r��%����C`�y��1r˥c�X��d�؈����'��Cq�zb��k�g'�"s �s.�r=	�m�������B����u�3Hv���X�>�x�o��]�������

0�.� G\ڔ���tT��³؆����ܖ��0W�s����*���m
j	�^8�{�**:�	Du���0/�[-��wE�b�k�J�7�B�<WKƒ~�y�hx�)�uV�Wh�A�1�����q��[^����~��\'��n7�f�۷W$H�̣x�d41���N��q�a����q�|�||/����я2 W�͆1�'ei3��S  EM��q�c���O�d-1b�#����O�Jmoh�;3h�ۼ����(�Z"Լ�M�.�~�*H��F��1��oM����0)w%?P��
�O��gp�E��:�x����D��v*���;�g#�N��P;*O%(�'�.�OQu�Z���̝�,�|���f��91�yF3f�*<�+x�JL�Plcgn���w���܎���FU����xp'M3��jS��q�RmY�C)�j��K�}�_���x��rʷ0
��uYM�@�fu� ���y��k=�Ӧ����_H�������*?;�K=�D���� ���oU�ϣ[�,T'��CA�&᷁��Δ�OT��.���L��ޤ.�&ҵiU/�!�ǌV��!��|S��nӬNXo���'�Vj��t���]c>Y��j����<%Ic+�7�!�[.�֡����y@�0֤��(?8aK�*y���J�>��:����vK�C8s����)��);'}�[����X��8���CRdP�>���ϩ<��(ЕcPE�Խ"��#n<�W�{�?�����P&Q:!2-,CA>����r��Dc	%���(/�X����o��Ci�ig`=/�`���DiՅe��8i���Y����tW�Vb�����7SgH2)׹˲�$�3q5M�����-��J����na"��r�E�l*=�_�=���n�� ����Y:�!n}��dυ���IXl�E�H����8si	��E�!t\`��@ �N�=B��3+Xh.��-/�}X�������~Ŝ⤪��U=�t�g,[d��ڐ�[�P��tWZ��!��H[�$p��q���t6k�ʟj����%0b]�����ȡ(Y�ĤE��l҄Ƹ�`�L�k���b�}?R�2�Y`�|)���Z��8��2~�o�8Q�Z |t϶z�~�����+D��b��\���5R��GZ���~G��[B�<^?� ]�M
v)V_x*@���u��S&3�W|}����%��|XH�)Ҋj��ɾK�>FL�5�B��Q	?t*�m:�����!O)b��`��q_��bKe��h����'�~���.�����_A�^1���+���·�k���ж���y�;S%k���m7�t�W���'?}y�6J{n�U�3L���l�K_�4=2��>��v�̏	gYUQ��~�~��#��?�@��?��ǀ���) 0�,�	��f��D���Y�5�vZyY����
ho\�(�m�����ħ���?ZX3�5�<6��]��gE�֒c�C�*����>ẙ�|=Gk��ئ��.)����9:'�I�ܚ �ߦ�T�:#"��G�RD"KQ�"j*��Tfj7������Ŧ ��-���S�Y-_�/:�=����Go���R�p�*�z�O�Q��` Q���w�7fX��7��"�h#�+I$������B|ץ!��&�ZJ^s���^)>>�s�3n��3B�DZQ�LA�=X}�Z~��l~�6���v�,�N��)L�Js��l��%Jk	c�D�NTY:L&͓��A�p���,�e�����[�4[���I��ĺ�Fj�R}�ڀ�d-��By���/�ڌ�X�:h�w|�f����c؅n���
�ω�*�Z̤���MY8O��%Qӗ%��9a���.I� ;p��&F+�>�L����Ԏ�v�?�=�L73c>���|�\�Ŧf�[�y�O�+C7�ףuP��T���n��l��T��փ�h�.J���[����$0b�!_�z������ĭ����TC��f����.h**�r= ��R�9J���xHF骲.�qH�(�Fk��x�n���<-`?ٴYժL�at	�e��-�~&*<?��µc��k��O5CƭU� ?�D��!�ILM���������#+�S�v��7v&=�/�*��%�m��h���r�=q���^.�1^dj壞'�e��c/Sq�,�G�������f��W�cܾn��<5��[���E����d$��R��� \ ��,���O��61�������>'Bi��p��Ҋ���kqU��_�![��A$�4}��~��F>e^T]�m��c�5:E�[n�R�m�;�N�`=$�`����h��٥��*�|�T.�z�a�u�y�t�zq ~��'?���|g��A�w���v؛ 
��o�{�� '��N2�F_Qn��d�'su�L��CM�Pq��x�!U�
���a'�Ei�S%����� Jޔ�*��}cb2��,
�P�kS��1BX{�4���,f
�/�)ƅzl8�T��[SԠ�i6*f�8B}�  >mQ�g����[�N�M>i��5Lc|4��6�{g@�!�P�<� �q���Mg���r X�#L:}�v�74�
�H(d �R��֜�V��2�5�!rR���>���8�3F�_���z�����Z)����=֗}<@��OaC���,��������,�搦��ŀ��u��=/@�(6[��`�Fs-��V#�W?�(�y{F"i�P~
8�a�2g� i�����A�[h���6?����gH*l!O�y�����${�^�^ZA1��e�di���e����&�|��]����	ۆj��O.繥{(P��?6�*x�w�1�t�����W��f��{�����Cv��ub�8vn83z"�5�NXH�/����7�/,����U>������!A��1�(��q��| 5�I��j��_�¬d2��qB��R~ ��2S��=i��f��dM4�[��g�zƈ,�$�j����UPX���zb���C��Tb�;^g�6<����,Q*`���'R�R8����M�/"�#��4��+�]�k!]N�3-c�m��.j��y�b�ja��L�~_i�+��_v�Y�A���4,C���r�r(9�n���9�P�e�Ɇ�,�2:%@��B��eAÕ}S:�Y�����`z�����5�\��vpzԥ��	�ހi����c����^��Q�lt���?<�`aоH`I�h�P�re�� ɰ�&��>P�i�R���t�5M��:;WV�Ԣ�O ��j���	*|�oI;�s��J0zN�ٰ�=��qi�QR�6n+|�T!����L�j<kT�'�t�m�.�>��\�w�Y�P	�];���3!)��C:?����,������;��+P�B)�1f��;��9�������d8r���$(����OK-��p�X����Zs�?)LteO��4�L.�
c9�F�ݻ�E��q��f6��НǰΒ����]�-~Y�B}��N��x@f��2��nE�4͆0oLŎ@Ng�d�+�\�W�7��+J`����ͧ���<:LP#�3�11l���O�9�����G �;ݿ����&���fw�׻�h���!�R9C	<c!�w��Ը�� K���
� �w�`���O�U�=L���Jw0���L]�ƚ����Y��k�		��� �n[8%�<X6>-�,]��.6]�l_��1��!
�����"IH�Ťu%�R�f���(#�.�>������/&��'�4�ᒷl�j�Ş�t[ߜȚ�k�5���y��ֽ܏�F-"c�o�7��/.Z�������p�[�V��fQ �H \{���uN��9�z?�v��e�UӘ�6]bT��w?e�.`p�c��Ԑ��������D~��;��f42w�3���ȿ��zן��7x
�B3L�����xR�Kv�M�&��j_���W���{�V�&�Q��zdQ���=�,�{��-c���p5�r�c��F�2�\!q�A����b`4���{�<й�X�&����V�}�2�Έ����y�*O�;ORf�O��y�L���L۪���v�~����t��G�H1}�>&̪CėLz%�!�VH� �+��?C��HmZ����3IO��P��}U}��e��F������Sj�C��x���#�:�{��D9�F�mA��sz4�d'�f< gy���r��	Io��E4��^�b��Y�88��0��U�y��#>�~1F�;Z���|�U偘�6�?Ԗ�­�e�Z�dK/�Ǹۨ�.��4�8��фf��K�
,��m���_�q����WO���K]�|I��O��!%��`/O���i�ާ��s��$�1�S�A)=|Hq�|�3��裆�K.-0N�Ϯs4o��6��M��ЪYl�gh4z䦼-�C��O'�= 9��(��F�L�ÅbeCʿZu|�9Q[&F��?c�I�ss4W�"0��`$���pXe��C}��K�.�r��iLD:n���ml�n�*&d���K
�|Dj� `'�A~H��]}�eNT���`����|��y�LC���e����cQt��A�d�F7�����Iy�8S���Q���1�G魛%.\3V���zxȂ�n$.�~�8%���K�������R	�{L���3�{��o�!�Yzv��ɺd�elV@�K��a�r�`�ށ�)?�F�³��L��x^u���]൫7S���$7I�j�#F�oO՝�f���#j��;������a�}dNB�˸i�#�m�3ⓓ��B#hv�Dqs���^)^��y�v�I��4.���6��5�`p �R�=�#��}�mY&������1{s�g�&�c�y��+73��^{�"��I}�����Ϙm���8��{D��Jrh�+��a�����zs�G'j�2eP�&��N�X�?$Eq�a���tLԉ=��M���r���Lo��d�B�"!)H%�e�_�s�$C�Z���mN.{P��5dwf)���yeZ���7_E����E���*l�����-#,T`"��~���z�{Xu<�%ݐ�����������1����N�UOD���:�s�[/$O�vtN�Dѿ��-nL�5�W;]�E�i��cy�urKT�
��:M�J4��
�b��4;Y?l�V���DX��,e�FeO���BИs�\�X�~Z��g��&���
�h0���h8�jM���j���]�)Ýj!uas���;�<�{�-jD�^��>���!�7��C�4��"�X�w�:r�����f`QP[iu����g�91zHS��@�]�$#���B��9����D̒S���"
�-l�����|��ID�G�"��$6�<�g��A�-_x���za�+	2Ǳ�Y&b�yXny���w����8A�Xќ�)~�8�uw�XX���y�e��ߐ ���[7&�8b�tW��篑�=L�
{8
�-�3��D��z �vc�]���˞�
J7y�n�~n��t:����(j�ī~����fº:#�R`;��*���Y|u����Vu��"�	�/��/@^Т�t�=r��q���1��?��h�K��.y��4��q�)�~��3�%XU���A�}���ݐ�cxN�5�t8� :�Do���?J�����L����٘9�O�kƶ#�O�W����Z5uJc��F��+6,��썸�_�\E�F��T����7��2���)�pRDߒ�Ϊ���]�����M����V�⺒��T�{�%�jF�H,��(w+k�s�qUV������D��5W�� �p�Rp��v�\��Lb�t���M4���w�-�N+>�>�TxEؾI��SD6�(�Y���-��#*GKS
޲�����?pj�z�:ϴ29�+�-ҏY�I�b�9H�H"EJ�U��Y �-�;������ ���S��z�i��wm/o
�R��[SC�0J�t�k�*�P�C�����\��I
,xw5]n���+�H�����8���&�%��K���Y���:Z�%{��;�z�
��ԗ7�Y�6����u��1�kZdA�H��c�!�v����v	���b"�
m$�e`�gR_���Ԑ]{Z�8&��yՃb���V�X��jZ��Y7�MW�Ζ����~a_c�e��L�$JV� >��?�N!��];. L`��O��t�#��#�I�Ezב�p�ޚ�g��hE�?(~֛�<�Sp�^y���a�N���{�z���Y%�l.�"������}&F
�&�xl�6g�(���]���SrJ90Kk���d*Y!���8b���i��#���]@�1	��v������4:mA�l���i.m�A)o�I.�b�d�d9��:�<�r�������3�4��5|9hr���ш=e���wm ��%1�'�T�_�d_���z�3T��D��jc����ˁ���Ln�� k�q��M®2��ʮ��w:a����ي��Aqy?���� ����* �f�a��S��n����	��ymW�*{��1� )A�r^�����������R���>��<}�R'�p���~/��wa�۠��P���1_K��3n 2�&��Q�ƶ]S@;�s�f��Wo-�..�������x-J��j�+�!\�)X"�����G����ey}��=���y�_��w�¾���w����D�ԙ*Gn�čw51�d���5\}}�_7�/�̃���'��_7S$3�Q0�I8y*�F�gApQ\��2��:�\I�������N�V�(��M�,��n�+I8$����g�u��CW����V�i+�ݨ�g*Ճ�V>�K��s�% �53
�Z��g]�2L(�p�/c������	����̗���Y%��Bԝ�TB���� �Q�&�[��t��t��	�u���Bz�`MdA����9�gCd$��B(�Ⱥ,��n�*�)J�`��߿��.�B��� ��SLp��MrN�Ig���  A��v�+�Ww���S,��K-���S+�*8N�)z@tT�d��M�7����K�8�8|�UMf²̔g�]�� ~/�i!�cZ�3��|�]㎙�g_Ыdtb��{/����1s\a���n!�Ь��n��f�z���	G�)"�?E8����	M�#uK��$�o��˴ʯS������n�`S���gj��m��Oz��K��ѝ���֒տ[������dpwݪ�J|Y��U0����%{[���K����x�-4˿mvMN��}폝�01�����u������mv�)ޘ��G6�{��ȇsvH]p<�, n7�(�&���i^jx����y���M���9�_�><�f�\;�J��M�#z�w�]�:C� ��vϪ�W�"��v;��(,�aƳ��^k��x���݃���^2����Z���U�����hp9-��ˀ��(<� o#�Z+/�B5|��>�h�Ҝ��� ..����*zKO�%�.ʘ�KL�t���!�&����i����AQ㺜 ��;+2���������%���O���B%Z[b7���0|M(�V�&D��(4~��I��zo���'RE��{.u�oy���bdC��y�sN[	��͆Z)�Į� ��+��"1�T u��j7�]bY���h1��R���x#4��_?��Ēp̩Y����w�4�x�+��޺�!��c+6�F��ZAi<��b*�e��𺎝���%0[9���)0y�MI�[��`��&��[a9s��=��� X���a����/��y����La4K�����[�F�CZ�{q���7���u�$9�8ES��U\*��]�¼u�Jj\�����p0J%i�*j6������Nk�����O�=3U[�b��Wf-W�]���ۺ�C�c��ǔI���6{�C����.�wt�X�6gd�����T)9�<��\�jM��ܑ[��c����g�	�����L�j)��J�xr���*T��P-��yy⎄��d5D[�{Na�3j��U�:��oyF�(}�*��V(�N#M����į��0�8��chʲ{F��ذ5���r�_5���X�z�~.�p~>_��)�(�%��������oM�0pr��� >���0�� � ��ZBn���.Ό��{�[�2�D��sa����j)R��ۺ�
!����������Y=,&z޴j*�际��s\q<�f3G: b�������z���*QF��F���0&��-�����Ǯ6w�!�?��y�)�#�=	Vq�)��t��%��L'\Ƀ<��0h��k��ŰN0�朦�BAp��v�m�GU̦��QN�9��p{s3L氙��8�m�;�܎�-Ag~�<P.��O�ۿL���<���jd�صo���Ң{�3�O��+C>+��߰�L���<����H���Wd�2L.�sd:~h��������%����l��l����27��	5��V73*T�B���VS�
 }�h��1c��QW�a�3�k��D���j�h�׊%��TD�(|�`q�:,ݴͻE�A�6M��#��~�ϓ"���m2��}���x�������g��4w:��"Ėrx�D\{Ke�jo���f�듲��9%;hɄa`�b����EQn���$��<��7�u4����-/S��m���P�< �#�~{�V�
cӛ�@~]��6�;��g�f���-��(ai!�OW[C㫄?CX�G�5�a)�L����C��%�*l6Ī)�¢��V:��A<F�a`�K*��V���4Q$��v�8M�����c����\��t�e®��aAZ�a9��}ʄ<���#��=�H�ç�y���d?͍�$�����v	'�b�����ޅ����N�~�l	���F���bT�J�
��Z&]#��B��Ԙ�_2�����z���̸�)g �Up���:`yyݞz�O�3E��9w���IK4�wW�w�(�[(s�z����x�?x�cT�@��}�>� �](R�upkLB/<蛆���$���c�.�K�;��V&��������j���D]5���V��A^�J�c~o��s��t5��/���MZN��장��}!���ŉ���H�F�p��SQ����p�c1YU�{��^��w|�lN"�	�n����8ݡ�`��*�����9��˔���=X��pS��0jN�Z���<���0`�ƌ��}�f]:����L�K�L�R�x`�H�"�Xn茻â�^�a�(�+��ĢGr�r�mCF�`��~�x�^����s��U��c{=Ƹ,���/���d~y\! D3�h�L?>�ն�t��l]�;jJ �r:~Ą��/�jA>�K�gx����[�'ȊIp���Bu)��w�Q���H�fzB���D��7����������6�RuKȪ����V�βV��x�o��0]�d���w���=Мu�ho�[r��#�8�7D�i̍��^+��E?�"��~���G�!��:�]�2$k������d�`���zR	oy�C�`���銃���h���hl�Q�j��Tmm:�YN��K���&��' ��2D3B�.�>g��CMj������o#o�t�42U3�hf�zϐD��F��@'�K����޵*+3]�b�
�������8Ft�<�(��rTúw��x�q[�L����� �9�4n�U�ZE��j�k dB+�#ΧF���8��p��b��E�Ʉ��t��#h�����(	1�6��7�pAA�~�^��g��n���4}����>�8O��z����xZ�#]j�]�P������^�叠�&;>�㇓�U�w-�73�!@�5�:�M��3.&��Ӈ�^�[�ϥ���z�����Ū���^��ڌf�gT޸��]�X�$�v��m�n�yX֖ˣX�J�T��n��`@�}BM<.kȵ"��{Prm��)��A0笍z�=Cc�j�'C���w�Պ'B��W�w��ɄdS�n'4��%z��'D������������ϻ>��{�L�#ӏ{M�Һ.1�sd9�T/��x��9f�$d��֋1o�����~֫��13��s��'��ƒL�uc�d��v����/sn�d��!�
��(�lD-E㖮!�C��Yݜ�����������c��Z�ۆj����LUc#���'}1�/��G(��>����ٻ�@~w�*�v�v�x�Jy�_�$p#`�!M�JP�ě"�ik�ʷ�/x�v!�=��pZ"	l�,b�T4�g`�u�[�B��e�Y�a�w���W��+$F� :��H�JB�y����aY�4��x�������ʓKH��<CC��Q�D��R����aj��&���67Y�b�{<Dؤ�bCf����D��:^/k#FkJ��w��[R_ɏ�4d��ў��!��A8�b\Y�Ƥ�q^�\jN�DI p����-��r Q�GW��A��kc>��I��(����sx�EgU�6��Ls��,�Dt�`��v�a��L�g�~�3�����U����f��ʈCb ']��M"��ؗT	��!o�̗FL��P���*�DʡE�`��̈́O��Ի�Xt�cT�F�<`�ߩ��w�=�������:��FD�5͎6�e� {�Ճ�<�$�&�����.�>hG2�V��O��[���e��4�x}��
i(7�昵:��u
g��Qف�M1k���Vp���3��v4AdM8ц���,��>�G ��9���	g ���2�\�_ȡ�!�.�A5!压�R�w�b�� �pTL(3$��\J�K����nbyz6�����/:T}5��Kou.�=T8��3֩�i�ZB�3wR1��c��r[�wڛE��o�k(*	?�*��f)|-76G2��l
ݾ'ԛ>x��I�w�v�z?A�-MQ5f���cJ-���z̬��&��򓘮�ՠ����1;��0���e����%���w���Jk� b����Uq������������A�,��ڹ��W[�)d�9���&\1���m�_?Ϡ#��x�
r<�Q[{6�g�EI����Um��g0C�0���bL���7y�:��ա2%۸��M`L�ں��yϦ���&�4sI��=t[l��F&^u?�pA��S�d|��9,�i�l�Z�,�.�V$����և&���?���������=�fkZ�����X"s��淚)��И3Zՠ�Z/��+n"�W�9�q@��G�������q�z��5���'HF[M̶��T� $,�]e�L���z/����P��;���L�Z�h��'�@+r� *���%_�;�����2�IK�#疘�%u�����g�<w���MO�? �2g�P��2�S a��f������3�s��82%m����w܂���6L��F��|o#�lT��ZWg���>�/�q	��l���!8�FPZN�k�݌=G��3��2��2�/@��x�D\e����kg�j=[���j����\giy�$���l�/�[_�pt�>��M1����������S	��aJị�.*Z��`����Lс�r`<�wD�������C�+S?�D�}Z�f�Kc 8gYQl�F����M)>T�Kcq��*���6n��@?2FrW�J�+@��*&dE*?�3=7��T�7���I`�Zު�<T��׵[C>�{�K(eن㤷^/�+��� )l��)�����	��J��g����ڿ|��L���[$���2�S  L���+��A���}e�SN��/����0%�5������8�ߩ�y��������U��z��m�ܜxbQ������h<�IŅ�(����X��Qʍ���6/Jv��{eq>sO�4�t����z�3�+���Sy��\OW@��%����|M�↘*������©ʐ$E�f�v�r���c�~��h���:"��xl�8�Ao������@��!M�x �2B[4���8wPw
c #�������H���d���H[�	ǥ��b �"<�  �"Jz+�����*+P��>g��9���3���}���J��X@,�g�F1a`�J��l{��gſBS��Am.t_ufA΅�9U��<�"��\��egi��c����E��V���"e���h�!|�G� Iah����͝�9��砏53ݲ��P')͙ӏ5 ��9��3����K8�'P�O�r����g xu����1b�G�bэȧ��ဿn��x�$�3�bh���[6��2�L��n�XG��[�~��m�,���Z��t�F���YF>˪���(�,�$i�̅[�L�ŖX+�J�1F�%n�Y��֝�n�����-���c��&~X�]k,��|�©�bX,��c�],�Xy ����Wn�b�-tkY�T��d��U�c����1hR��q��YzL֝�W������h���Dɐ��)��R�M��;��#�P��,\�H#	��C�>��R��
�Q���w��w��cV�=f�vj�LCZk�W����k��rp�ٜVL��$���N��f�zN�N@�=O��5'J=OnJ��snX����Y�S6!�38r'o-o�WQJ�[Ȝ��Z�x���%��.km[��/ۺ��O���>�D�r�{�'Ԛ({���<����h�=\�i~\��ca�z��L��.�;w��|N��o}
d������f�UޫԆ5v�L�lOJ�s
7��WU&�p�b���Q�"}��~�=}ww1�s���q�񁕑���N��tu�o�s�+id��'&�p����d��9��v3�:S�3w�Òi�sN�8/:��a���9�A�P�!V����=�V�\�⢿�J��6j���[H1�|�W⁷��uz]�g7G�#	� 0�ٮ/p���ԩ�U��!'��5�I�e}�qn�NaMz5I�}�h΃c��z�r1��bp�I�޳����Q�{n�i�]>�����`��g-m�q�w�ǩ��[��N1<�h�hv~B�����#��/v)yE��z+��2��ǽ�
D����7y&H�Bg~5+�I07����*�bp�W�A�"�Q��]�G��SvP�Pj"Q��#,��V)TԱ�7�P}� ��R��|(i�5���-&m��䷑��c�"��1�E��f�z^��	v�1�fKd/xWG�ڔ�\�ˠ�@ӻ��mp0Iuzs��]� =���A�Ah{̒a;=�#4��s0cص|�/�z<ȧ���vH+��T�c��x��Vc@���4�/��GUI���!�J�����+�d�zA���"*���I��Ǿ/�|���	��[��T��X�d�r�0��i̤�+ԥӸ��nT��;Ȫ� �y+� �n�Te�a�ӡ�}�T�N�} �xY[��/�ȿ�����i�=�C���ݙ9�W� �Mo �d���	���Bg�'�Y0��Fq9i��9�n溺!�m-f��0L栧�;�_gG>��w���[��	=�K��lչ�e\t:.Q�T��y����U�o1���I\�˔����2�ߘ��* �qI�v�[eC_7���7�,�g���l"��~ ,��yk����T4�e���70�q�#/�^�n2�O$�������$q��=��J���y�t��F ����n��"����uh%.��nI}�pUۍT���w^�.��Q�??�70�+isZ4z:^��DS~��[���E�>ƾ��Y� (�$��+�{0�P������D��D��t�`�.��A��p_!o���)�:D�H��p�81�
�i	�5Vv�H�X�ө�!m�L�e�C�q�z�rA< ���f�ܧ���4½`y�`��HQV��$X4fa!l+tU�m�y&.u�Q������h?E&�(/�2�p�����%(����z�e�ǹ��P�w���UAiܖ�i��J3J ���j䬮�${����)������Z}�%�wu��J�-�ko|�p�#���+�����ݾa�DG���6�&-��l(.W�j��X{y�XbqU>L�dܵ��3��*��&v���s�Sʄ�6m�wi|P)Q�YW��H��v$\������ ���i���=P�I��N���k[�1�0��g�3��	GP�y��^�����_
	�
6���t۱~�Q �]��qc*tJz�G�m.r����fM%K��c��.����[�B�s���$Xe�KϤ����K�F�k���R�1/�Q<J�`)�[�p��)}Z�2_'}xR�E�X�nʾj�S�_�L����P-��l-vU1��k�&	"�� ��������7�0=Cx��v�_�@�λ|�aUyAٝ�j�Oj�w��������u��u���Γ��(ή�@������:Y�rQ�}�pq-DĨH��R<��th����u�1	������qq��F#�z��5cB�� ����|¬U��OT(�=p�8���<�j��բԛ��{�:���MJ���?d�n�W	V�eF�6wmmJ��6D�q�?�F���x�:_V��;���6z��8�7�TW�N�4�'Kw �Ŭ@Y;ՃpB����`�t�_SZM6*�
3�X�����R�J�8��(�P܁�a_F��{�@vm3#Cx�Y���Sd�������T,�ًB�VЀ���p��¸��ݘ[���Y�v��	0��؍(>7����F��j
��Q1���[�yI!G��ӯC�9����-�~�]](
L+N�]�Z��K�W�S���^)9X�S��욕%�e�"��aD�8�Sx�e�ˋ�4i�S4��ckE#T��;p����b�S���s}W�C��J%��;��7M꤆Ց��chN���S��}�Ff�}HYN�$}#)��t��p�ƭȽc-�����,ڗ,"n�&ٜ�\)ӫ��)��x�����f�D������TD=�0nG�eR�)�EEޟF��"�g"��kda��b�ЮЊqK��#������Z�9p�Al-����P�h����Ņ�C�-(�f]��o��!H��LF��@�P�V�#ïK'�����{�q���W���<{���/�>�̒5=�l6�5\�TR�ZӲ컁�B2.}�3`�R�i���
����H��Ot��%"�a��g
����6���N=��U����.��J�-4�
���t6�){������@��\7��ψgy��Q�2��Y[�$���W
���W1��a�D�A��h���c�7��	Ջٮ;C�+�me�\'5��O�[ �a\K�g�>6���T�P{�\U�B� �������[� t�e� �dba�k@���a~С���T���_��]`�,����:'�<"Ȁ����l�����ѵ&>�:�oC])����p�=GSM`����,�.��h�^*O/�"�] �I������yyOiэ\���;! ʦ�%��u�@znQh�"EĽf�8ı�u���}@b�]!<v�]��A��N���Q��A�蓰L�s�F�mCp��nQ���N@Ds��8��m��^���B�B	*�ߏR�p-T��ˊp���>�|�{T�r�-�����7&�$�5^V�kH�kz��7R@k�0�k^8�:(je�?.C���v<jt R�W����i\p2g��?�T��қ�m�����b;H+z�L� �	�3��%9.�m��bd��s��&r��X�De������+F{M�,�;���*�ۈ9��|�X6������	bA�J<ҞFVV; o ��6��	��n�k86v퓗ۉ����#H]�I�H�D:R��`T�7M��	�sr3�8�|u��δx��s6��챇�,N��X��-#+��լ��vH��rB�� �� o��VY4ܑ�31����Н����(�2�j��tއ��ޘ�)/�f6K�D�sˡ?��i�Bn�,�Tz�SL���{$[�mS\���ԉ����xY�$B=�Z}.�}�R���vdY�G?�ԍf
ݿG����|��+^Qd�+ڳw� C��<�:���^��U쁁�sĐsy������L�.�# T�o��Z`�\;i�l�m�%v7
�i>��ճ3���S���eN�lD�����)�3��=�Uz���D��*㢜�HCܻU��:�Ӷ�VNJL,��N���Y�(�L�{��f��X!,�f4�l�۶�`m��,���)D��{��Vzh�b����Fm��0ƭ"������D�̨�[� ��<�j����֔ߖHrQ���bD���a����v<d�ջ`Ǿ.B32Ҡ +z5���#ot�9�Q�_�JLL���x,d�IѠ�dZ�{D��g���	�?�T�ߠ�h5R*O.߹�\����/�]e�-�:��lW�a�G��iYu�$�N��1�]T!`P��0�k�?p%Ҫ��a�%����� �Ə�/����U�z�S���S#>�D�ڢn��,x9'�ym�4�f]��=e&\B�*/<�-�Fr�t�^b������/�a����EQs�E����WKG���}���+D��߾�m�t�l�uב�V�K��(�תL�^`Cf�E���Y�b�xGߺ�5N>kž�Y��s��ܡ�5bg��k�2�]�@��Hp2<<��wP�-�bFR)nE]X�G9g�osw�$�S�`~�\�^��U����M{�i.Y�K0��u0�Ī�Od��
;�Ӻ>�|/+.����oA"t�����=w�"W��1���g+�>�B}�)�����ݎB��1"�G���y�q|�䪽�RdF���\�N.��h-)�,Lю;�6��/F�Z�΃T]H²�����Q�OR�A��e�N6˩�E�@4�Tnif\3-M���!������D+{�	��eK�N�UB̥G6&���*|vJ,H�8�|���Q����B"}�5�h��:U�OQ��Z_��3���!�}繢����0/j��k��t����KT6�c��~
�
|Vݠz:��`��&�	 ��h;K�C��P�O��f��x?�T�^�q��o��f"e�� Fu�eJ,��;� Tqh��EA����#p~@MGJD��~�u�\s��|�ES�$��腝�$g���O�'�B��?����7�K V�Ù}��YgT��VH� М�L:q�u�V�P}���W����A6�F'����s#�嶕��,���Y��}�X
�"����׸Nx<5���:6kvq��Y��41�|�;��-EF�^^�s=���t���K�P|�B��"����Ȝ�YwN~�f^���3Y�}5�\-�ě��H�1¶�]P3�2>,���Y�c\�g�c���g8��Vb;��s2��<���;@��OI��O?N�=��"Y�� ��bۭ���bN�q�";�� �R$�~����+&bI"EdӢ����ɉ��fT�#�*�F��w>��td]��W*�u��Ŭ+]|#m�%"�A3d�Y���Y��i��~�]�=�ȹ��_�����y��4@��'d��+���P��E,�n��p�{t�)PDD�E�ꭾ��.��PB�;`e��+1�j���(\@���SߟKz1���O�S:��P �#� ,���LE�Mi̚y����8g� �2�X7rNV��=Q(��#�Y}�"&�,���fԠ��ĵ���%�1~-�=U��#=5{f-����x_�+
C��F��O����k����X�	C�E[I�h���ux�9��w�]��&��"N�f:-I����q�D�=QƲ+�w@���~�c|�7��U+�^��W�u���~a$uA���zk7�UX_��\[~��� �������'d�����$���Z>-rcl�o+%ݲ)�TY����aն� �����`�<���|��P���d�� �����`qc��8���:�IK��#v�{�փ��3�."<Y��|�[�i��)Z7�5o@M���9�薳��H�S��*R��>�S�y�5�������(�^��B@�����@�DUS#�����g��)��'*�B�-��wT��Z�ĵ���x�I���!�,�I8G�TH������
���\3s����$����~������>�[}���X&����^�~li�;_?)�.Z� ��u1
rW�ȏI�l��P��B��xo�Q$��aQop�U��ts�)JI;j��,�sl�j����l����SvZF�~A�(��<���Sm���Z���޳����d�X��MP$�`yx�%�0�
��C�Z��M�UeaF��ޘ�����I�&���B����f\�^�q�e\-3��E��;?/����	��]�<@�;)�x�$���y+[���Q���L��lu!��⌃�C��j�	�ԡC�.)*�J,���_��,��P��=e����h�'�`e0��A��ߑ]JH��C��0����|��5��zUh3���K��hZ3ƲOG�/�u+�Z:�5�1����dؑKz�.M�@��S+1�<}K�X_"�	&�#�j��s����me?d��B��3Ug?C,W���>�u������Ic�+xG&��#%�5~�|�J�%`C)�_xyeZ�j�/�k�q�P+�.a�5�x�����������8ՙB7	]u&�.�H���:Bס�y`�Z=Թ��kC̈́^���x[_<��gM#c�\�-/�E$�."�^�Q׶�������i\f����֤�K��&!:�d-�����ʡ���@��W�����f�m\�Ӻ|t�?����jA�%��{��W#���+C�Y����?	�ݷ� u	"4��5D����M���;�<�����e�b�O�/�[����X�8G���s���	�D&�
�:^2v,n(>�@��:�L�)��$�+P����t�� �����5���q} �:<�-�)�㖆����!�2ix��-D��z�^��ݣ2{�7�ȼm7BCǆV(#�bn+�]�x:I��f�Kx=� �"?�Bw8��ں���O�Z�	rAo`� �3��bP�����IX��x��+J�Ex�Y��
��l99�y�����g���h��Eջ�AT���n��M?�q�@G�}���d�]�t�E�[�U�p�AH;�=��D̊���Pgt>D')���Q�[�z<�rH��Z#�H�\LT1�d}��y��\����1�L�*֦=9����]��ˀ�J$a��Q��9g*i��U�z����̠���f��¦��Zo4 s{��&b�图w1��h�/tPr���� �͠����s��S����!���K�̺Fx3�|+�y�&9�t��܋'0G�1�] 2�f����$���J@o��I�Q�F�@��O%�
.��4&1ii#:_�x���j�V%g@���s0��PmDKy*�l4�����s�)�0�MPWK[z0$-�0��}_�ҁة��t�N�?c�@�y����X��H��Wal@���ޤJڋ��(;��n}isF����%}�-�jM?��P�NI~	'������yN�:e�'��Tqx�wu����ڑ�z�������-eM5X�`������1��y	Il���Ú���-��a����5B���W����0�W)-�)�g�RA��<�p��K�vq���W$U|��)R/�hWw��bS����Xdw�F�r��՜��x��	+PE}�F¤�b]S6=?�6�KК��+(�����Ѻ�2�G\��Q�<�9�(	�`'>;;���q�R��)��<t�M-'A���k��T�����C�2�)�_4�v:��.p��q���u������#i��msS�E�Ŝ|�(S��(�̃;�s����,�!��v�-�װ�;��������Q�X��%ü��{pO^[:���&I���.�+����r����#G�fG��AV\�t<�dKp�w����=ġ,�����@'�ƒ ���7a(�0��s��+Ĥ���)��'Η}ɄI�)g���������F�	[/�	)-�|v���� �C���]��u/~;K{��2�"�7`��~�?uXQF�T~�\P����2<#�=����[sQ��L{R�\f�kVd�Y^�HM|f���k���)��e��p�����Z�pdl��f����։�ֲ��(��}M&��G��K�=^"m="��=1q��^J����m���ca��I��9�c��F�����2������^�2��x��a�sY/cb<dX��UW:s6(kq����>�f����P���c�q��Ǎ�_���5�S�]7W�Ot�hx�����l��"ؽ_)��5O�#�3�~X����M�٦�bj��.�3���?�Ǎ��^� ��CV:�1�g���E�H��U4 ��d���u7�!V��o��v�vX�+��5��,$� �I�(��cۅ �CRf��J ���r�� ����۵j���磎��m�� ��h�2���:6��Y`��f;r_�4�5+P���4z�����$f�_h���*�2��GI�!�J���ݳ�J��Ƅ�@�5[q�LK�Uk��V�3���]��qu%I5>Τ'���m�d�ǦV�s�}�o�� "��+�r6���]��i�f�U�c{Zg���|��?�����.�Q �KE�95�v��k�~'����q�:��H<����0��ħӳ��J�WZu
�A'��%y����T��&�Ҏ��&&1|
�q�y?�j����~��8H�ej�w�5#Y=A༃�)ϩF��$�l�g��ݬn��%�������γ@�q�Y(����u~>z>����v�p��P�>�$��׽>�^��q�5�ۈ�RXv�S�}F�~�dj?Kb˧�Rt�k�TӚ����i�Ã�Ɏ�9�:�$	nr�����.��^��o@�}��o �M��F�A2��:<+ �sv��f�Ռ	C�^|Â�( �x���?�LI<�傜��y��{�e:69��e��s�E�f���������.mz���Ƴ�[Ύ�<8U5 �Y�������2�[\P�G}�������;�O��iӘ�hL]x&��7?�s�U�G��ȧ��K_�xƉ�����|X\�
�N�^�Z��2��1�I���8u�ܯ�?���O.0�s�!�A���,?Jb�D=�Y�a��X����eXͣ���|��	v�;A��԰m�M)�̶d6��B��0ao�V:�\ؑ�a�n(Ȁ��펆-ᕤWu�.׀U����G�P�Np�K�Z�ή��+���w����N��f�o4���
�HM����޳s^8f�4�-��n ����q$�"ǌV~l:ZY�bs_]����=�aN� �Ơ����k��O���� 8��h��x��@��Z�u17((�T�kb� u�x^YW�(�u�9&���KȮl���2y�~��U�{�� �m�����0"������e���rR������+�h�?Wp.�"�7�D|�1�RZ���0�p��I�p�i���4"����Qy)3<I,X�r��h-*]6\��	��g�O�o�__"D{ʆ#����m1�a�r'U͞8KU��1��=��*�������Y�+�GT�R�7$�1wOh�G���/(��+�D��gD�>��*G���	����2����!��]�Ə���Cp#�Z��`�f�0]��7�&@�_��Zn���#q���D�(On�u�Q����^��z�5�T�V-���3-�SaV�4��X�k(�ۉP$}����&J9�_�@�`�Dy�(��J[1Cq���o�l#��/� �����b;0�j�c�n�b�[(�g�#~��䓘U��MK���Զ�����@j&�Jr�Z�;�<K�{eg��Ύm[]LW-D}��W6*y<��hu4�is��<u����/vss�-'��c�q� �ȉ�!��A�V���Џz�)�����������7J�B�r��<���W[���V9��G����YTe}�V�Bɭ��" ���^?o�_�h{o��]�6o:Ǹ��������G�J�jI���[T�$���޺\���~�PO��22
-ư\���k�	���ϞT�\��e�q��25�9�͇Y�c�6�]�/^i)%�SEk6/6�?~@l�Q���'v:�"�46c[J_�>��,/$�+�=��hj/�<كâ�v�0��S�VU��\�ڊ.�jN�pm�Wִ�$�ܿNB��xX�GX��4�\E�Pa����O>�|9���T� ���D���F�������t��r�c4��}:F���ff�����%�`�Mˣ��N+��<ڡ��\��0e(y���,��"c ��\G��&��U��&���^+zYD�Z$'����4�����	���h��˧ob(Ok��i9� ���0:���c�8WX��*�5J?�҉Y�+4/?k��D/��{I������}�"�$wKК�]|�xd��Y�ו�u&����U3�>�wf�_��J�t��]�Vk�%}b��ot�Ygn����Z�Qhz�f6���(o�]J� _�<2��8�E�_���N���T�IM��k$�IV�B�S�o=���2��d>��,��B���&��g��g�)����B	�52+��]tX޿�3���Ҹ�E ��*��l�f_���u)|d��
.�'�+-p�ފo��M�0��溭���Z�jm4-V8�r�t}5�����u��q"!�[@�?a�G��(rcY��j@yԠ�_�6��>�M���]LQZ�A�G�d�����VCY���&�mֽ�� ��^4��Y=.��>�{��>[��Fi�u��]�qM����b�]�m���w�{Q��Z�/P��^k�j�P5���J�Dr"�|�*�L�6��NC}����3�.Ĕ�P�a ]:Y��)	����E����W�ZQa,m��s�E�x���!�-�:LU�î)؝�m#ۺ��yVC�R>�h��us�r�t���cu��x�8YmF���#���o��h�6�Q�o�2��Ț��*1ʶh K���&��{�`w���,oe�ѹ�h ������D���ĽNQ<%.Hi\�x��_�]L�G�)�*f*F8̜V|xn�B6^r�H����P��XLK>�]yD�>�V+�T�R9�^b�#uqhe�T���-�3儚҃���{J�o�I-`��b6��UV!�J��ƶ�!� �.�Q���W��AEb3�Y0��_Lk��H���i���\���شYJ�W�Y|�
C��G��2�ώ���"�X܏ �!���e��[���`KR��PY�#Hύ;%�4o�#G��(�r�#KҔ�ڎ�!�Y�c�f槉d*�CQ8�K��d�Qa���^�x6�A�Ę�5��ڭ�Sǃ����Ox�����&l�X�/��˜�*��q_�^͙K���R$a�Pް*�c�ۙL�E�7*�C�Qi�8���V����v:��oA�8�0��=�|�F�_عqx���q�Ϸ���X�Q��ϡ��Z���ӧ6�_0P���B��c�����f|@gͣ���	����t
O& >��@s�13��Q𘽸��{t��UG���h�c����/+�x��P��:t�� �I6:g6�D�;<%��$�+���o��OmC�4O�[�:w>�R�;��Ժ)Ң��9�.��4�a��0jYZ���_�T�"8��5<���߮[?æ�y�l�b��@�̓\����V��:t$[��q���R؟�Y��<b�<�����"Y��=���y2Ĩ�w��7��S����ӆg(<�������,˗*�,�Ӱh�pF�q�$8�H��߆=��
���C�X�H�6+��	��Wk+p�-J\ӝ9Ά0Z�>B@݅���-��Zf��E$-��	p.��b����������՗����)�2��V1��V��I�g�C%^�ڄ[�����U�@��r�'�1�cq>��f��_Vs�>���R�P�T��X��H8X�a~fM����X�`Oe�9~d��Ls�Y��H�G���6��$$�������L�F_��(4˼���������oZ���6�.ȮpL���i�4���h)N�9�f��o.�r��m{u*�-��dY�;�[[/��g�1t�v��ӂ�B��l2�x��iCd琰
�Ѱo1��S.(%ؕ;<���xÅ�Y����r�M
D���b��ؠ/�b$&�a�knT�}ĉ�`�`�#8��zv�Ŀ`(o�e�ϕ���l�?5r=����8Z�j��_��#7�h�����)m�Xr��O�(_�^�p��@���x�Wlȭ=3S߂�Y�zy]Z���F�z%��oR�w>7����WťO�Tn8��ޗ�ޭ�D����3�[:t���G$�6s{�c�c�`(�,}hI�i�*�2c�7leԽ8{ɷ�민�͉%s��x{�Q�QJo�UO��=GZ��N�����p���J�ؾ�9�A������Y�	�u� �������g�u-�ܱj�W�(�ͧ���khG+�V�y��
�m�%{y�|���Kh
����^��ܬ��l�4}�\[�qa_REn p>TaGJ㕳�����jO�w]�;@��PY�ѐ��oi�Ń�H�&�Fy�����?T���O���h�61���]0zP[Lu�j<�\��P����e�M���g�z^᫘B��6��,k|�i�/.��la|�����*�f��7(-���N�sp���i�Ŝ�)D�1��t����/ہ|��&[�',9��
1��%9�8��WH4䞾ŗ|��>H3e<x��K���� �f���ȂUї� ��fH�ح�=EM}���Ȫ�4ۊ�k��w�~^����I�=.l4��&�.�5�I���E@����<9$�j����'�:�q�b'M���%c�m���O��8��J&2)�<�"Q���w-
U��K>�7u�ǁD�6�Wr���YҐJR�/}��&4�@���*b��Q��>�P}�Z�c�U�U7�"O�=��!*Q�
�XPV�J�)/�_vu	���"4ȷl����w��5��]Ya��B%Zf
�79������|��fl�;@"�X%�tt������x�WΐK�C8���j�JJ�ϿLiS�yk
��-��\Xx��υ-?L[�CA�o��q�F1�����Q;��r5��d�S��:�[y�e{h�z9��M^Oj"��Q�f���Hǖ���Ċ=K�t	�����}�)I���*����v:i\�"�/sx��jH�R���`�\�]�
�Q�T\� %<����{��=,��d""�Ыx�<tiL��H�\���WK#�C~?'�ul���O��N8Z�Hb1���r)E˟R�7����k ?C�>%?eS���[�,`KѬM�Kunkp�j�# KF(e?Z�y����jX��� �BuM�ڈ}[`u���wy+�Oo��M.�/�fS�4�Ei�l.խ��c��֡�8K)����J�(8J�{�,�K�� o��(�y��$	��/�����W����k�$���ʬ���IX�/L9���o��©���<WXW�S]�\�M���<"�e�P-A�}~��Y<�����1K���
�QJ	�s"S�O��|Î\����^{��`a����\]���p堢S$}�w�O��Ъ����cf�fj���c�����A�,��u�ƬE� 7CEl����g�� {��"D���0o�	�O��uY�K��<A���-�á����׹�cq��@*�:�V5�#`���Ͻu� �k�St�<�1->'��rCB:/m�X��Y�MLE�ꇓ�Z�i����P��X��w�|��"]n1(�4xӋP'�&~n�{
�38 ����%�l�&�4{U�-�e��l�-�V9/�Ft�=�r@p�@�t��P(	���8� ��21�D"�r�5����	�mK(��Ĥ����ޑ���}�����۟���xPyd�E"S�c�`�MP�bT.�@>\8-�!C~��,.��Q��2cI5�j9��x��㹿H�$�n���T=Fq�p�ïBl7�����ׇ�"��?���o��Cm牺_�L��z����h�j%Si���U8���Q��`n:�<P���2qk^��uV��||�����4� /@x�k:��7lXBz�6�Ѻp'�x�/�Z*�� Nu����:PPPޛ�IL�]�E��G�k��NY��y�t�~a��W������^W���D�@����b33Dc�܂ĪPйN�\����bm�Ṡ��QHD<�G�k���^f�R��P���Rzo�p��v�+�lj��_�H^�rG��HW�1�~�zOa��ف���`�F}��P��Z#y=/��:1KdY����K��.s�zţt��A?`��;�F맖0�,��t*,~m���4��0��Ox�0�=���(>��lk��7J�h!��>��&[�����3��[S���r��:C�/Ja�+����Mq��pW:F�>�bkp�'��b�Xޖ�P���*WYqHw���i�j�xn��4�O�����3��B`��e����r���7�OQ��Ij�rn=��>$ �5 ��x�x��(����ɸ�8�}���M2��m��"��!���)��p��k��+�S1�y~�q��z��
��OY�qu�/V��DO f����F����KVU��_
-$s<x+Nؕ߆}G���˼�Ni=g7����Ȋ�=%�xs(��LK ��gR��m��Җ}E�O�H1�=�.e��yG5K�*U�īE/����%�s���K˞�)wf��?�R��8�����;�"��z�*�rh㬺�C�كh�N��fʥvVFv�r�����Of�@ʳ$2G$i-Mb�I�a��?~R�W��'��%5&޷5��C�T�N���V�g��,i���/�HR��,�np^�Z~�6f9�J�
�XH^=��_�ԓ�` ���^@��0e9�������ڶ_�K��^�<�Y8	jA����Z�ie��N����]�'&Dc!��<��їȲڏS0\�����ь+CU�yC�������J�C��E������F�#o:��� 4�!j4u�ȌGX�/!�����x9֊�e	>�c�}ɷ��r�E�k�n����"}�vRI�LDKA�>���$,��5� 	>��-[�6�m�	z�=JW[̇��޲��x����I�@�d��|=�ԖP�(�QZ;I6;�ڇ�˼21`,�����S�${j��f����\2���S�a|���߶&e��:����/ �
$�"UkZ���+qn�m���_}�k��%�?�ݗTY-:Zӗ�M�tݥ��6��×���_zUS�舛Z|R* 6D��-��0�r�|l"'�D>�Sd�J $����,��9���e�8{[�Vӑ�z],ٲ#�