��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*�s��W����*��%3R8x�l�a[��_oS�3���
�hfAX�A��gF�k$N!�_>�Ł�����ߊ� 5"}
���I�L�VB�y�(�hf灭X�l���q��c1[i��Pa"LG0K?7�<���5��F��nuӰk�X;^/�]q04xj��W��<n��D�`�j�"^���Q�̐���-v��Z������r���t�J�jK@<��n3q����9���˰���!P�> ��D����Ҋ�p����6��ryP0���K�˭]����8n�N��)�[��Qⶺ�TO:d�s�o��e$�H�����3�Y^�r����Bxi�Q����BY���F���Ra�vS�}���R#��zljKݿ?y^��v��k�{�ڀ��E(u�"� B�0��.�l��b�/�S뭦�:A,}>�N�I�:��ZO����]��<[	:_ԣ4��u;���vX�=?G�uǮ)&���
�1�.ƛP�?Ԏ`>��bl7k�zL����o�4V��� �g������
���;Z5X��؃,����)��5�(F����^�e�쌸Qܹ	�"��AvU���w���T���΁@ś�lg}�v����~n9��O�׎\�u���B�v��h6|獰��&�-����붓@m��T�H��'^q���S'�Fȹa�of�֋�G �M�k����X���p�dK��]%�,��BΗ�`�A�	�����ut�JU,�J������A�u	���.�9QR�t�POP�
�K�<��e1�nC�v��6n$�;q:Np�+��

n�>(���K�1������à����0:��u^!J�}[BH�C� jEL�����n#@T��]V~3(*�/�ѷ`���� Y� L���[�X� ��a���講)k� >":<B)Tg<_�Ȇ��0)�M��@e�J�J�{�w��{���߅���C�0z����4�([-��bws|�M}�N D�_�HI������F��\��\ �ǵi�����wd,'��j��-Q'JR�>%�����&L��0UJ� �H]_d��y�e0F`�oH�U�ć�?ge�'���
�h�����u]K�G��Ys�޽���ϓ�Ƙ6��iٹ	h:Ȧ�o4���c�3�m���x�$@��`t���3d�M���啸�_�f�J�{GB5�-�ۋ4���/_G���f��.��w��5Kn����f҆��t��A��v��S�9
&T���4-4~_�$X���d����oqH�A��IM�����X�_X�t�j��}�AԈ�X&�	W�c���R��R��̓Ӿ{{M�d ��b���2���߻�X D�����X~N����4�sj>���M�°2|ܬJȈb:�}�U�[�ּΙO�<6Cܕ�h��p��,#�lt�ZMv�k����;����ʱ2#BT������[���i�y
s{���9�=-�{�;u5���`�ùBv˿��	P��Z���"�:��ݍ�L@R��%E�bM��D\�pdmĕ�2��Y���Pcj�}���	�)	�1�v�'���o�/{�Y��EW�I��П�levlw����1�������S�Mv��|�~7���P�E�ts�p���z�"[�zg�l�gm�llhSFf���������w��~rsὠ\"$��"����Az����T:$��'�H�F�)��{�e�a�t���Ն���������u�[n��n3������{̦9��HF��󨻧�q�	��\��s9�l}��F��s_�3y��1ba4�Zl4���$��-Q%	W#��1
�2\bKH�e����P�d�D�;�<�g4�U����ǫ�VD�z�٫b�[��S��>�	;ܝ�h2R�ꐵ��q�\XE7;����8f��of	t��i��(]��=��=�D�A�2J"	�U�_��PRٌN�9��<�x�ܘ��^�U���%�r����!4NQ��$U�t/�%z��fP��2��f�\Sx���cR�"��^�E����7ANi3��#UM����w����6r��uG�;a"/Eoo�k�HR�@G;�����Z�{�kV)8)��!Q�ϹM*w���qAOp�@��F���X_��3����ܤ;t��S�1a�����~��l?���6Sс%�Og �h�й_����#���¸��~������Ic,ښd���C��f-)h�tܰ�e�����:x�,��9sڽ���r�.$j+o��<.e��
9.��i���E^����1�_xı�i$�}���fR�kn8��1��B����������=p"P47%�Q���s{�<J0<��aL᝙��;��)2���i�^�@n
7�K�ݖ>]ۭ���go���YD�K�0�G�}�����/[g3Im��+��o�R�r�[SP�cw����؂d��NqP�,�[OY���V��lG��K��X�w������Իs?�mso���y�6�:������:jCTT�*1?=�nt�^G��p�{��	��&_6�*e��7v���^������W�6$0lǷ��������
���dֈ6��ʊ��(�m���K�2־�{�3�HC�&���R\Y�0�tI3^ZS;�n�7U�,�JM��l�It%pcW桙�
K�<�^��tP��a�:��3�A6�H���ħ�s�LyW^��AQ����)>��<v�g7���T^.��q!ٸ���,b��u� �����"����rYۜ�����oS��J��H�B����3�S3i�j�:�R3��.�˿}1�sRa��J9�v�7&X_4�?�������q�4�#+�X�S�Y2�[�k���!γ��M�<ŉ�_UJ�D�F�afY�z�^H�,Wd�iA��+Q�E����9#�-o������M0A4˳����Y>d�Z���|��L���e����(���.uq(�y�I�@����{�x٪u�v�5��]�K�����
�w˹���:?���*]��k�ѷ��.�_�-3��ޖ�(��|��#[+��aJ�{0��<X��"���9 k�s�����tsd�R4P=�[G����k;��@|**݄���b��J����&o=2�p&��lH5�W�~b��}&�c'	�v��v�Bg@s�o1�ek3���W�O�Oy̳!�V�pk"�2>|��
d��MMdhֵ7�9T�v���+q�[0U��e<��ʊbox;��[�|�����*���z�l�pv!�FVI��BcǱ0��̕'cC�+�Ue��ܔ��Ǿ�
���E����k�=bN1X��x卧M��0��*��m��Ъk�����u��m��>��#�x1��,=p{�T��Qn�:�P�*"E���eO�[�t�.[�ټ�.���`�NL��Ƣc�E����]��·��t�]��kS
��i���F�&�R��0�q�g����[�^mc~������}y��2���P�v[,f�*Ȭ]�~��W,t>��⊰��#ϑ�m��9�]�}̯��M��ry`n�c�iT�SɬYu�#�va_��=�U�<7 �/����P��D���5��L֥m��A�]f:m(8��x8m���~s�&
��"ԗ��C�*2~�f\Z�����i1���(-Ow ~�5�Y֨VH�	D�~G�Ah���$U��Ϲٙ��y�X,?z���>��g4� r���|�~��� g�b�w܎���Ȕ�YI���?�nTey�>��<��B}xF�,ULr\k�Q[�
�!�������,g�������'���]c��M�P#ԬtH��8���Y�Z�fue�_1��u��A���NY����"�B�E6rF��-]G��P�$^�ir3�݋'2�2�9���wk�4�z8�c��y$K��aƶ$��Ѽ�|�m(*?�4��W?��t�*�
9�IĴS�LY�D� #͕~0�g8H�ű9��M�"70�D�_=={p��I�+���2�����&\�N�W��n��	}f-?���5�ԋ>��F�&�XDK?`q�u�����TZ8Դ�J/~�l�0'�C�lKi���n�-��Z�:�_����aZO;�LH�:�R(���^<%ۿ�����7:|`Z�Rc&3qc�ˏj"(ZNz7fс_���s���0A-rv�-� ����bA`�Ҁ5�[o��Ly�7������p�a_��J�T���������a41ZF����m]�JxO�՟E��I\��_?��EK��)fB4�<��W���M�'�Y4�4�_�CܰAvK穼F�~AQ�/s���ڷ�䭮�q&�Ch��x����������������<|_����*Fm�g�=�nJsE�ӆ{�RZ矪�2���%2�@� d�G
Z�Qޥ{���[���;f�1��Nws�e{l$=��c@��8���P�T��nyJ-F;�?Ŵ�p�YW ��m�\��X�V�	;'��>��ۏ���K�Tf7�����ͭ�Yk����%����b���5����k` �������6��A���H��\���ߏ*)��kń�t=�?{s�=�̉hZ9�f�Yb�_�¯�O��P������*^�{�[G���[\�
=EF�+Wb%� a�W�j��K��ot*�*�6,]\�W����h�?g6c�T�/�ٲ3-�`'�dG��lTI@��)�����2�E��:	OR�j��wkx|�������0�n��{�YgT��I�,η"����
M?�Z����3�!��CMe5X�P��H��Jq`�ԅ�QU���{�Q�m?���VY$U�v!�KQ2����&e@z�2���K�;���f̚�gn<�bM��	S<P� h�qy���%ܮ��w��N��Z�Z�]gsc�B��ļw���X�
"P��v�Z4�"Eع*�}�"֫lV�A��Dg�/i�F������Db��p5SYkb�2���Cɾ?wLK^|��	y �.,c�?�#�N��"��o�t���v�ocܘ�?�[�I�����^��3�w�4�vۢ�ΧgjE^w7�M,���r?v��5`oO{v��w�̨~A�e��
r�^?��p�m�I����6Tr��P e���g����P�N�]\��žį�-o�`�$<���$�}�<V
S�D��u0-Q+��t6�1���;�i喹��Q���yD�K��HȆ�EB�+��m��3rݺ��Zi����'�?��W���aCxs����)����	0�����t8�����Fj��ҙ���e�n9O���x���+8vۺ�n�*�d5D�v�=B<�=Qta�ߥ7�|�A�Ҿ
KV���qvR�����M�78fY*�}~�:�#���*!�?�x��Π�x`��R�F~Y��x���%�'ĳUl$ٚ���z�k�C[�K�]S�&�1��4�3Z��:3��C)��HY��V��/�"T�T���j��oB_c<�o�Vdp���� |����̎.�Q�$y@>��o��T��ʠ�וx&���K��P�|%��MI��֊��]0d��"2�/�0�S�k ��R
��O����If��җD~�5h�GqF�$~��S���x��<C��[��<pR��He� ���B�i�j�ʐ����f݊�)=�в%ol�U�wu�����-�.!�s�w	�nr����§���k���p��O���8d�^�V��t���W�R�m�䶡��濒 G}bZ��K0�Z�)�t=ᭉ~i�T�#b�ܲ�W ]�W�@��:r��
���&��5}�gL97`�'$�c�i$��['��[�2i�+�������EUs�gb$4���Ҳ	�IM?_\�h�\X�m0Y�˛�h�%�������}�uo�b��YX���N���T����0_�O�����Cg<I�'��=*l��(�
�xI=5�]�-ނ�
Gc|USĒ8�T���B��HX�(M̑���bM_N������YZ�B�f�%�N�Hwl�6���%T�Grp���G���/�:+S,v��_�D���J�N]��i�����mЮf��1)t�Y����Ҏ>�t�ߩf �ҏ>�+�I�#V
�'7�񻟞���l,p��$�o���*!��N"Ю��&f1b4�-�U�8��z��EQ����m_*E�; �c�l�<�X�.?4x�����/L�=�5
e��*�����$v"7���t_�����)-���!�-���Z~�߾e�m� .�����Ǆfn��2���~���	i�@��}���В��>�Ui�YO>���E�-t��g5\�(}�\_�@Z�>C̷�ബ�>n��?·1����Gb���%��w�Tb,��#vr6�ЁV�,u���aWk���L8���
b64%Q����R���˧�K�e��dhKvt*B ���%������Vkٗp���M�;�?�M
v"�Z3Ir�i�=G�23:����Fޞ���V��z��6VF�9����C'���_�Av�"�����\jADQM:��!�i+�X����nW6���Y�K�]�רY�#K*@��m r��k��t�^V�v������;tk*8&*`��v�Ӊ�f��u�{�s^AG��T��y�w��(9hIr����֋�lK��J]��Ȩ�a	ȕ�X�;`�)ա���	L�u�����)z���	V��2�b"�V^[ǿh���Йu9C�3tZ���*dA��'�y�.*v�V�N(�����PO��UZȥ0����4��>$� H>�g�7�~D�"�����"t�<BY�c�"���0$��'ѷ0��ZGԽ�D�U([�[t��
D��C�M_d����s����Y T� M�_��E�,^��< �Z���I��ІP[.����m�D�f�=�_\{�����:��e�x��ɋڥ��e#�aw��:X�����E^�m����v�GML��?�7Aӝ�_�x�7���/���9ؼ�3Vׇ��0��� ?'��G*�Y�Uoq%1��@�r��f�Õ�3�8�g� 2��j�54�o7\ïWpPP�r$���Ñ��	�\]�4�l�j��]��;��ͤf��Nڮ�9�4�[}�ST��8!.�JI����s@$<	;Sh�Gƴ���]
�ĉ�p���θT�{�6u�_����/�!^�����T���C�Ek�>.A��4�|-�/$�S�������TO��)��xi����Z�=��X�v��Ij`������D����9�v��I'
J{s���� __��	Mo	
�n@u@dV�5w���������LM��W�6�������]m�=+�r�d���τRwOo�����V���\8�٨.ܬ'8�;��5�� �i Ps�/�af�i�gw�+�?�mY��א�(�N��Hޱ�V�((vި��C
�tiT,��ɄkZ�6���e^�+D�:�xI��N�9� �d��K�qbZR�=q��Ŏ�E��SH?]U	�
͂T�#YfӸH!�l�m��S�ƨ� ���.�N;3_�����	�C�&����I�����W�������������å�q[�����E����.U����V�.��������~l�6F��C�������*�X��R/���Y����$(����R�B�cM�6>��O`X��ҵ��%��Z���=Qִ���M,pM�妙i��%)X���^ؙ"(!V�C�8���LV�&(l�WO@۝)um4B6�J��"���\b������9i-���x�"^ۘ��ϵ�Z_QΣ(�b˴6��8�!U2��=��]]�?[D������ ��a#� p���	?�i�v>5:�z%�7�S���3�/[�W:كl2����dK���x'�f.߹[ȏtF�h(\�7���2��mbי���6/
:Y^׽��gY�i��\1C���d ~VPwDg�Hn�������3���)�a�vLܝL���r�~NA2 2G:��t��]�<��طKT���Vq��ߓ^�~9�n�:í^2�-�PN� �%��L�d�R�v�ݸEch� ����g&��dm�ן�3nx��`�<:q0�FV�"/�H� j�X���=K���m��fB�o�S���U��
�P}LE��K�HQrn� �8������!�_ƌU����3�������B���������K���Ɩk$ra�H�"����\(\T��6�=���|q������5B���R�3�W�&��:�N�x�g��	M�T5$aT��q���<T�kvp����]]�פ��D|2���6��[ i�oE ���N�fvzg��Jr�d���/��^��0+9����J���a���ߍ!�z�1>���݂�B�l�"�X|uj���
�֜x����R�����v�皨�r.���'�<SgC��	��1�'�1
n�F�g���w��9'W�Ȟ�&�G��%;܊� Ï!6��yϯB��0ʀ��?:؉�g�^���6
�V���SQ��\������-�VV��E˸� ����P��Qj����x�H�
/��m����3*����.��c�щx��mT���3,���9�We�ŗ�b̞�^��^qs�H`[�uy0on�7Y�d������Ҧ��P�9_�ۃA���i'�|�7ȃ���i�C�9��>�-�Vπ�����b�'��/���͢l����B.yLLxI[u1���\�_$���P��,�m}�2 /^�'
@�yp��6��ʄrJ`11�nB{N9�����
j �c�_.1������$ ���Д���Sg{e�\��׏E��F���ܧ�$�|����]kJaƮ�d;Xc��|f�F{3
+�cT���߮t�� 6���Y+������O��"�B���)���!�t΀���?G��k#M�;�KKs6s���*��7S�����Ƙ7�sL2A��M��-[��K! X�,��f��M���ݭIYSTNh,A�V;8i~5��Fe=���8i�i�Xt^k���f)�-�<ϩ���zi}xmy"kّ����v.cj�F۱�k���UcApq����G��5��{"jm0g�/�.
H�f�r<2���������6�H���j-��#���8neڹ�	uX���;j�F� ����Q���Yce������"�v8P,�]n�_
(Q}�.�^��?�	;��������Vv��},φs�P_��n�_���w�*uTC�Х��4�?U~Ѣ�\ݨ	��i����dii'h�}c׈�Λ�qϾ��]���D�%ȷɄ�!�5���������h�_9� |��f�~$t��]�	P�٤/�s8�ME�Ot������kB�/:�u�0̎��6�0F�C?u;���X�Ķ����}S��V��ǰp�Cg�d��*K�MH�>�u|a2�	�Cy�������X��ϴ��f���o���|Y���e�J�׀����sn�v�������5l��$��3�zWj�t*�[��A �h.t~Lk��?=��$�p������Y	(��(^M��%���he4����ٻtOk�Z�`I��Z�
!���7�%l��
�|~�_��N����6=S1;��v��������hMi V�p��0�5Q5z��u4�5�t��:��5i�-`��0(XJ���Yإ46�\Nt;4�žƽ�L��~����, �Af�0�w&6N��Ⱦp�x�������9J}�Ns���<���ύ;s�~�yp�u�`���f�%�r6�3����÷@���͢�I�,��*���~B��N�v�����\���#5WzH�?���Uָ�9�WZ Fsv �imsK�'Lc��F��o����P���i,�sD,w��2bǮ�$5�|ج~����Çb���WL��]����]Uy����6��ja��~ʶ����;����ea�L�&�3����n��B�!Wj�n�CT\�D���r�
1��H��u�P��t�ll(Rf[�a����%*c�$7�CY�ދ��6�������K.O�z!�x�(���e�Ky�w2�=
�f�����\�K>��&�5��>{�h`42D���<c���o"O,�kT�7�_fmQ�RH�}��Q�VSq�*�������{F�Q�:�}>'�z��i<ylI���)f^��"��7�u=\V"@�2�ZXYY8ܶ�w7�u�E[\�������ֲҶ���	j��-����ɵХrK�38�Ÿ�����9�v>�1���Q����nv��k(�Ͱ'��d;����Q.�˞��	�#����؏O�	��T�WS����.In���n�+[�@��� ���'���Oy�V�8�mW�v��5y?����9QL�"4UF>�[n);(x�Ϊɤ�4��f 	:�8�_Ä{��LVU���dw@�%P_�`|�^�ϥ7.s��������L��顁^���Y��P�ԀL���c�m����p���V<C��:B�ŷ�����Iq�=�	�����flg��ܒ��Y�ʞ�*�I�y���vp&��ڻ��G!�ϧ�a�b�tFQ�דR3/o�6w�{�6e���A�� Y�����Q�V��t��N��빏�xoZSu��e";ѯIZf���|�����D���\��e���N���,u�v�J�����ۙ������hg ՘p}A�������z!ۿl]��P���[�u�(�3+tf�GM��	��l	�R�E7V��C��:���Ė�"�:��Z�G���8V�y��X �l��[))��+K)���!�/x瀚���?���Qqomzr�L2�$~1���<�T=�]+��Hh�r�g��I�:�j�{��q��`�ƇӔ�'�l���׵~��m|��s˶�9V��yW�������\����<��4����\�QF�J�1K�C��j/f��L�X$�~'i@���r�]��?�	�5����6�T�%�!P�G|��'�j�R��꛿����b2�]@�\�=�Q�U�{�s��*�H3ѪE�U9�E�����#�z��N
��v��p�RӹB�<z ,!��;����x�������8�Wy�|Y�\�	���3+�h�dh#���b��<�J���*iyQ�]%b�	�/6���Uګ�+-��C���j�2ƍg�4BL��X�ԙ�k�ޏ2��r��ەP/�pt�������>K�� "���k^Lx5�����ǚ�V>�M��
8�b�>�Eሬ.�w�דA9�x�ߘ�2H�J>R�2�1O�Bs�e�t�b����X���F���+w�	 g�4N\]l�A6�ƘaӚ���*��	�1`�ڐ�C�(m����L%��a5"<����6Y��%==���;U�jX�&�\�RpJu�&H{�
G5qj+��`�jS���U���%�n\���8v�9^ߞ0&���ˈ�Iu��[��!O"^&ES?/J`�ƀ���w=9�ݕ!��ȅmu�C��dG��#�$��y�蜀�ch�0���%&'����+��D��qo�$�����D'��*ݞd��v��D4=�_q}n�jbr;q=����)ֳŰ�[���2A�B7S��]�.uqyg�2�&/4o�#Δ�����r�8M4�[� �y�m�٨҉1B�-�d3���Oh��o��b��T\G�МN���K���Sv3h�����#�C�'ې�l�u��|3�B�ѿ���q�o�F[y<h��Rr���kM������f��L��q��Q�9��à ���}�Yb�aQ��_]լ�Z�da�
G݅��+\��Ѭ5\�(�P)�&��HR�����i����������D��dkzOt�SO���ي�qF䢫D���kk{�íj�L_�l�Wⷛ�.��/;y��<��!����_+KE� ���N��C�Ң�+[C@��D�anCҧ��q�v�>R+��K�f~�>']��q�	 �)�Ƕնx�k�]����B�x)$X���jSW�X�$�bd�Ӆ�7���O4��XW���=����d�b�#3�
��v�U
�^��P���ev�I�eڒV��Y��R�����;��<�y�G#K�%�	%xQ4/�7�-Ҥ�K��E��"	�/d�ɞoEdg��XƢ��@��ƴD����}i|m`4ǔ1p�R.������c(��[�ag�J{0�ϋ�?����R<Ԍ�8H�;����7�Km�<�O�V�_I�i�/�%nj�Y�4��k#����y�.�-��n<ZE���󊵳bf ���|ѹ%� .��i�$�6�"�.	N�?>�0�=��֐2���5`�[����W���7;)��Lf�H����Q޶R}���}�qLka_^W��փ��� Ayu��2�\��s�X�k����s��5�rU��V~Veo59�w ��,y�]�����5�3��YZ���N��إ�HIsR��V���g?8/�E#��O���k̶���~ ��8|d�#ps�.�v�q�!����d��!t]�~oƣ�s-Ze�%Og!��'����IWN*u���#L��$���^5�A9x�G��zȝ�p`����չ�	��qM���SR [�z�`��C����?�vW��Y�Y�k8���_M>{%�	��Y��V�d���=]��9r�cO֯r�}Ⰹ�(�Ð�	�愄ȥ��Dwس�D����fu�D�L���m �J	�O��2�X�Ap���8��L�=v�����Ar�X�p�C��}�"��7�h:�����i�w��P��MW���h:���.&qߥ�##\r���@����/X���8�v����a^d�A��H:�?���o�d�tA�Q*�[[f�3O����ͽ��������5�Y8��)�O������]��w���"�Eq�P�<5�B=�{����%\�֝(��ǡ�"�K�)��L���_�����+M9�A^���zb*��*�|����E�5�5�_�st���>j%�U�J�q�Pv�����b�5',ƹCk���-���&�s%:�ϖMqN�ZOaJ)�/>;GV����3����l���h-����5�ʖ��O3A���W�CB�zO��Ď����K�=6�Se�[P")Q�\`Ǩ$J٫��6$xJ`ο��zٌ��I���,�&�q
�T́i*bt?�3.93��!�|��r����8�'�▮Ԃ.�e�vJ}r�@����fI�WFAvGH�f^�eNlLSƏ��-)�K�Py���U�����B�-ls]x�c_��~8�i��bʳqU�U߼$*�]���;;j#��8���<�¡���
%�s����w=F���֦˫��aj��B���TV����?4�x_W����^�l���;{��^b��&Sy~ɳ����Vd64�'܀�i���.֓dB'>-�;鸫|a�'"��Í�1�ˊ����{2f����:�#�2���{�҉^��}.(�D�$���A[�����B��;4���b�3v�X� �B9�b�lO��Y��`���H��P��9��kԉ="�T�<���Ŕ�A�)W#��0v��.<aiۓ|�%���<��{-(̺�[��6�j�Ƒ�X�����9M.��8��H%@-�^��\܎-�O�/=FZ^���*E��&���"$
wN1��f�|HE�4U6i�@�`G��j���~�c�gx��HB�c�Ele�H��z�6�6t2��8r1��,�G�dX�dh����;ZF��IV��%�j쐆df�3K�cR�
w�R߇��=	�,P�-��(d�.�b�͙��"���]���S�!r����W�ߜ������}��cev���@8�R�$���ݶ����bSx�WBz����	�,J���9T<�7�;��~���|�;n*}`�Mr��ȴ��+V��sYi0�2�����kΆ�.{P68(�S��Í���Y_��?�-�n�V�~$����s	}�\�����/Z�W�2W� HR���$F��"m:��_�d���^��Zz��%X=pR�J�Q��\���_��������\)��R�h�i�CJ��l��B]�#YV�I����// c�ʛT�����f��n$"��ó�і�@|u��Ez�,�që�z�m,��ZH�m�vo�(a�a}��I�(�z6�	 Q���W��l�{:�x��W�@,������j�O��7Ty���V>�.?�gR���:��wẚ'Z�|ۢۖ�G3pT�Uu�IFܼ���neΟMu�M���~y�"��4Ԩ��8�*k����o��i$M�=�UW%g�R�7o�A�@q��ehx�����Ƽݧ��X�a��B��ZC��L@��ɵ��d�Xi=�a~cZ�P�a���V[z��s�T��A��s]J��+a��������V�yָ%�[��A1�HTP�:I�I��cFn�<��8g͉��v@(�?t�}����ܠ��?u���g��RY|f!'�K�%'�]`>*����(��#�b�0d�����,�+�㶏Ž�L�94П�ᵃ��J
��q��J���Tz�V���ěF��y���~���/}!��չ��ݐ0�4he��ZXV�k���x]z/*���BL�nۊ�>ZDX����y��9���;UL�x��]�v�b[b�E������/�S&��A@؍��G���t���B�RC�ec0wL+�����~���g��7=o�w�=�LA��t���&&G�ٽSfX�y�l`7X?����p��P��jPnd������#�����emJ-˿D�-�1�:k3�x��j�]H>�����q���2��P��L���k� ����SƎ}�2���l�qjB�/i�7�!�%��VL�S���(.a�Hdo�؉�H�MubkgZ���ou5D�]K�:�sb�}�e���EyY	�r�a�+�0�#"=�G��F��
��/��lN��o"�}��Dn&�DPH3!ΙC򎙠�ytn�����JO�?}��y|���c���4���z��@�U�6�s%/$��Px�8�� Z?����^%���E.��Ɓ����q*������G�����&��NZx?�|�b�L��S��X��X����� �RaY �
|;<���=���b��v⏜�� D�`�"�-�w�[h�N���q���ݰ�]��}��d.\jP�Kq�%(,tZ��|(0�Q��0T��YI���P��,` X�Tr�y���ed��#g�ezn]�ih��օ$��M�q�<��DN�a��jl�Wp��&g�@�̌r�T�w*��-ˣ�N��+m��y������uЬ/%a=%wm�~�EV.I���M�c��~[j���y�B,�X�"�E�)�y���z}^
�6 ]�7V�a��O����_��2��a�G�Q+�?1�AŪ.]_(�	���l���QE즇e��WR����E°�K�i/�Ξ��;K�3)ƭ�Cށn� ��v��6��%�o���3����;���{�T�������9��PE�D�����t���eW�*N��p(�>����Ӆ8�r����i��Ns�	4������`B��rF<���2��K��x�fN��7���$ĳ$��H�h��H��<�~s��M�ct*Q��nm�)#)�}ř!5��7h@���w[��5�Ii^b�G�É�ֻ�#�>z�	��0�������U���4q��pF�A,1�j�v���+�?E���=ml�xX���o x'��h�
>[�ᑭ��U������.p�?�D���;B�BkT��?����'	��sI�:�V��LX���DN����gZ�:`�Ą^4ǝ��@[��`���,C�T�h�?����7>�u�#��Ӣm7��J��G@��ò��ȋ��1�,�
��G�����3S��Ľ�jĮ�N8S�?<��v�cV�Z,A�7��P�2�J�B����}g<Pˊ�E��kX�����ї���K���^���,h�*+�O�a�[3D��K��!�_�'�������\�ڳ��I�L�L�28B�p�H(O�ħ4t�4l��O·^�{�>��,�OtD��<HI��s���K{��U�':�����˴�Fr��_82��Ko|I^�����gۮ�iq"t9\��U�t� �I��0xG0�^/�8ä����-��<V�͖{M(��9���Y��d��R�&��o��`� ���K�����;��#K���?�P����um9j�M��
%P&�!A**�vN&��G
�d��d�����æF2� f)�i��)g[�W�@���Wv��c՘��$M��#c�- �|�_�D��@��r���	��������Bϡ�������p����^���/X�x��1�4���L"�>�+M��h����ܳ����T�������o�t�"-��M6�i��u�l��� �
�[�8��yB����?�sad藅LJ�-�gQ t����p�R�!�P�N�r����m ������Dzj%�+�4
nW{#P/�dJ#�+ث��$3N��Pz��%�.�n��V������1�QbN32���n˯�P�"a�C�`AxqN�\'3 �
������H|�E~h���RWR��/юec�ܩ-?�U%��;&1$��5��\�I��˽�F&���Z���**���TZ��b�Mr����MY6F��X-~�X�&�ǅ��A,@�q;#�
�e��������+>�40���[�oQ�+���w7�6ĵ`���H�V��� �I��W���G����e��n����^�v�=�ʩ5�/?4U;iZ^[1禵<����q��7Wn�$��L%ۅ�q��锶Шb���-'�I�u�C�5}���\���%;���`�Z�����c7=$X�x��4{���t](����>�[h3�	�*�Ј�3K�y׊���r{a
׎#�]�����X�,�	Y	�&����P�D������5@|���ڛ�(��X48)������b)/��V��ĉ�Pkc��F�:X�B�M�&�dKw�KlY�I4��ɿ+�I~6�ٵ�sѭ��H�� j���T��^J��'6��u���\oA�����H�̾���\�V����u,��~DjXE{��#�1V~�!a��'��q|,��@E����F��De��GO�mO�a�W!��9b��P�I���#�z8��Ma���Y(�N5	�����I�����/�v��K.̳��RiB�.���t/�B�?��)7y_^!!�1T޹S�(�JFZ�nk�U��{A1�iׂZ�ۊ��@�g�]�yy�����'������_�6d�XOc���9]��%�	G��R�!��K@���5R.�_<|Y����$�b�N��mAZ\�M���Ρ�W?rN��w�M+��=�B-��F��ޡ7e�1�w��-��ťl�.0KQ�=�Q%�L���:#�H���T�b+�pr�/k�=Dk��żjW�t�a7\��	63&��sP�1�)�	�\7 ��B�z���`@�8���O�5�9;�ш؇M��Y���H���:�����ԭ�\%Gp��Z���n��}�P:�n�0w&ҵw�t�}��H:^���Y��Rh5|B��t0$l|�
aj <KY5R'=9�������r�b<����w�R��Me����`���4�>�S���h���yV���ᖰ��*v�n�A�?r�ӱ^&���q.����&@��-D��y����L�̨@H��V?Π�hZm]�F��wL4zU��V�pM�u��ٌkbX�U�MKFqό�(f�>�g9F��6��Ԑ�^�ph%]�E,����Pq�A=�.f"��\��|�4�$s��k�}eh]E{�
Y�Dl���3N��]֜�{���x)���(��n�`�m��*��4���H�z`U*�P&ؿ�@��S�&N�<!t�B+��Q�\����7Q��Ay>�M�:������.��BG�$����P*�Z �8���1m3n㯙X9k���|�)��z����`ĝA���A)��;s��x2T�AI�J�o1'K �v�}����l�&���>����b���lC궆��2筅li�v�vt����	8�-�@�q�`$:p0L�Rv���1 ��YeK$���
��k
��E܏
i${���m������8��C���mH�[m�HPr��0����,F��"��ē֙��"�
�
�d��a[����>��LK�]<Y��Ĭ
��t�����|�c`�Q�{��^#-r��M���9���@�[�B!�'�,x���r6!R󃙯,qe�����p��Y��Z���;ZX�1pJ�q��/G�)!����{�����Z�)�̵�$�Y�����N����duߖݳ �7�4�����8,V�r�*l �q	�Z<7�D3���r~���;�:=����d�H�sM���q��(�v���ջe^HrsnA�,�oY�qߩ?<�!�Ua?�.��n�y��t�����Q(��&q�M�������k�-�L�E+tц���m^d/��j+ߵQ\%}�q�� y
\��ڻb�B����)Si�<˺/�Sɣ��b��c����}9��8y��*����sՇ��n7eZ�*9f�?� �1���� Q�k�tR^Y*��a|�G���(���e��!�LQ�v���U-l"����;���������Dz�!�hf�i��GQ�,��3�_���,۳X�H����hf&�؆�iPd����������<ݛ������% 2V#��l�]WDp��%e*��و�n-j=�AS ��-����{tx���V��$�n� '��~k�1g�w��f��K�ZL�i��F*���h�qT�}���+�g���?0Մ�W��FN%���J]��D�\�7�%o� ¹��)�N@Ƶ���z��>9νj�&x2������f�m�N6���ɇ�'�H=���?�t�������y�������/����qS�IkJ���+�	j7�v�q�u�]�p��O{B�X}hwMrq@�Ķ�J�P�n<T*L�6@	_@���i����w ΀��ώ���g�`�K�ßxV�Vt)?OOu��O�(K�5����x��[F�FD�ϊ9�	CN�	2��G��i[���a��ګD��x��-e���^Spm�@�E�ǰ��ьñ�018�w��� l�V_��4��&���:?�/�5�K/�bNDaBz1��~��
�k!�K��,�V*P����ld� H�/_���<fe1�S��ʡ�°X�XBC�~�E'1�E�*�`[�C.c��~J���9_]{l���ڕ��*Fi��S�At�p��q:�C0乗�ٱ��4��^�|��h�b�ٔ$�hy�+�Gx�)�߯3Ս�{����qc!�FU�~ǅC���c��v���yҮ��!7�3�/��S�(�_K�f˳(i��@����'u]�JT.����{��<����Z����.^��I*�
�%ڙԩױ(�#f�L�H�M��z$M���+߹�_?�{�}�;�R�c��6��AC������aq�,]�<��-����ռ�;��R?����j����b���z�Ey��fx�:$��HE���|��geX��P4E88	:�5)�N<"�_���D:y�������[B?{�I���]�7�^�m#�O�Mܡ3jq�<���_�xV~�k���� JU��4�����.^[m�0�oj]���O�΁�9/i�x�˱o�L/ex̉���/��ݜe��Ǹ���%��Xa����:Pi�`���"��c�`і�;0�^��S�ﯪ�� ��H�l*4��G��p�lV�']	39�3&�K2ޟ�a?��N�ذL�c�n��AS �N"����aW6��A��+C����Q���=�3k1��F
�*�p��G<	��~5H���5����.Ш�v�R�F�fV�
�{���k�l�2��Kۏ�묔��i/��JJ\�I��pH����n�G"x��aA G�,��:�����
�G���#hh�q`늃 �vj%Hz�S��N�yٻX�X��e�	�HB$�M"�����r��+^���3��}-6�|�wr)Z↿J��� b���8�F\�m���  0�V�qf?�0�d�;�T���.���jz�0��������J(�8g�xz^5����u���Z�w�jR�\�z��N/ �Kx}!BEwݥ�<������T��#�i�o�bV'���^���x4*������C*�:��S��Y�!(>j���ig�Q���d-�Q=T]�}j�/`%i� 7�e��y3���ru��t@ڧ��.{�NH:ĖfJ� I�jma ��Ht{�fh�vA)��xNYy~�� ���v�>&>U�h�w��>��i���<�w0$�bZO�EϷQIX��Y;jㅒh-��$����H���lʁ��koF�6��8Sh�˫am$�fܞ�X�)��-�L���t��Wv���rLa��|��t?s	�������%�"ܸ��>�)v/�7�����j1� �e�1���~ie2D�����x�S�(n+�7�O�`�q�= ?,�����7V�~4��Z"�� i*ȟ�14���w���g?�'�Z��p��SD��~�f�օ~�6l8{�9ج�[Ɖ�k�h������S��U�cT{�]b�bu^��j/]��`)����&�XQ#\��v�!��J>2Y	���V�K���<��*	�g���HW��#DH�Ulq#�	z�n��S{�`yp���]%v�FYW���p�i����9=̭��dT�S͵�]=����P�bBr��j��i݌�$�9z�	)#�����R���lݻDW��^y�[p뿫@\���q�[9o��r�,�o�9\��0bޑ�\�iĠ��O+r�{oK��Q
�a����<���-r7)7��n��QH�c��v
��X���;����]qկ4�s����MDn�3ɐ�B���T �bq7ik�<�ǂ^u}�#O�p?�<�(W�~�-�����J���W�Xz�\��Rh�&�}m��T��B^t�/���nVB��_ژM����a��K4����h��Z��J�ȣ/X�u����-9��ށ�Wط���$�[�־O�c"�O򗀫����Κ[=�XK�|�
Yk|�T������|�Q
P]c#���Ou3�Q4~ �1*Ҏ����a3tA$$g 5a�f��3�PPR
�'A�N�	f���x�Aw3��6���jj�·�TV��la����F�\�&5�tjIs��[�|��Y=%K@��.�b��%�����	�64�h�Q0��^�6�����Q)�͖' �'��2��,!�B�P}�v�����*��<�Ճ{�����0�	���F�D4R �1�0R���ӵ�����O�)s+�D:Gx�.��V���g׆���;g��J�+�	�'ߑ�>?HB�6�1�[�����G��93�����|������G۴6���/H<6�(y�0"���M�asf�u�5z�j�� 3k:�^�S�a<����˟9��-'��Q���o���piyԭ[Ȫ �=r����K��t{7Z� f\+~2H`����������+��C&�}��0m%0��mo�~��j�K�#�\c�B���N5�f"Ώ�}g�����sն�Q�D�2X�5���#��#_�~l������"MT���nL���r����.ֽ��R��b���]I�-i�o�$)�Q ��8���z6[�{��:S��R�̒�I��(F�� g~�g=��*�˖;Y�C;2p͊�z�� _v0�����L9�%��}�X3�~Bf@d9��ފƋ��N�_��v�j����H;�xp%��3F�3����a��4w�b>��!n�A�Jw �#�U�m�'��H��F�C%l��E�aV��&���?���8�4�y.!f�6�$��;��H�9�M�A�k��%����>%��lۚ�+��$��e�2Y�G�1.j�ʋA�t4W&���iv�R��8W��1"�� uX����1�#��ogo���JF.�l�r��?�f��(�i�@�z���WJ�2;���6��n®��PmÀ���6�����5(=�Ki8�`�&W5�/���j��K|�DU�ma�q�T�oUlabl�1o�؜��"��w2�jbg.'l�9�ޜqB��j7a��4j��bC P�b�Rp/5>�]*��K�0�Ӄ�n�����L���;S�fʻ����i�`s8��Ss�T�T�Ȉ��<Hg"ݫx�mqs�&���a��_V�B�h��&��������N�k��F�}5�*m�^���<l'1�����̩,p�p�ŵ���� �W=`�\�9�u]��tG����*��