��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf�$!��k�� ��,�uT.|���Q�]���*B�pFz2Xt�t=�Y6��H�+���}f��s�4�2ܠ*�����#lo��f�27�������)�|���j`�9;�g��4G�_��T�������T�ػ������wט ��nwD�R�.�p��:�[�D.ۍ����5��eܻG3V���������xIeeZ_kc�2*>���u^M�����&�Xr��-w����)��c�<�b輵��3������� K���&���Y*�\eZ�����|+�M��PЗ��)�a�jI�k�5K`J���.Q2��	�ҵ+�4b��)T�G�')�?Ի&	"N$Z޿mu5ￊ:�|	��lA�X����vLJ�J��~:d�pn�D��-ȁ ��
f��%\r���5�^��ז*w[�h����ߔ���^޿�dR>��V���d ��1>�6��q�~��U��ϙm�x�D���W��.%W�d"��{s�ry�joO���p��b2o�b��C+�
� �_��9GK�QLE�Z�C8U���n艤G^�^HZ���	�KKc���w[7W;ϕ�7�q)��U����l�jF��Fm�0{����٣��=,���|��i`�!�5o�����ܒ�Q%�:~�F�5��ş��gQB����)��"�D��~���X�Y��S���"���l$s('��R�`�t^��N�C������l�lWW9S���N[����tܴ�͵8���k�xY�gf�d�%D�UG�1q���2��|B'�I�[tG�7$��#o\b��g��9[��ﮁwM��sw���/�;��t�I�O�&7��l��~]9}Ɋu�26�ظ����� _2h��H�n'��������s*B��\� �[s��S�2��7q� ��"�bx�Y��s��f4����A��`���*!.Ԑ v�X9����b��	�;G�0]���C��5+�.�垄�C���ٷ0��b ��^�����Q��u�fl�׺ƱK��i��q�^IC�kV��R�2Ǐݧ��p�ħәU&��ݟV~(Oa5|<�һT��>�Y��W�$���<���7%���V�\-�-��\�SWV$B͠�S`ϗ]@7�Yߦk�����V�	QE��|�Y<�5��[����\�*`d�V���K�S�h�"t�2���[8Y֍M����PRӧz��)�A�¨��'K�|2f����`�&���p��w�1$��&��%u�}���j�%U6i9Oa�2͢���8e4�X5f����5�"f��f	��I>9 "��/�+�ε��Jo��`�����~�^]�U,�T6�ݷ%Jy�y�@hIM��/����hH�Z��Vr����֫�I;�mA�U.����9~�pyv�#&���b�������K8{ո7��T�n����uFʶumb&��*� ��Ɖ��4HM�{T�qa��Ll�|�+%��Á�8���f0Τ��P��/Y�|,����h�	�z��V'odĊ���-��1k��G��T'�`��/^�|0 İ؝��z���e4�_�m�s��ՍS�Ӕ�4��x1y<����$ҫ�i��4�?0��.G�ե����E$(�Na7צũY'�#Ñ�K��;����;)��
�\f�7�ޱFF&|�O���.5qz0���UZ��B�f2��$�
r.�׳�n��pFAТ�#IX��J}��El�(c��9�O�+<PG5�٤�+e.�� ��^��@��4 G������f�#j2��,5�h4뫽(�^T�S�����h9Y0�+pn��S�r�����g��]�ϮϦ�ܑ�4G��5�����-��N�������L��ĩ������i4�E�ļ�� P�!0��>E�5H�<�1s�A�d�KFS�?��A��e�5 J��)��D�|]ں_�Y��NUѭ(��A�̍���	�?WK��QAXVE��9*%�D`Bք�