��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�j�uh� ��!��3{(E��;=N�LdoyC�`*0Z��-ut- �S2�"������(� ���( ����|=�kI��7ke&:�Mb����������7so���[��Nz��D�,�x��
:+lŦ��������EP�߯��q�-x�r��ц:�U����	$�i仾�=#q�+�d9��^(��&
p$���{�`!���6F���VB�lu�@��t&���/� c3ZkЕ�	}�L2�um��3��}@�*���Y4U.�Na��χ	�i�	`��=F�!�c��C�M�:����="�u�i<5$9g/.Zk�  Ќ�,ٜ)b�J���������A�y���-��YEP
��8Xq��-��)���T��oDX�
�!��t��(x�_�[-2�%��|M8��nzv��LvEe_���\Ԛ�3�%c��VF6s��J�Z~�=�w�s��^�VA�Zz{�<BfK����������1��C�i�����{$���������U���0��R��EiN}�0�0	�����j�c��4t,��ȗC7*R @T�QΙ�q�f���L���x���ǽ�}�Y^%� �}�(5�\�	���R��.W-5�ww�XT1�뉳=H���x��<A1�k���ln�)]���lH�n2g�<ÑY<�]z��7��s�R��.v,�o���UR%��M)��A�eEEeq�^ L��L��E g�/�?k�־��ٜ[���o�4���T]�_���4Rף\}�7�>b4�߆j�
$��fP �L�����b�'��qH�ru������#�&������X?&CK�i�$p�ݥ�c����Y��
c���d�6j(�@$c���8����i5��} "Q�|���M��"�ŷ�m��u3�*�9��l���Ib���	�-{�/PH«N��4GnXD;�����������*0�y�Ĵ���1�����=s\�n��G�"���1���'6,�}���b%�v�r���U�z�D��ٖAG.{V<��sv����v[�޶AH�܋�w�=3&��dI�Q���N�Q��9��	F~l�!m�D��2Mk�bP��j���j1j��� ˩�K�����{�p8� u�n:�Ҿk���W���i*���.qq��8T7	9��t�+�9�[i\��5'R�$���O��z�ؕX,���"垒kD�g,ٚ��^�g��T ˀƵg�Ȇ�.k�D�þ͈j7>� ���h���(>��B(p��nֺ�ǿ���^]� �m,�#p������ ����{t\����2�V�u��OU�i�3򥳬̮ -_�x8HƵ����è8-�l�������</��5�M��n�Y{Y�D��xo�N��b��4�l���ň�����X�%����S��6���f�	�V���e�8�%�p��w���9����}m���z��XU
�������d����b�i�&��+|<�E
a��e�xs&���s(=�$̹ob��3W�wL�J���뫗m`�B4W��%%���^�>����ʩ�j'�v������t�d����]��@�j�*����)�n���6_�D�R L��/���<ը�o�W����}�s�`�#O�+�~�h ;^���ǅ�7�Ô0u��(L��?��5���Vǧ�i�"eT���#:�5�3_/m
������*�q޼h���h@����.�αAD�ygO��~��*���?����ױ�|�@�Ҥ�=���"{2��?~��5����8FuM3�r��������#z/��#*��v3��T2�����a�f�N�>����aic�u�m(�ԧ颂i��'��(zg+��M��߈���2C�5���2�c8���tйRX�����D)'*�rf�e���}2� ��b�N���N�a�)�j�7��bKP��V��{��h����ơ��)^�sjo��]�V�Rk��~A5h�Ο=�q����{Bq�Q�7J*���k��� S��vM�S�ˇ�U��W�;�5��ܷ�c|��dN�nP��Ӌ����Q�/ы!���(�]a�ɾ_T1��5����jJ���s�L^gʻ-¥&� �f�_��%�r�ȏ㵫�tu�W�w���R�����m�;�V�:M��*2$���f>�.������q�LOr�1����ڂw�0������/���b=� D��i�왆��J��hu�{�#2���� �����4|^aF���x����x_k�=�9�֔����p�� ���Y�ٙA��gk]Ϝ���ʰ/���
�_D@-w1�.a�,ˠz��iU��
��}��=s}�tmo��tw-܌�g�BB�!.b+w��zqR�D�-r�\�Զ��d���06�1��63ۯ�-L&�%��l���1��e|��<:,O�F�A�Ĕ�4�]B���9��{[X���?G�6�ҷ�u����vs9/0��9un�a,��H�r�̑������hif~	(�3r����BuO��b�c;���@��}2f��_
b�w��?��)~
o3���%8U	�K��M�f�[��?�#M9�6��9���z�$�|��_��#��4�i�r�A3���t�7D��\�����;��Y�Ż�?{5����(m�t�b�1v����\�b�1JX�p�=a�b��^��oZ��SK�P��eB�~v-���a��Lx�x�v���NX�;�y3D��AۛH�T�O'���~��Z�=l�%ɇ�?�6*�ru2��1A}�9�о�i��#��~���Bv�7X{��#��l�g��Өa���������Ո&�f�v��O����y��Ě�������3)X��c ��O�=�qy��!�;fZ��6�^��2��`*��ͤ]k����&�Ç+��ȍ#W��h}�+���a<��[��\�A����W�����v�ؤ������'22~���@�K_	��=�·�T�ߟW�SU�jd�>��۸m��=k�O"�Oe�+�ȅy�@���Lѝ���1�˄rOE��x~T%i\>�j����s��������M�/Jb)w[X͡\Ia���0�n:um�YsMY�C�=���#z��8\K�C�~��d���Tڕ�?{QF�����[�
�?��m�� pQ��d���
�y��I�a���>>.~[)�?��Ѭ��{U��FK���ɤH�%x�eA@�2�t����{K��ǀ�{���������ְX�NѷÈ��P�s(�O��>�p\�
�-��F�|�;Ƒ��� 8�e��>?�Ze���ш*C������Y-���� ��6۪9^�ѿB*2���]���֒#20�XC�i}m����T�/=�ʃ����apv��zo%�U�Z�{��P�v��n�I����o�Fk����1ʸ��?�E�����]l`3�|]qu�N7�;�V���\bNz\V���,�]�
9z�Kx�$%���8,n$����a��ܹ�� 'M:K�jw���x��;�{��H���eK�8�۪#��|��r"��)����3�zn�Ř�v�zutz��0/RULR�2SH3[����6A��uU�s�1��,��U����>�?K/��
�S1�Ũ�@y�ю�8?d����2�q�fQ(z-�d�Vl�4�siC:_7b��:��~��ˏNǑ2�{��y|-c��k-L'(	�^��
����[i(!(���@�C�;J�s�y*d�/�Pd۫�Sr�V^Ӈ���:�SZ_�w��ef^�H�<�e�U\n[�E���2�v�D+}U	Ƣ�q``E�Y&����-3�&��>%���V�
�;?^x�қ�n`[M
�l��������&�a�"鵘8_ o3�_��3ǭ����a�x2�2mܟ�)���󩴖COr�n�]0o�^}"��A�Ȓ�y������,���+Z�)�^�莓����Jž~�E�����da�W�~�l��N��B.���� �Lk;nb�VD_D)�� BȆ��͆���w$�� ��Ͷ:n�"���E�ˏg,�X�\w�f��e$�L����ٲ�V���}���Q/s���D@ԡ#�-�l8�f���2��;L���Y�\T��dZ7��a>�V�@f��jmo�18"QV�Jo"i����$�dY��3��m���Fh���]D�jo�t�Ă�=��sϢ�m��F�}�䵜��?Q�[Ձ�0�?-d�Ll�1�c��E�?+�`D�6�O;�:�:ېi�צl;�^y�)$����M��W×0'��O]х�P��"4��A��.����ŀP(~�&����K8)ئ)��l���m�&P��"}�O��r��ϵ��q�����{U ���q�C9��G��IAu�,CZ���GJ���J�D��Ł��%x�-�G��yС���:i.���&��-�;��/U$^����(aILI�"�`4W��d�P�}1N���jұbN�8�MUǷ�~\u�|�)���c�1*v�ǰ����S U���Q�,<�+��<����}��`�g�F��5��s�=������SIxo�($�9,8��]Q(���М�+v'V�I����$|�v��86�1�/�ؙ+�xi?^^�d��lt]�7Ș�4��_��xpLe�=l
~���k��!��1��f	\��hU�[<�� ���3®���p]� 5R�E�� v����P�ZA�:����6}��
�Q�����cz�W�t��<�5i����p�3��j^O�!�BF�N�^{���Z.m'b�F>���D�x��e�}���㻍tx�a����'�h5}1q>������3<�Y�gn󕚁��t^,v<� V�2����cj��Tf@�t'��Q����,�^%����dZ����ܭl���(+	���w9�����w�fvl����8.}�<>ʼ��)h��\��8:Ͳ�ߗո�i��~�`�j��n$��	�DZ*�3՗'�GTX{��
�t#�Q�KBԎ+0�+����X�@� ����/��5df��8��^ ��S�+�cS�(J�j�<f�x=�E7RY��]`^d���ُ�V���VTJ��?��	�ʋ��@v:�PħҨ��,_x�Um�N��&���F�" �q�oW��NQ�3.��,g���Ef��-��F9�,��L([����vNH�8i�7�6"�K��~�ih���t,?�4��-~2z�/ʹ Ŧ`�{mԍ�����*��^�{�A"��QJ?$���{�T|�q�H�h��W�\����b�+0���6��P%������ �j��|km�D�b):�ĳ�w�98����d�,0 �c%�_U����"�X+W��'����@B���Z����x���1(��s�\e,F��ؗ��3q�z�����]��7���ʉ��t�#~��*3*�n�k{/�%+�.]�M*ˈX
����)��ZƑ��u ���E�@R$�	��L+ۙ��*�e�x�?�]�t���z���1/~&��^�������cY$.��/uH5(�.�~�ϰ�!�M�ѹ}
�����D�u�9Β�����=#)4ú��� p�t%������^o&�/���Io&���X��斢�7?�%�a�Z�3�����W�Q`��i���\]�l�K#Ko�������s���s�#���R�Fܜ�7Ù$�����/fW5�}f�����!�蔿a\���.x�LP��LS��-��؜�;��rQ�}+j�M�[�fBAؐl=+� ��׊��i��J�3APǒ�==�>�e�:�m�S�z���v�5V�7Hʌ����pw�3Q�3�`r��$R(�e�a?h8��BxG�<:@���� /H�����z�y��?��:�0��jb�|^�5��q��X+�u�K�ubک���hj�o�#�ƍJI�]iG�g�w�	�wК�0��)u�N=�6�RWi~����?ڶMwΰX`O�3��B�t�e*���BYO�7��d�wF	JEV�$#�ƚUF�86eMC)?N���u�̛�]�DH���No���g{k��**�ާ�
n�y*A�Т� '����J�D�6���d �i��	n'��yQ�.���i����{i�Q�go�]e|fČ�CW��9�~�.,�33*�|�$�F)�2z�|�K��e�6G�bbw�]5"�y؄�%��J ѷ�DL�W�rVp"���&7��g� �0���.d7�蔿�x�Tm��V�S_;a�Q]1
����:��a�!
�?�c�$�<pd}�y��C~\l���� z�r|� g�Z�M����>y��6��<��.Ew��oX�/�����L ��©��`�Ea�ʝ�JR��q�$j���b�$�� ���YFM�1���� �F�Y7QDG�|戲�>F��! �yoR@�f�a򞡄i�4�
H5�'W.��Hd�K1y�6b�����>y8�b�^B��8z���9�L���2\�W�T��D���BJ1 _y�3�l�HO1��mt��>��@�Rb�����>P�в=�Sͺu׎�uƒ���}����˽p{�K��Ɉo�p0m�c���|�"�g��l`��<�%�+�DŴ$<;�#��O�y�����W�s�����C�'<J&�nf�Ĝk����+�.��_PN�D�{M�O�����F���1SW�]���*�o�����5�|��%�|�V0p+����,%�e�K�;���I���h(�_�)K�M�ʼ�_s�8	��_�6���6�R���}��D� �C���OҟWA�'��1��rKiFt�����^�)Rh)z��p�4�޴���B����3+���F���f�
��Pi(5�̾�qC���v���W3��O��u��g���#��[N���C���$���J�� ��c�ta2�\����WZn#��aҾ�� -�5��k��6RUEzڏ��5��L4t|�+���Fn�x��?�<@�$b{+��������	�m2��fdjƸB|=G�j�t���ā8.ᾡ�pT��|C�)���e2�$M�4Ŋ��n�!#o����'oM�X�^:���jE�P1#�f�~��)E�WH	#=
U��\�}���:IG�E�36�$b��3?�<!;�tc�]��iW��"ʾn��n�4Ƭ������$dvb��(���>:�*�]'��j��Co��Dw����֔`BCe9<2��!*)�뗁��^H�S�$���I+"�G�P�R�wqNtAs,6x���*�1��=�s���s�l�c�|B��GY�GF*������FrA!��<4�V^8�כ�m��_����]oD�6
�"lDr�D�p!�f�ߵjt�����:��j4�,�̫�����iOV1>e��e����?q8P����Bkt���T���	����Z`�^�QQQ�0��/_n���fu6�n\C.��(��K��s���8vUw��NJ��7��xU�R�dj`DR�v��f��n��ä�t�Q����x�O� %l��Ca�a�k��$C��
rnӢ�a��R(�yx��;@U⊦���MuMZݽB�����i�����X�Y��Ï����-L( �+s�H���h6w�S��U�6�~!����L!���t��[�X���%�+�T��YY��m�hw^Ź{��U]��kju
E���)�*z5�uoRx����,��ϭiw�C.����%�@=ͽD��L=2��6ZE^�����f��uN��ÎJ�X��n�pO�[��"�j�1/��ڜ����76r���c�^�������ށP&y��a�`p�c//՗�e������F���Z��Jϰ����b&~��^���b���#'�����"]�0�@�A��K�/|�#���ٹ��!h�\�$s(�;�u� ��D�SD�|Ug��͡��~vKa�U�z�&���X{O�S?_��M�!��p/ ����{!��X��, U�6a?����-��jgu���Li�m^��ɏF��O�&���$`��\�i���Qnf������X\ֱ��9��\_p�$�g=P�<�2ܪj���`�A(��P㭘�MX沆��/�k�H ����ЎRB�U����&��FN]����1B��a��e�������SK���>����?.+�_�Y���e�Q@0��]�~G=�|��ޖ���#�)�s�EO��b���B���������|�U�p��)�d�1�W�]}$rP�yh����:�n ��_�8Į�$��a�+�� k�o��"M�]vO���UzO�˩7%�s7�ʑ�Y�@�'{}�|<�^k5�T�ץ�Z�7�f��Ԝ�mm/! ����¿!\f ��q����+/�.�_��Ht)�Ʋ4�X�
@�|��c,ď.�Z�n���&�tC�	��fk����݀�>j��e�=uf��B�$�;+,q�&�iߓ�>l��\�V�	9�0��"ҹ���Ť���C���y S[���u;N�0�6�vO�*"��#�k��f��,�_��
�v�LVn�M�݄�HT�l%4)D��
�\I y���hA�⒲�@�#�,�XF{64�Xو�q2��z2��uN���g���+�;���3c #G�����0U\�^ �_�j"m�B����fS�F����>�,;гpl+Oo���-�l����V�%f�$�'Ow�&c@e�A��qgm����͡t���Dab��rL*(Hd����?�w�I8֓[P� J}G�,3q��1|h8ۺ�fp<S�L���o�9\����r��&ة#��L�	�_�<�!�_�<.C�D�6"� ]h䉳����B�����\�`�q�:f�>��3����e�^�J7����@��}�Y*�q�#��*��P%����"9���Ƹ�����	��_n���;K��q�ˆ;v2�B�N�#�7�7}�����y+-��A~��s4�������Mw� [�h��ۑ�*��nC뮢T�_T�x�f�+�%�����S�"vsSG�ej��������c�ֹ��,��CD�{:������c�Y����J�T]P�������u�͂kZ`��N�1u��}�m���ĵL�������>EW��s~p���F��(��r��oӮ-��I�[��-�6�Vr�2~(�ߝ٣b/�g� o�:
'�mξ�]C�?-����ᚿD)���8zk�[�F�%�QcoI��e��|���]��S��{��n����u���)��0;~��i)��Y_"��u���R!02��5���/X,���{9"#�u�EI��7q $͚oyvQ�x�Z}�wո��dA���qdK����B��!"�M�P�ۧCJ���Q��������D"=���g������<�0��]Dt����eJҞ�Yds��MS�J�_��<TqW��>�|�.d�y>wԽ�S��6����˸Yw� #�p�v�p���J l���<���P�б�~5��!W�^���bmTq}4�~;�T,8|�e����jB�M����N*:�j�����x���8��-�'��k]�Sac�k�E*u����6�����qO�����w�ѩO�����3ʙ�:��J���	8B�U�
�<�=gΔ,�ln�P�3��|\��'��y��4�p���gb��b.��@Uߢ�jj�OV��ۊ���OCehaK[Vn��	-����5\�3�� ��;b�7)�`t� ӓ���%*�|"�k�DhƤ�7k�d�W����Є�`��)�)PF�j&�i�L�g��>�f��x����:O��dI �I\Rm�N,t����p�RO\I�|h��OTf��/��N���M0T�$	��V�`c�ō���2tF����U%������v6���3ܻ3�W
y�=E��2��&z-1���3�a�\f��?�K2�f\|jɀv�L
*�l3��{A�p[�k����U_��M�mc50k_q�#:�ۮ9>澫e^[m?�A���)��6ڱC�J5��f$��Ě]���*��h�0����/�Y��Am?f(i�r&΢KV��4 �2�q�m�D�Ԓt޻>�UQu$w�wR|�J�%�"��T��c%�*�K3^�v��i|�&���p�f�ؽ�ܘ,q��se�E����YO	�K�ѕ��ڟ�}�V����.|��.u�z��m�����/��L��I+ųC+=�m2#A�}e��g~�Qx��Zz��o&�:���Paj�,��n��CY�1�bW��c�+�q�!�jr�٘g�W	�L��(��3���.=�����`Ox'�w���ԯU����~�DA�w�+u/@����D�����vSXn��f,8�&V���f��|��+5����z�I��P�@T�D �SM u�n	�3��5Hk�32A����F�I�aC~,ָ�)��3�|:��������MRjZ؆A匈k�xAX`�5tfwi#�W���+[tY�3��4ж/��DMe:Xͅm�ʠ�DC�E�^<P�@R�$�)�m����163CC{���#���0���r�����(0�����7�dO�@�}�-K_h��$�B���`��q��+�V�����z�Ojn[���J�)�Pڡ��l|	z+x�Y6�m^�o�8+XFX�W�C�.��p�U2j���xA�l6҉�r~
WP���"�aV-M�ޥn�$N�QL����;���Y�s�����3V�l7@$�
���� �/��(�4�f	�d���yw�ĳ*��W:�ۊ�}���9��O�=xܰ�z`��ŢLӘN��J5+���<��g�z�)4ׯsM2�c~	#��z*N�������ҕ]pв���ӫ�=�$���8���e1(	�{J��2�h��]2/�:�w��K��g ���s���d ����,���M�^��o����`�����)��{������R?�(��;ݐH|Ĭ���X���ǳ;*?���B
ɩ�T���zOq�2J����a��#&�U�I3 p�_�E��ȮV����r9�6i:��������������*"�Q�AQ{ĒH)�X�P4��5�**����3`��y1�HЮ6eY\F߈.J�\�Sb^�#`���M~���
�"kS�>��C�������) �v�/6���]�J��p�T6\)�)H�f�7�,e&bH[CL������H�R�?�����������E��i�z��s��ŕ�*`)ñ�{���rb�1x�2��:�o61�,8r�X�����y�WFkM�=�$=AF�)�ͱ���ϋ��`X�i��8#fòێAfʚ�H5Y�ږX�/t�Bk��h1�Y3�&�V1{�G���Y��-��;����T;3U�g_4[�K�����h)/`���>6�)n�?�1�X\����#A��p�3�S���P�*Ⱥ��y�����d�6���or��Ĭ�1z˖l��\���i���ȉk÷�';rR�UH�I�Ċ>�M��*j~9!���(�dpoU���Il{��7vA2�AV�ss<������"0�L�ǳ�2�zVg�ިz	c�}�AS�OI�([L͔��ł�p9�v8㜁1-���i�GAu��F�[%�BChU�DFv�`;v�9Ox�����*@ tB����R|���ݲ�_$>R[|�{0�Y�<�xX�!�+�[`Y�9����k8u�؞�K7�hi'��R�Kb��y:���Q;�y�
�s��W��=�d�HS�n�I�}�Ml|t���f�/��,D�s�B�O��ˣ,��qlGͅ����&�������j"�q,�1�t6S����Yv� ���zA 09�2�4�]���ؘ]�3���ߝ��Dڶ���S�.�f�m�	*!�%F��>�do��+����[4�+���h���y��A,�k�Y�δT�6z��>i�B-�Mٶ��-���4_S�>ze������](�dX��9HgS�2��[�v��YL�;��!ay�A��d�S7_�G��!�xo�L���S�B
�"^����-p��I�CոZ���i�=�~��n�>����(��h��1�oOrT����ncj�.��QhS�;F)O������RP��'����
WS�/�=w��q�0��9d�θ���3��2�y$���m����Z�fX��̦��r�9ZEF��$�`��6a,H���U�gw�$�'Ҏ�&X��Q_I���DE�ojU=��x����!��:�����jn,R�wr� ��bk��آ�&���y����)����E�"�~B0�lꗾ,��Sh��jq:�1�=���Z+��� ���z�+�2�^�|�ӂWCyؙ��ʉ�a�����9O�������RKl�,-�ߪ�����fU�������}��c�Hv�c���S��Q�<c)�A"%o�*�Fe��Af�3����S�3'�g��D ������خP
��%����Z	��#�$c���$|f����7��=:�R�(X�R�&��n��>�o�p�����	����l0�t>�fr:+�J�w�?�{s����NMO�8�>ă�����%_�V���S1�P|�ސ�$���Sb=�j�-����76�k�c��LB�^��v�_Vf�U?�r�>g)uEf+v�wqz ����v<C�:���g�wO�y��{Y��7�(ۉ��u��W#�d�x_ ոo��̕��Ӑ@q��H)>�G���W�l��NC��(F�@�>�vB�q��>w����z(^��m6�9O�=-��@�;���@6�H�C�Nlnc�������DjI��_K�UF�"[*��@Q��~c�x���׼x���9��`4���ʋb��b�ԭ3���M6l7���|���H᰼�GԆ��9l�-7��r�S o��"h�y�c���������#���u�N��<+Ӈp��>&=���l�k�|��8�0�a6{����I%�=�2�3�u�4X?��?�r��}���N�+�l�U�bk:j)�I�T��=V�eԾˤߓ\_:�A��ڲF��R`^���Y�IH�*��D���.�tQ���
�s�
��fc׎s�k�N����5����T��p}�\���B9�I����W��ϋ��@���p���Uj�G�� �E���e���ԋ�����t��4�5I��\`_&0;ɾk@��%��YR eX8���Cq��y�j�x8��d��O��G��V�	���A$������8�˫�N����j��;_l(��%쒩<���jz�F�����uU eM��YC�~�|�P�j\)��(��Ѥ��r-�q魲�:�LR�N6��[R�zXd�~��7��"֛b�2�zR(v	�嗪3D�/�=Ĉ��3�����N�O�����!���`�����LEv�5S)N�PȞ��l��ΤA�����JZ���S�%ز�%�BI ���%f
wfhM\��tb�q�e��� K5�m���N�w�n�.�'kfp��,�����������j����F�dcΑB3��]�/�W�K���?+���֏}�&	�7p�$��c�_wU��ҭ�E�L&<��ų�������;۹�T��x>R���T <��H�ˋ�+	�	7�1	On)�_��Ldc	��x� /N�X�>��k����q}�#|�浚�5;��p��Q�¦�A��Dk���(sW63B�;oR�6 ����P�f}yγ�줭I�7ܕ�_)7����X�@���T`��{����q��U���!S��)2�,$Ys<J�goT�H�I�5J��q>K["��]e�(��Ѵ&~�P��w�Կm࠵�<,�'�̈e���G7����z��/��1��\�a�f��7�5z��ĕT.؏'�4�q���:���$����[�Mvj_��6Eړ�=9ѧS-&��,����h믈X�q+q�#1��C�0��	UT��p����Ђ�!���1:<^T<�H}�m�Ry��?���(!
]�`���* ���� ��rX
���U\����W	���J|��1Ӟ�o�乢O�!��1��=����Z�b��S���)sy!��x 6�,�;u*�r��N`�F@�)�v<��3�>��x��uƤn�q��=�T�|ߐ.~1�/*��2d��(�WΠ.+�bT�0qi�8n>�g[d��ż�ƍGD"%�s#	�G���X�ŠE�b ��Xf.6�Q`�؁��<ZJ�+%�s⚍T�r����$���:/�P��:�T�)��]|ǟ�ٯ5����:��Hǘ�g�,m_=y3H���[���R����<1Ic��{��� w���rk����3hpQ����$q�Jo�(R�'ڭ�zG���5�`h���t�(e����9L3�e�c���0���s]vz�d.�C�n�RV�b)3�M[ߙW:�# �R���W�#�|AI�X�|��>6 �`=TN���ѻ�m��$-�9ϥ<ob�yȑh
��M��1m��x���|�b�슻���.,��)ࡁ�G1�������~Rr�03�sWU��Ԇg20,R�6_]�J2>l���4w��G8Ie�&3Z�x���i����4�����C�ۜ���/����������	mi�M[n��Q���6��E*��u����Տ��K[ Ye���'���J����|��BseR���d-"_@���aulDXD±�YB!���p�e�pGo��5Kʃ�����!�j���B�M|���{BRt�L�W�n2��ڑ��jX���*^[�����u�$}RN�R�����)X;(Ԏ�l ~	!G)�E�)}ـyQ�� �)��sai5�2�"���ӣ�]\�c��W��/���������œ�V3��!z�&(�l_f�z��3�QG���CPTz-��
��]�pn�q�&=�*�@�Ь 6�ΐ��C�N|��%����Pkk6��<��$P�T��y�Ն��wrB¬�i	ɛ�ޯ7��S�ORK�Z���\7S�e�D�_����g��Skp��9����v�r��和���2�:�����~�8[K)��o���r�w�p�h�	�#p�	t�� ,�.�6Q�\G�~ƱJ�,AbA3���S\�4�9;�F_�X�Q`sCk=�������'�Eiv<|,-9�U6!;B(<"�I�T���ߙXpXX�9/�����n���$G#M�??B���3����WH@��N��H���u4b���䅺�^��	��3�>�4e̢ ����ۜڪ?f�\i�!k�-c� �_mx~ɝ��?ߪGa�d�Jp��㘣���dv'���8�Iq�yv�>�U��)�߽_F�b^�Q�Gu���+O����Q�$_Y:���+&�t��W���c`N�-���������	h��y`s���H��吞$t�s/�+:I��ۂk���<m���	撾N_�㿳��ޢ��AH����B���z���"'����*�o��ҫEnB�������_e��o�Ǽ�)?�-�����1��'5�ԪPj�i"x؄�hy&������i0�E��G���-�+�p�n8="��si�+=ј��$���6rD�P�i9~Yz�
��pb�gdyUI� ����o3�Ě�/O�pˣ�L�t�Jb ��J4�]I��:ȶ�š^�"i�~��U^&% k��u�Tӊ��[�iG8�5`���~c�z��c3�^�Q���N�� ә��`�y��9��O]�Jf_[�a:�uBH�w�@���{X��]����]k(�� ��4���Djl�~eFD��/ѧ�Cvu_ɽPK�O�u��:l��́����)V0m~sp��VoI*�[m��� %P�: P-�d�N>`#��#	a4��'<�]�G�I����Qd��дN̽�i�nL�Ǜ1�[WR�]�O��x��{5�L!^daD�x*���NV��΁�A
�����G�j� K�j�g�!Y�>�;b8E����	ZN�H�r��zKӷ5�����u��W�g<�&��mx��x�P�;v�=�G�|M��L��[���p֭*�Dɱ8X1Ku���AQP@-���hY4�9��ؘJI־��46� ��|HkR[i���F3G.<4~��W�U�c�`5������Qg%�Z�QثV��?�[���6W���qs��%�R�FW�v�H|����J���#����E�զbź8��4Dۓ���+�8*f�|	�+������
ֺy�	�Rc�#��BܭAs��
�e.V�g����R���֮��h��s�{`��å��6t���S���V�H��)˫��p*�D�{c��ӌ�ɠ&bH|�(�B�%,�
<p��' �ɣ��20�jsA� �2����N_�y�@7�����x�L5$g���/��>��Jh縸�����$����b�8zW�������{t��w��a6Z��g�U�/���PZ��Ȕ�<���(�?���-��v���8��c��M��%�;$�� �S���((B�r���{k���7���7P�8��=�J�ӻ�r�ї���P{�-�q�N�I� <Q�̋�"o��B�<%\��b����Z��l�	��ZyI�d�g򫶍�����Q�-�o2v�>����E2� �����\��K�MP�h�H,��[����,5G<n!)2�8�� ~�7K���~�/���@Q��E���ҩ��Q�,�N��Dc��3 �x⸒.C/�{޳�-�xw8��\K��X���u$7����+
(6����jD��crn�Nq��g��V.��� O���!=&X��1i���.��}�$�5	gwf�����!UO'&��
��U�uc��8�k�7�dZh$�+�qQ	��#�5�y��夌���g�����)�g[	������.����z�G~R./�l��ye��.�/eD����<T%E�$�Ƶ�
��#��e绉����d���t� ��]��z�U�/�k#MC�`���UC��ꝦS��g����%!:S�r\`�5�� �y��?�:Ij6�m&^��c�rW�U�8����|E�9��ifl�L:U�c�O��W%��ZT\6�Y6\̹����/��(����;�ь���Ĥ�T_�����:�{����`I�rg�H&��MLB��\��v�HV��u �g�H-��d#&��[J����C	�<G��6!�x"�$�P�a�A�&fu�p�\���p��4��_`��l�_�Y.�*$-��	����tu�?)WN�|��K|x�䑔^@��Y	`;s�)拊6{(߱p���W�#�HUZ�$�W^7}���:���ĩ��|h��j�l��dBh	��^������}&�ͧ7P�X���T��=)P�B}'�c�)���i�$�S��'X�<�2�<Ar��i̋贺x`D�`jĴR؞V����@�Ռ?�N���R5��"�e�,92�)��w�GQcQ>����][�(]/)6���l��=,İ�y=Vqv�@��q)��U{�Du-4�,��۽�����������C���/��*ۓ�?��ŋA�������ERu��I�=:��G�k]Қ/҂���J���Y-;e���F��-�������n���R'yZ�6��� ��?ᘅg!R��p	B��?��]�\��W�dc$��	��%�\����);a�^�F�@��/}�Y@}Br'� ��F�>!G��%VN��4�W�1�S���}��T��W3X\�#�L�_eD+&�ap(�Z��ĭ�3��Y$F*���	.��a�M��9�^1-zN|� ��F�����B��ꈦ�2	6��B#7����m`�*�=���v�v�#�<M$I��_p1V����(J�6)�(r�͒Lqd�߈��M�|��I��B����nQ>�x��ꖆ�L(�?��7�l�*�=�������?�I�]L���	~n�)�`�3A�0�/	7��7�,ρ�iL!F���(M�,
�}k3��m|.��3�T�tO�%���K�랪^��M��b�+��D���?瀊�	���N�o�}��D����{��)��y���� �G
|~���)Rh,�#B����d�0�ޗFS���?��z@w�~��İV�'�/�s�X)�Ù��J�r�C��� ��Z�C�?�Y����tr�[�icJ�q�D���&��fi���@� �£e%o_
S�`��Ɩ�0��;(�)�c�%N��R�2�d
jW�e���`��E�@��0h��:S�,]�G�eA=���n/u(�7#�� f�O#�Uץ���\�*�ɨ�1�����Ѳ����Q��j��i�ÈܒI��{���kw ��|��%4��־I�q�	Ot���k|�x�ߵ�`Ʀ�����n�s��ǐ�T H�ܞ�CE@X�	��JI�� aA�z�eT�(u+26��ߦ�d��9�!ϖ�w�ƣr-�Uw�1�Y{uѬ�C�`b�ń�/�8"6���{d䞾��;��C��v�(�'�G���³��bLO������"�J�����F���P\gEv-�s�8��U��@Lܟ�W����Nu*�o`��������=9^�����%j"�;�;�m7j�&.�~����j�)�^=w(Q_ڿ=�!����`��������̰�{��7��[����k\P5�1�H��7
��MVU3��x��Q\kAt��1>�<E����5Dh0W��5~)>ӟ�Z���?M;	����1�Y���(ۏ��ͷ��k[ݢ^����e3�7mV%&$E����W�K�����Z�O�(�w��C7��hف��z#�H_щ���P�X��;oH�^��Z�^>�C�*v�w����� be>=�C�T�~�&��r���+3K�c����'8��\eS�ރ���qi�=9���+oC�:�$ruO�nmn,Ъ9�J�A '�|2: .l��M��K�{X2 �f�������
���C��!Q���I�ye&_k$)�X�TUyy
7��ߋDl
?�+b[��&*�g���Ξ_Nr2�A��T`S�r��#��+A"��n���U��f2�� F|�<���3��:�8��
 ]�7o���[�M���O�`>��V����g����K���_���V�d\����r�U��y����'V���*X�>A�US�NRh�:��Ns���:�������������#�;$���X"����7�-}�̝
��@������-��{�OXyc.����es�Y��7;�TSN�w�f_6^��$���uџ���!�ŁlƸ&��6�&��Q���ӻ�:s����E���Ts�H��^iv��'k�kE�&�X�X| �O",�vF�\���Ld�Vd��3��پ�SI��P�Û�7d({!���P�T;��fs���J�+��
L��}�W��ez�Q�3D��z:�+��M͟��,N-���Ce�z��r[�4�v��6�s���0j��W5���[e�sB�.QŻ�tV-A���J�j<'%'�[n��S}����j�����hl�f9��u�xs̅X/�H�O�����ww����i������C)T����g3�3�����*���gS�'nt����w�{��o���UCyD��1*|�fC���.����J��"���y��l��vJEWt�n@������P����?X�l	Xޢ��i~��G�[��K�	�_:��I�k&�����*�ҶqW)QQ�uZ�g�2��v��ݧ��prN���K��Hd#)����qd���}��U�~����-�vA����&nA�ؘ\���T9~@Yd�Y��
�r��_`A/G?f�V���m�5�t2��]��?������O&�kH�l�=y�$'���-^sڑ;+�ُ��i��ņsw��)	�nd�*r9�'���Ro�#��DZ��6�C#�|a����F+���Q�ةQ(e�� a"T�Zc>�$�o���R���\8P<�9����wP��B�n m�I �v�
C>!=7�O��O�7ʚX14H�Y���Q�=D�RU�oÎ62>x|U�n`���"�B@�G��8VӅv��(z�=�=C@�γ���v?K�M�-�ݿ�,QH6�}����ZP�C����\�2��oM�l2Qg�8u�3�ș	U~�se���l.��&q�?#��y<*��:���a�Ъ~�ۜu�sc��%D�ؠk�m|>�q���,w�a;Rz0�u՗��hc���4�2ڱKG�ݺ+�..$�S���xj�{����[7���;4ɵ��Gb*	������4>~z2ď~�S�F�~�㶣�1��/.��z�X� D��������#�W��Uy�B;D`�`c���O0ժ�5�K 8,���*��󱝑�_+=�~��ӱ��޻�џ5�\`��8����N��/��L;�"��M���b�셴@c4��`&�g�Xs����o�;�0!C]}U,�R����u����o�-�)���8=�@^�W�yj��TUIh��df��Z�c��R
��9ׄcDǰ��4��Q$�q�7QWj��k��K�Y�����H�#���(+7f3B�÷1+�0h����4���#r;X�B��o�g�8�≋�M���$��o~g�cK�m���}�A}��\}Zp�,#�D^!�x
��j��נN�LL�T���,��H�e{2����Q�����h��c8ު�����?4��;�W���{�F��1��,$J{P�?��˿���<�{�n���t�C$�[������|e�d�$3f��g�X(��?7�k����(ND�/�no�%D�v�ξW��$]s׈d�xTp�+�*���Ie%�]����YMC7VO�m�f �v��.H�5���<�%������y��7T����^(p�����%��0�dU�)�a�g��M���XR�8T�o>�hA���%]�� �p:+5��m|W'���H���H#<*�ݭ��o|�P��f���و���{/I��d%�D�Ay�J���j�UB��������$�@ɝ�����ڡ��o��rNǾ?�V�L�ia���(�Y�}\+�� ymp�����j>�6���o!��Y����_ު2*]�4�c?r!}`���`�2�|%����55�Re�J9v9��W�H*���}Ao������W	����>~|�|���$�o�7�"����#+?�2�pI̲�f�&|����!Mq����Y�>X�#�D�}#��1y-ӪUgٺ`��{E�>7�H�hr�N�l7?z��!�I�:��@��=(T���.?�n&Gag����w���?﷧�#/��Ƭk�f��,�������(zA#4-�,�� Բ�JчGW�Y��������9!��d��$=��"[��2�1���~��Z��;�cR��˴��;$�.Ś�VO��R����X���E?=���G�,K�ܲ�k�aTE" � �My����GK~�#�Y��L�5�y6�B%K�6��{q�~���h�없�Z�Q���$՝׆g2<�! zf\�;��K�	�ۯ�e �Gٺ��0-+�g-O$�6Hoj�_��:�$8�z����P�����|��v���a~�A����)D�Χ�b�y��V��۶޹<�)k���7j[i����\��l�S%�4A��V�$�2��`��xCr{�u%) ��xމ��꘨U_�mhH��ɉ$����K������'���V̵ť���1>q�\�D;�+0����#����0��a�^�Kutĝ����߯.^�������pMg3�PT�����}iGp�_ 2����?���T��d���x���)�Rc?�ҧ�����z�Xe�k���L��Un�Ҋ�մ�dM�ĵ�N*&y� =z�f�&O�o�ܲ��5Q�%�;Q�˹��74�5?M��=�L��ef���ڵ�İ��f��B�X���(8G����)��QWfA�P�HQ1�a��5؜��5h�v[��B���V{O-V��>I"`�ǣ1�,l�~��W��h�t�Fʷ���K{�����Q�v��X�nڴ�J�f����!���Nm�2�K

X�K�b@ݢf� �� [�I��R�_����0$%\��jۣ+���.ew��L)�����o�_�8�ڰ���o��-*��2��ƌ���Hߚ�0�i��ZE�M{a7��ma8Wp}l��I���=�q�;���j�$f�%v�u��26pP8}]s��t�ڛ.�����z}��|h,����6w��J/���}oo����E���^o~87�i�F��eZ�����;E����}g@�@�zn������DJ|�Tf�p~�Է���]+����Čc�ʓ&J�q�H�� �.�̼PAL���[*;���0���I���R�i���>�� ����4��u�lt@>ʷ��ͤO�=eQi�i�!Mp�ė�+�����T�����YIG����=D'�t�W�g���?�覻d1ז����^03�g��35��,z�䠥��=0I��s(�t�j��ί᪭T�:N�-p�ua˲��&I��L���dS���HІ�sG���{m�佘Ԕ>]�?@n�j�N�s�g�֞�Y�8R��H�E.G��迷�!f	Ij�����Q����Z��{ˈ`����dtzJ���Ss1���ݣ���O�92)��`�"aEropjj�J�U�Nk���\;w�w`�yءc���-TL@>���Ҟ���q��nar*C�C]�.�=3i�=��93��M��,Ƶ��Φh,O�G�	�Q�Q�hNf[�q:}��b!mfk�˔1��`�����g㎡��,#5!��Rj\q��q@RI�Y��j����.1�U��髩T(�3��Y������>�1�"�}���vB"���Q����u��,4��O�s����ٞ+$�6	��PE��`��e��Zpv�BHҞ�s���|�5e�4�
 <��CP5-r����T�d��SV��v���'b.�o ���%vJ!|U-���>Y�N);�Z5�
� ���T��t�����Y���a������Y����4�����g�ף���R/x��Rg�/M��M��!��x&#�W���)]�(���Tq����[E�b2�d������Oq:�-��Ao���d2}���ֆ��/��6�05���t�m����:��`rʕfy�f��
�8x)��;n�3i��SosM	������G2������7G�0�����,��
�i��T���-��6��"HO�l5M��^!ib����z��-�xS�P`
�PIƷ�x@��7���w���A�c˼ K��C`){��į<����@O=�����j�C��7�"����(�y�V��Z�v,Y��,���P��J�=�����$xP�f;n��"?�W�HP6p2h�c�����4�vm�"\+D��d�Zؼf�M�/�o.w]��;k.՝�Ӓŕq�w2����s Ӡw�%q�9D]2Qr��|�q�M1G꓂�=3�2��X8�UyP�So����0?9O���]��>]�^�$�Oi�;�ҭf\2�u�F���;��\w@��|2E���� ��(��\R���I����I�;X�԰;k�>A��Wۄ��7��,h��,\��D` 29`�1�ASY p�w�97��-B$1��^����p�ֆ*b��h�Vce[|�=�)A��di��{���J��CB��N|L���_�\`&EDYp$�)Tw��,D���~�ݛa��@��X�@� ����JLEh-l��Y'�H�q+�慊�2�n��F��H�+[�=5�B��a&��k�7��O`���*��Ѷ4��+�S�Q�&��t0����r���5����;��/�'
�����?G�.�^�H�ι&��Zĺ=z~���^�v�sH��D`DJ�v>�Y��G��8��T�Z�.h���(s4v4��S�Uhr���\b(	P*���1)�-�	��H��p9twq�IU�1�h��;`��6�daEۼ]���7^�*"_��Ls�֊��5:"�x�J�m��u�Z->,(b%X��-�A4!�e�Y�PzC��XN`���'��)P�Y��l�s&�h6��>vx��)~N\�Q�H�?�;ڝ����~����ng��g�J5&ݿjT��(b4Q,0�@��L�����jZT���o<x�D��N=Is[��h%���,'_�Rԩ(qC��,��⯻�� �7~ߺ���o��}��L2b������i�$~�Ŭy�s�N��zݒr$���5"�A�R���:����d8E��]�r@�o�ʖô {���q-j����Uq��M��%�,G3����ҳ_K��,�7v��Ӳ�w��9����*�fp�o������x��E��if��|lw8�Mܼy�:WE'��V����g]w����`���{�d�'�{�]]�jml4��HݝT�!߻�/_��%��,��ADH��3=9��v0&��\��o���r�֜Bu�o��)9�l-���]����ɢ�\k� �Gv1�K�6I�'VhOd�l��˺�$��ԑ�8O�QR����<���yOOt܆C8ԏ��a���&"Wa� �L;Où�m�xm�����:�,M���a�{'�-\+A`��0o�)XQɭ�%_���EI{3�>%�d$���%SyBw���\N�x򉪙�\���G��k��TƷV����:)��&�ౣ��:�Uv�8�"�it9�6v0|ݢX8.[��s���9"ȉXyT����כ�U7 �z��AO-	��A�`~|�Q�S�7�g6ѩv`xa Վ���}z5�/2$�t�P?2���P3�*WJ^���U���ϵ����\\��ž��t�u:��'{���d���v�XZ�"9X4��Q�<]B�é.6j"�*�T9��VW���}1I(Аt�B.�O���V����SE�l��Qy�=��{��+����������:�d��b� !�9_k�t=����Ӷ�� %�x��ｽ�����}Y������f3��8��aQ ��8�]
&� �a������H{���R���Oq��?w%�Ao o�)�(���OK���OH��/�յ`؆ͮ��e�a�(�
�,{^�m�A<�j\V�՘����`)RsǕ�z���g�QI�HP��2�=r	ɥ����iS^��Q��h�HH��ܨ6�u�����x2,'�bL��Ls�pS˟c�.Rė)Qs:�����C��'#��FM!\�)ئ�t�*ɿ���r�/B�?�i[��ڿԤ��#ײGh9���N�C�a�G0
��z�^�-=:����8Y����1�2�I�ę�3а��	��	.�+?L!ɧm�C�pPn��Ra�d�(o���\����x���ܠ�O$�cL�,������Aa����� �!�fV((�)�^;�<�;w� f�j�+	=Ь���bN�}sH���g(�,����n�v+_�i�Hh�r���R�#���d�n\|�k���6�w���ׁ�	��O�"�o��J]¿��H�ϰ�F�E/Z�o�\XqIs��E�����v�B�4��׃�}��.2I�v([�z
Ǳূ8x+R���3��U�h�����I�ٔK��'��@�z<&��GH��~�R("�����7�ʐ������D��hŮ�Df��s�L�K֎Sî�N�{�?J�s3�+a�'�a�rLŌ%x����"{����]��&Ȫ���z�����b^�3b��W<��kd�Q��bY��B ;2�A�8D>�&��v�#]����c*�q���B%��^�YB���f���+`Z0Yj��<���Ś�_�ٕ~oY����iOxL��r�[F��@��CZsH�Z�KWk	47���q�.Z6A��w���L��{�D��2����x~�~�z�����$�)���QN����S�W�f8u�HpO�͸��!��`��P������ak�~v�cv)32�<��p�)����/���Sx��~�k��+h�+MQ(�����4h�_|#/������oKKj�ǵ�E*�5 �S���heK9E��*��GD��1(��،t��}���g�h�5/�[�-I��I��͸�]Ы���Y����J9�=�Ҧ���"|���~.�@S+t��B�'�3�1��l�~�/W�M�E�R~��Ķ�&�F�% \�s'?3�V�ϨΒ��Wԝ�J�Փ���h������z|Og���ܴZ�^/ހg�e�ҊOhD������"k��;D�k}�U�[�|�9�\��\�ҸN�%�b�e�h�e�^ard����"�	oˏ�vy����)M0@/���g�hd��?��_��แ;֌ n\k`#D/}�W:W]�	5���� �{�g ==,ن+��k?�ٺ"xa�xi���:���f�=������#��6��� 9c������{X?��QP�a��C���3b�#7բQP��e��_
ENtEŊ���D��V]���s��7�Ɛ���a̦fҲ�oM],�c�oo'��(JY��.�ZV=^Q%�&~�،�Q�g�s(T��C�S������\�U��_21#�:�h|a�VpǪ�T���<�ݠV���t���s5��w7k��Z9:�C�;���+�=��K+b�ܰ�q���W����Z/��uK���D7���Q}UV�)gNO�$��ʟ*�e��\�9��X�M��'���v"�]W����%�|8����k�-h/����z�п�������=	z���"�}X'2tvY,Cm����T�Q�R1�o��K��s�-lH�������R���y_���x~��(��+�<���������sN��H-�wY@Z!��cPU�{�JT��������l����b� ����qA�����S�+�G.k��݆ƥ�Ms����<V3�C��e��M�hd0�뺫w�mg�)�C%	 -�B�JTR�wa����l�����뮭P��-�)�@B7�nO�s���t�ē�zwm�3�5=�鉣rY`��L�`�_s|���}���$3�ۗ2բ���:�?��w�!9�~�21V���J'�;�aη
��⁐u��0DB��
��
���]�*
��3~jp�.)X����%�^���S=n���@]n�U�Jq��/�YV�p��H8���@ܮ���� #@����k�M��H݄[/��~�gQ󬆏��vR�yG1�O)�ݎ!��Y񣋁,`��k2*7�n��eʸ	��hl�J ������eM[�ay'D�B.����Sd��� �`*�vDP���F�UXk�䬴>��8W�+Tl`��e[����DVYa%��)NJ>+q2�� 0����=Ǻ�1z���|{G�	ޞ¿�/�7�w�1٢~���/	=�h}n8X��)sDD�l��`�4(q���v�N�"�%��o�,�8� �
�
�T^yz<.�|@u�m�nw	V����N��!���'{��쓆�z�!����g�slF�6��a�t"�UY���^�Ș��C�*Y�H8��W�6�|	[Q��#�>�aQh�fuwrmg���t��2Dɂq��{�?�Y �	Ъ(�^VR���m|D������_zLQ\�+v0_7\!�Iʌ��Q��v�������Gt6\V_�`/霯�V��ԕ���ӯW�M�`���@�*%3I/ ����޸R�3Ȳ�0��0Or�,��_4$�|Z��fP7�BFmΰ����g����q���$���0�^@$�3B��R
��SЏ�ń��H@ѰO l�_�Q�/7��� ��7ͷ�{�z޸�:���&���ɬ,PwIP�x��w>|���K��F�O����S@웪��?��}�q��΢��7y��1�Cp���v5r�/�N�*����-�I�����{��^�H�oE`��m܎Ԕ{@�G��Ӧ�,�)�e�±����|���
���
PƼ?4�-\�~�j�c�cM>��0@��Rn٫��~ּ��ue�R�O���Ģ�r�,Mρ8_�{���ZT B��8�����O��[���\��B��h��Q� ��	�e��mo'p�1���A�?A�+,taU����}OF�2�<8���`�jR��t,�^�3�U���C���JW����`�*����Ţ�����ڕ��f�#�=H��)��|jHU��}s�@XĂ���@}cv]f���0�pi��J��Q�7��%��ȭ�`��$>?�k�����T�YI���͌���o��m+];)Z`4l����xX'+u�d��)�ʮ������U�zvaWZ1ņ@ϧzΌJ�|�z=�Pę`(����lYn!��X�Uu��T_�ּr��H%�D�o�л�V�;���w:����ל��<��9�f)�jE�one?�1����@SZ�*�F¡�\�!
,�u���X�TWY3���k��G�䒶�Y�QD
c� ��$OA>ZOu�.�	�����PU���C�J+��b�5��ݑ4����xU������ѥv�U�v�(a�o��p��Bh�K�	�T�X���'41�o.¸ᜲ�nV�ۻ�T%�R3Ƭ�:��',��L�?J���7�<9��aS��T�r�� Zy)s{b�8��>WY���`��h�4D�5h��7��7�ڕ��tX��CP�w4�s�6�q�ŭ���UѰ�¼iᛛ+<!4@c�󾷟���v��c�Ӯ%�j��JH�3՝�X�7��ʖ�T��u�4C�`�-�։/q՚��r���X��VuzW;F���bPb��@���y6)��Y
/�J#b�����D;KH+��Y��lg	į:�sXTp�'�yu�7#mS�,��1ŹB���]�2�3���&���5f?�~�eG`�	55��g�N=N��M�t��{�U��dZ|�B]���5I2(��$J�����;��c�u�i6��� 7���5�W�ٽ,ZV�ć�1?���z� "X�$i��Q�Ŷ�@����ӈj	S_��<̯t��������Y T�ڢ�@m�_i��8��0�~n����� AO��;C\4vƛ��Z[<3�#B&�[b�}�I�;Y?)z�p�z��l!�{����S�����k����A��c�o�%�������́�9r2"��jN��L���lGTB-����'�������r��iBl��W]�4�%d{hꐴ' :�2N0^��tu���V��D�H��<����D� /�A��^>o�G���$�!ݣWt'.4��E�L�K���y�_���%�|�k�Vi��ܐy,vPt���pG_h�<g�~T9Ao���j�$�ŵ(�"^�J+�Ƶ�z�����OQ�UF�~ǧ����U �@����&�aq�D��q�UǶ<�sP�qAA�@tȋ�z���TsV$�z
N���9Q��R��^V����}Mf��^��bV�-=����F=VSLO�q�;�ε�0����֋~"�Q����Jy`�!R��o^�3�$��}�����2W�pm%��h�}Z����Ѯ~�M�cJF#�!;�W��Q$�	'\IZ�1
.9:3 qń�֪̭���AN����Ɗ��x�溾Xw8$��ʹI���B�F"�H7��>��bU<1��Y��C�IiC�R�y'° ~���H��q,���m���k�]���D��j��1QIeq�zM�׍�IX�_��-�N:_�c�aз{Zc�'˟��Q�������h������4d@{Y�G����O�g1�e����CV�j��y4n�;�Tn����)����գ��1�/?��h��D�ZQ\d��uM�ե��.!�3M6�c2����eKZ��)�Z�b��	��4j89"�e�&��W�� �pH�X�jR���oD|(U.iľ��O���+���xs�m�L��F�z�o~X e�R�}��([��7]b�.ϩr���2R�O9�<di�5*�b�ʿLxn�Z*C�K���KAF�O�}�+M�CK��e�z5)�R	L��3���=���D]v�n,"�%�\b�P�CP[$��$�+�ҡ��� ���f[�8��Ω$�F8R5��L�\Y����H�o+�K\<��|`�w����+�
(�Og����Ʒ����#?�e��T�r��0�^�$���fjEC<r��yӝU˛�)r���]�օ��������zr��T��*�u%��ӛ-�Ȗﾊ���.*0D%B��J���2Ȱ	�a$��I8�����2�ړ�*O���������\�9�̭�%�UXS}��b=��5c?8��ZlPt&��v��h�=0��ѩ�P0K:��R��� '�_� W4K-+�,���2!�q2�\���>�f"�����!6�}�d�-^.y�JBY���G�>�3��NҬ�߫��w�Q^L�Lx�W&����n.�d�P��l���Up	^2�� �-�깣��H��%�_���*��l:�"�7D���1R����P319wS�ج���um�x�}H�-3�қY���vX�P__�؍H�
�n��җd�[�D�O����"_����^)E��GGo�@�����5�)�ko�cyk^`���6v-��*\n��w�g�v=�qA�*M�S@.G ��,dQ��j�<Ӯ{�˩�:]B#'���i���
�՘�>��L|�s��.�R���s1�'��E��ýc�kXC$�����5j���є�u�ۆ}1�z9�'X��Һh��蝎=����tg�e2%c�蓫�4&�.W�΀<�9�6��������l��)�|��N�����UMz�0�'���q��of#�
nG:��w��ZS}��6����5|<�;q-�I|�>_Z��z�����UO�f�:UY�~@��v
�֪��+��F����V>[)~s���~ߚA�6�yp%_�3b w>�������� ��\0��@���0z��^�� ���GSV��t�}O=��/R3�C��#�����>Mk��^�9�g)ư�<�DFT�.����se�\Or�xU@-��뢚xʆ��u}��?w?�0��Â
X�M�t_Є��bѦB�(Pϡ�^�$����º� 
�:����˕7cװ�|o��Ӷ̴<-#+�D�C�ߴ7�*���� ���,ɐ��ۼ�u ��4)QtjúN�u/`�o�)���o��]�&R�	��M����LF��K7�o���%aޞS�;�y�\��L�������&��ۇ���ȍ�i\��N=>�Z�Y\�y�Y��O"b�����4JW�w�0�:+��6cl�2��W6+�3�I3���D������ Ud���t�b��*ܒ�
n��M,_]����Z�&�;� ��i wj��}�+���A�g��׵+:Dg{m��h�.:��C�+Y4v�3X>�"��Կb��8ϝ���e���U�<�c阮�c�"7�����>b������*4a��9�4�0���ڨ	��Pi�|%ֿ76E�����L+EĚ	�����\0\��F�"�P�5�em������e_�{w׳��˶g��G,�U��7Hh7��Xp%�R-=�/��a;-Co��q��F)�eA�H�ն��P)�@��l�l����D�((X���F= t'�LH9.@%B�y���ggʔ"v��M0�*׮�C��l䏝�Z>a[
�O�_�d{�Zh]Ϟ�'`Y��+��_���ot��+�[�=��!�R��&V�&�Z	�G��@�3�;k�Hf����i�rD)��E'��@o�V�2��������-W
�^�[��b��&��S渮B���T\ryPA���ͯ�u�FSs[vk|�/����/^ϱ�N��A��tX5��|w9��E9(��qk���~ �m?тA�6v���~$�1�H�
�Pjп�1&�U�\/W�toڴ�V�t�`/
lu��$�g�k���ī>�/�rAǟiq���n�	�� A���8�K�ݾl�=�Cѭ�m#8!�{�j����M@���LnNQ>��F�JN8W�U\DY�6�:���;���k��^M ������~�F�S�<(a�Nh���s$�i�+�\�s��u�q��
�U�(�"�b�j�&t�(w,�o��4R�r8~И��7���ͨ;R�1)��f�H��"�ns7�����c�)h��f�AQ�'�������J�����Y����o��I�蜻�/�,���mʽO�[���d���ṻ/B���Y�u���&ӆTEµ�?xw���A���[����0u�C9�^�>&��!{���hxzNjl��l=+�s5{�e_jJ8��r�3��^y����@����?�ˣ�{�Ӡ��9�vK� ��ک熢w�*�0�r��	��U`���3����bW�Y��5. ���n#%R��,��_~����Ձ��?U�9�j����6�.KI#g+
��5��;u�х�h�ڎH�Q2��r!>��p~eH��D�?���IY�.aڡH-���D��k��3�p�����a�XI~E���]޶x���fE�fyc��&(�,��:Z=�I�% ��g�}�P�^�`�'�y��p&DJ�����g�.1�~S��ϊ��w�Zb|،)ά5���C�2��l����m�i���eeiCԞt�T�&�v�\^�H�z�g,��Ă փ�����hW��-�'�sB�v9�H��H�R�n��� '{D<BF��[�ؾ \8�˕N��j���93cF?3�����ޞ��s���֔�v���s�����ՂT5(�w����!��y�!�*��XcHF4&��]7@S��o���mn�|[=�fN\7鈥ח�;S�ʦ��Z�+:����9�_��K���V���l+�X�l:�hn������l5<x'��^��ÕƩ'�a��mX�&x>+}Gl������4stJ�ʵ6����7$�rlY�"��3���92ښ=4���^O��!�E���-����7���r�o?lN�U��o��H/���jիN�7W�8��S��"�F�����[�-T�]�6j6��vCI�N1(��i
d��|�������;������6�X�볮W�ጂ�?�^H����lO�m
��N��lq��6q���-U�1�����V�������]�x����^���F
�ժ�L�/��)1{���8+����ϸ�s,Y�kߜ�Ob���� v�S�&����y1#[o�q�m&�6+.�tg3cjš�X�=�O#�0m�;:M��Y$de6ޘ^�����؄���)r�0�"�_��<:�vN����g ��;�V4S�`��&S�B�P[C��E�,M���rKmf3ӑ�@�W^՟��i_�(t-���D#��K ������V�!{���7�z�։�j,/�9��i����Er�v�yy`o^3>���簹���/'���X��\kH�	��A��t�������KVu� r���n�F��(���lЗ����0�3W��ڔ�v�:�.�~�tD�1&h }M6��d�w;��J��E��!w����R���!�8 ���,�[1��/hhe�0��hK��>��p�e��I���+��(��'�$�W���������DN��㏔%���}�3��@�r��'���
.�Ͳ�ξ8��`Z�mt�9m:hV�VuE�M͹���|���j�3h��h_���n�}h\�P��|�|0d>_���f�c;��g�t��l����ﵿR�e��b�Č��¶�U���5�5c�O'b�U�`���ª(��E*c��r��W6��L@^KQ��oSC�$��������H�i���;�E�����H3�!+z�:xPc�U]/Pmk�2@����e(�|���8�G���Jr��|�u�%��%�͢���Oe�\=����
����4���GĲ�A?
�����40@�(��G U�ƺ[�ߑ)��VÛZ^N
ʕd�'Ў�`0��IF��)�7���ݠu��'�}�ͥK`�����\�S^b��dl=��[n���x;!�[�7����R����o��O���Π�����4�C���u��`��♠��⪡�� B�Ly=�L;��K�6O
��6���,:�]��0�����������v�ﺡ�G�/;�o]b�%n��Jx�[��#E���r�| ��|�!����8��ւ-�6�V4��ݤ`�'�G,p~�b�L�N��B�^���V�`���،�J[1Ş
�̅BR̽m<�[��6H��om)t%���h�c`_�TUҋD�qq8�7$o[+������d�L��^�j/��H
��2Gb��H~��Q=s����f�R�u��	n�ڭ��`R�g�^��o��[s97%��i�ru^�,j=��Y!S}h&��,I���G��4� @��EI�����@	d�0xY�_����68\� ���./P���-S�-Li(1�s�ǌIr�ʴ�ʖ��zos҄l�@�뺞X�X��j��`�B6Bh7�� �^:URA_X}�r���L�u�#��>=!��ӆ�%9�S�cVo��i��<�%�#��'n�&R��Ĺ��W��v+'���v��inv�ڦx�ч��^q�kj}�u����s�[`B���GN�M{�J�=���� �Te,��6������s^s��N�T�ʩ�_���K���y���y.������!ǰ��}ⶅ�҈-���y�H_R�3�$=.����Z�����i�Q�y�>*u�Q/��V�͘g1��c�a%ؑuqLH�%�,❘_���N�A�j��2�Ł*[4��;8%��J���l�ν)���0��f��,�1���S��{��Be<��-�]��Gt�k81�:@��XK��Yi�H(w��Gq	I��0�ae��ᬽ�1�!M&$^�s$�	<�o������y^�5BS[u(!tICc�Z24��e{��� ��8�*�O@䞲���#��/��-�䛉oS����q�����bV��l:6��e���g�X��]�P'������ݑq@�S9j�ǹmdA�8��Mo�E�R���c�y4|fuoN˂�!_���0����(�I���f3�0���y8���ç�����sN\��Qp�v����Ӈf0.L�z�̬������� 3�_t^6�v�\j� ��9�̃6ќ��Q� �x|%~'���H��<:Tَ���#A+��'೯�][���v��e�b�=T�~��������#b*�t�R�S�>#�1�'c��5.��7�C.��l���K��c���3He=�!�����q�D�Xui�P�G�^y�U=z�1w�z�'dqʹ"V��IY����tWX��Ġ���;�rBU.T�V�ǣ�\�c�(VL���.3/�����)Y������j���ԛ��j��fUk�r�
�_�~D�׽׎='���2(�ȷ���-�`><�%���q[fpqh{?Tu� 	lkTe�c_i�ć���i��3+3s����^�4��X3X'�6M6��y�~6�/��+l�-�t���Mjy�����w��V�b|�=���ˑ�Sp��^�����VW���t��vJD�]�"*��6�����R�ź�(b��_d�e��cG���kv]�ƦU������rt~�ɇN�QZ��B�3��<l�VLV�ӊxST�e�%����>�v�0� �@#�c��8E�]9��;��'b�N*���ia�٩9�#�GuC
H�כ�����w���Pf�ۋ�r�,����v(��"�z��_�P�����<��y�P�[R5ڜGU"�D�K�ں|��/W�����@Y�6�����1(�3T���y���{��2=��}�wh��$�=)iG]ћ<57d��r,���X&����Qg��h�4�0�C/\�-�zV��eL��D v%Be�����m����������{��Z�n����_����!\���0R��?�X1L܈��	���������5�f���-�.cفN���3�h|J�"~Z�>yK��m8�0N��v��v0��^����p�#���V!KH3��Աx*(�FukfN2�U 1���8LP�P4T�-��ɢ�-,��A|�eοE�����s�B1ơH��ȣ��O�Yd�i�/L���A�+� ���[��\"�-*2͎�>]�'`��A� 1H8�ݰ�tP� ��c��&F7V��>�<��{�����y�0^U�V�U0�y�\Z]�3-�ѿ�g�,��Z��
L��y��*�VCv�vV�2��~^�e�"�A������	���_�T��b�y���f�m�+���!Y����dJգT/pڃ��Q���)ċ&�~ @��nm r	�ܾ�?�=�!y��Y����}ϗ�s�ڳ��9�&���.6��ޑ�$I+��>��<E���PO�C	�?լ��[+�I��3����Kt���j��~0���
��ǥրb�.��X 3���՞�-�O9�����H�������S�Xt��?S3y��ֽuؒ�t�K�;�v9����������f2�B���0�>ew�K�3�}��:TUv%��Y�$g�bvֻ�����A2�ٻ�@̪S7/�E
��-��ԷgM�}�ZS���g�.��H毅�j�)1�5���M�hk���݌�!N%������?�Z\p�����B��tz\��ZE�2��o�-�������"g�a�ԙ��O1�Luj9*��]�-���H��(SbD<�kH���O�����0�M���㟣�L�Fs�o�i"���s��ĠGt~�X�������IZ�Ua�5�ո6�K��qhQ����'P���u�28n�4�g�|��j��hS�O8�FA�O�#��N���Tɭژ[U7��'<�윞���q�p6�LI��+c�>InL����W�S���(_�d3��u�)+݆��+=C��/\!q4�{��l�%KΡM7�2ww���U���E:����m�.Qx3�b>�K��^�4�75�x��$�w����b�l�ŏ���~PG|�M�Pk��֍�ǚd(�?�Y��/%�����L�ڼ�
F`@�z��򡎓)�����7k?ٻ'�Dف���?���2�f�1�Y|[T�&w��H�rz
��M���C�e?��f[��I�U����u
��U�#]娬�r���T�|���o��h>NI�+��������+n��T�󈝪����m��Պ�ˢ�>�Wb�����F�®"aT�_5�@����ܮ�tO���^���<�[���������c�}X�������[f���Zd�$�`j2Y�F.4���`�L{���!o�~5)?ik��t��@���9+�Fh�o˻w�#�iY�U�q�TD�^'d:�`Rg�<��(C�tO��e���2��{mVᒨP�d��c(ńT������&ã���(����dBB�<Y�-�E��~�*��}x�\JC�G����*�.OT���<6-�(�9p��9b2�Vݖ��ePl�j!:8n�̬s�9e�gH�,]�ӫ-k�@ ��fV�:1���P�<1\�����؟s��~�>M�O�"$$D�����\v�
���%S:ҋr��W�b�����2{��h�Q1�n&�7� 3&a����H�
_���0}�FxC����?�'��#`�ɉ�a^��D��|���x������j�y���C#��W���!�}#?$��8;1/��+.�(��L�*���c�k�ӭv��iga=}����p<���'�M;;���r�0q����;���0�d�����*�N��"�;F|:<ۘ@��5+��^�8Rś��kAn����1��7T,oY����Bsu2�y+>G�=)T�\[���Np�}8����A��_w�Ƞ�s��Uo	=uyK�&5��F�3�4?B.i/޸�
c53�-˪���姍���� �'���Ǳ�S���~�̀#�g��yE��>p_ڤ�|Uy����� 4��mV,Y�M	���7=m��YE�&�>@g�(����	g�~�VUB������=�V�������x��}�X�%��,��+f�	(�D}tٿ_�.7:Set�Ʃ�_�]�����/��-�}���w(//�jY�������hIKqsv`����8eX,3�W�=��Ԩ��*S5S�l|L�P��U6���}��=Pxp��?�i���kܿ�+OBo\W�;�h����|c��YxNl��۔���1��$�7�[g����a��C�~���4��{Rg���}e��o,:Ƨ(��đȩ�LB.ѴY��OhO�bU��h�wn�x���Q,�W@�K��;4:5}��>����a��M��x�YL�uG�4�3��!9E���)��ۼFڷ�$�'�\�'��+��N2�"4T�-��`G���h$�s"ˁLyy�{Y3d�W`U�#�b�@y,����>����Z�����l��>b,�7�h���<q�]�F=%J��X��C_2Bz�ĐQ �0�����wKl���/����"%'��$��(;8Qܐ��1!��n�� ���@JDUJ��j�-(�V�-���W�)o:�z�sj�*�F��V�a ���*BYL�Rh�Ea�>ó�^�kl�t��+걱Shq�̋G%[a��ˡ�!)�r��p<'����aW�0&����V�I+�G}=K���oh�S�(w�Sف�j)�������0���p��q���0x��%'�r��|if&��z�-�SY�����"�Tc�t9�Ƭ)@�T)�&zbq��Ng�Ƭ��m�79�863��`��:�a��1QX"�Ü�B51��ּ ����Z��J)y�^���9����v4��j�����h13+�tr��ByRS�:ê�f\A�6�Z6�z0̨��p�wJ��&�$8�,=K�"x��+޿�cT,�j2-��9-�Uk�6 �z�u\V=����Jg�������)��򤻭��=�����ߌ�%~D���/CͲy�\����e7p�+R��F� 3�[��
��f��L��LE�p�+Q	Xg=��?�!���$�y�}����<��[1�k@�pp�1�/�ފ�ӭn(�Ȭ�ǒ�'���JN�<����n���cҽ�9�?��9l}����Y�l,�ܾ���틜)>$��E_-�M�$%��T3�ה�g"��3��y�+u�����'�J7�=��9|�N�#�H%Wfܯ&j`��7	:��y0@��b'�\��Bsj4<Y�d����c���8�o, ��� �XϽj��ٛ��53�Cm7M�t����N$R��A����c� ��J�%�V���(/�!c�'�9�w�b��;���>�t�=��64��u�8ҥT~�^*��PC^��B
q�S�5M��y6������ъV]��a#����[2�B� ��}�����Z��47��q�4�N�҂S�<.��g��h?Qc�������Z�"�gz-{�DU��ŞI��!z%e*�\�����c�Bҍ�Ѣ�Q��t��ͤ�"zy8���`&��1I�E�W��C,��nm�������Q�E����?�L����S�H���R���W,хsQ��އ�jPTA�mR6%�go�],��"$q�X��Wk�/�aYP�|�bX!OX�|K3�1���՛x8W��q���N�G����$r&�l����9�d��q��V�b��_����O�(��f��P�D�T��t�Gܷ���h3�[V=�T�a�Rͳ&���nj5k�&M&���Q�.��Gc��e��:v���ڹ�Y�<5�qse���G�=1�C�'�b0� z�q���/r��{���w�s�G�\
/HC����y��U`D���
=���i֋�����1����-��Y/	i���A�$����}Uai-*���ѝ��>�6�}l�I�(?!�D�P�h��2p{�dg;�E� �N}�&���窧���x��= ��dOJ��R��Dͮ���tz���z�~�[mFO�v��ZfH�S0)sƅ���4ɥ�s�Ibz44Qk���Zp*P
tj(��d�U���ĕNDD�n�K-|�x��D�T�:/Z���`B*�
�&�	
�J� !��9��rT=��[�`D�9�����c��t{ԫ��,��� y���rD:~`y]4��7��oW��5 ��@iDd��7�ެ�r�D+��IժY�f>���]��u(�X�`)0�Ɨ)y�^q7<��Z� -��(w[�:�9�r\N+�(k� )�{%y�����IY��N@9���Gy�����6�OR��,�E�{YĂY:H ��`�8Q;Ծ���1Z�|��^����RL�(tR4o���'>����� �Pnp��p��\�ϐ�˧'�	��0w�]��MI-�k���}{3������{Y�]&�]�e�kC��+��u�9c~CE���#¶�QH�X��#�
ߜ�˟i�[��dQVo��m�]#�Zr��æ�,�{ؑ���J!y�����Ѱ�bR��}�T@���k���<���w��0�eY�t
��y�{��b��ge쑇� ��L�y�d9>�D��d�I����"%G��	�lZ�	�z4-,o��gq��1�ܤ&���4x��/��j��q��K]�6#��
��w�,|�U��\���2[΀f�B�1�DU��6@���߆v'��Z��d�X�v��L(�Uk c(�q2dNK}�4��N��#�i��g��,2��B��h��VYa̝ޱ����9�#�?@/C��=Q0�Q_`�4�b����R�`-�S����������.QZ�&�y��</�k���2�"=î�罛�:@G���>H�M�ؒ�U<3��0�g����|�F���'����ĭ�W��&j���\��`g|"_��r(�dT�]�_w�*	br�m����T�c%,�I�}��[�7����SE�Ao�I���	����_�?��n�Ӈ�����n&�C�ɞ!JM�����(�Y.�홞����F��u����\f�}��K%ogŶe�*��/y�'��Wjs�`�k�DW4ɰK�;����7;�$ޚ�S��%��	+���B_�LbP�K���ǐ;�Al��eў¦>��2��kjgȢS�%;��.�|z��,����ܻV؛��Lg@)�TótGg��^
M�}b	�ˍ���P9���Q�5�u��ե��o���#�d[�)%=7H}�P�!�д�C�t��9 G`:Ԋ�}�������&��n�� ��b��w�����`�i�W+L���k���4M&�n���A#�5�#�Cj�G�9���vzC]O��5��z�S=�R�L�ɇ��s� A�%DmY�
k5�½yPBm�O{�?�g'7z�b����	�j2�g�_���
�����ٝ�8ͼ"�q�_��5$)ұ��T �}�`��A��"��T��(b3f^��_�d���:/7�1�˯Z(��e�2���XM5PV��b��s���o]r�X�sxi@���_��tʉ��y��2 � ���qw�j��P�i=��W1ė�-��(��W�DG�0zE�V�aSP��{_ٴ<��A)&�C�f+_N��G��=#���MR��=��
��"\�@=<d��d�C��2z�)V�e�xLa��<�~fƢ�����'�r�>5Y���s]��6�g����Cu
&D��u-
8'��uW��Sq���=�-Xoj��҄�y�ݾ�UI�s�zPY�)�R�C�	Y� �ٹq#��Lޔ������QhW� ��.�7�εw�{�y��6�@HB6�lj�b��%����8."������i6>��lcvk��<D
�7�=�?,�LWx���� �R�l�Otw6h'�M�g�{���Y�(��ZJ�#��6�S�+�������3�Fؗ;�ᾚ둍�[�0�<ᧆ������V� �����ݿ)(~�p�j�� �X����2�Y���=L(FR��x�H�kX�y�A�9��ע�N����ܣI�_�2�����9�5�~|���_n����ze���2gLj�4l+	�����t�Jm�^3�0*���bh8T%���������fXv�v<D(J��M'���n�+J���^�}�_b�з�$P�����a���=^&��37趫�7���)�	���3��������.K]���r��&��MG Q��0�ʤ���d���Px[C���}vw�/�d9��c��4��
_v촩��|¶�j�W�=�W���H ̘vx�旅v�i��7�s^�|��q��^_�&�iC�M����G�Wo@�]��00��BL�ǭR�HX^)�����}�+mp�]��1Et0��J�2�2j��ϵ�&w�;e���'��Bc�-܁Y/��m�"Q�v�lj����t���3����$�C���5p�3_�ۖ��E\(rf6��!��3�$�h���(��!�D$�]�[�730q ��_��f��Ql')�� }�St��J��t|�B&�}r0��~zk蕢��u��G��K���D�D��-)��:���' K�5��u؅���=����LX���ô��i)���r]�� �C�����J��3ʾ�W�* ��� T!XL�{xc�{�OY���X���C~�ׂ��0�װO�i��d9��#b�����jؚԏ�f�,���)�ӓSa]�w� �B����-'���F��N*�/����?Y/ �� C;k�O��s0�t;2���Rw��,+�;J~bקp���I��DӐ��!����cvX�8��I]Ǫ����8�E]v�?:�0"�ܚ@���0§�;!�\�V&�2�}ü�ނ������U���
�1�f8(a���S�;��s�ؽ 8�W_e�c;z�r�o��_ �����Ê��������*E� �O��ښEI��I���K��\�>�@n*�*` ښ��cTs�r�kJ\d[����8�v'�=�l��˾疹m�tsq�}�9���gǽM/�w%	W����W�����2�;�X�m�Y�R���9�A�so5�g_0��g�$-����f���O'8܂�5�`ј�xEo�RU���ƸuvX�;ǙlX�/m	� H;�pXƕ���-b_� ����G��x��<
T7��		—pVܦE<��LqʖK��@�e���b��"��T2Y�W���0�+�4h���^K;���W�4[�В��xrR� v+���eyWFt�|;��ΘE�#z��-6'�p�	��D"�n��9t�#�n"�@*iw8���4��S�R<�l4v6V_�bY�p�"��Ux� k�?:���"�.�j�XbQuQ���~�G��m��=ڠ:R�|NQ���<�n��NZ�
�e���R=���@g)kY�T
�w)kT��S�`~��䊶�d����Ҙ����5\��|='h�5��lЋDy8�]̔��o��d�2KDJe��T�	�';��*�����a�<W�i�.p���w\��(�AĘy\� �R�¸A:cl
#��wC�͂[e�3'�xH`w���tYU?�(�WPIJ����Lk��^������ܬ	�7�,�cJy�L�4
f����x@ �fF�y�U*�_R�MBí%�P�a��D<�����c`�:J�>5p-g DNހ[��z�;g"�&�rp���7JS/O�2��:�G�{Qt��Pd��	n�����c�6?�c$�Fq|"�LJ|���@���SP�u��ښ�Xb��"|�zO���}��O1G�&�:�A�	�a��8-�CMt�6���{r����$��8�X3�Z��2e��,z�MK��l�Y~�\��ģ��f=f/�G��G¹gX ���H"�R���w�Ċ��Kt�dV���� (6��۔���vfۍ�A�E�={���0�64���ݞq��� ���8���e�<��F�d���S�I�
�r˰�͘�8�ӂȿJ���m�ɡ'�T�Qn�^~��Ċ$+p�'�}�7�:*B��ee�� 5�ߦ�3kh��s�����-��.��#��n���O��_�RQ�ɩ�cL�|s�U����7�a��L�ү�
Fm��m0U"���O��0��%��~���>��F{ʊ:�����1�1����<�֏�J따�U�����N'�6���/����,=�l���/�!��'���%A��ʭ��T�1[�漗�F'�K��5~��-���2O��Z�,�@�W_y�l��.1x�o���Y�K��BbF�;"oI/��+�7��'��m������x���������Jn�O���Q�/i։o;����Y�o��f޵/��&�'�}|h����s�>E��;�H(�&�}/�U8�u}j�S64s�� T�fXј̋�}�1��sH���\4a�Qv�M�K#l�K������QwC)�_dI*�x����PbJOYk�q�+2���/*�=����� O�Cp��6�]�p�YKά��l��#�h�g,O�0�ux/��)��$��Г����t~��:�!���PY�K7+�:3;ʶ4*X�(��}�[���RFB�6�(��\T	s�x���
+��ip����*�0|�~�Ʒ^����?�����i[q�R��Gx�tMH��+�0�1Oo;����.�5��t>e�x--P���WK���zP�#��� \�Z�|T�(d�"����x�dי܅�H
�/���K�A�q�Øf���(�xǺ�����w��Њ�w�`0ӱ�����+ı��Y&L5��'i��9�*|-�J�?z�F�Fr�>�@�� ��:^o��>7܍�e�qU�m&J��-g/�} �4����y���<��4�+4�)g+�C6��qF�쒧ߵeRL$�ϦC�$ѳI*��JS�Xݷb��oT�*�y�5"�$"�S!� jK�k�aڜ�,� �t�L�Z��_{��ԗ��!dU���l�qctiȼ_c��3��9A;.�O?W�O�{c� ��"G#�}�_���A
��H���i����:/��=��� �M#Y GTO�v���ht��;� q'���#>W�JU$J�m�-�IM\|�\� �96�y�-*B>'Z!S�k2]�9���<��~�>��8�/�5��&O}$:�N�!B0��U�^lm=�c�k)�VL�l��^�U{D�wWqڝ	啥u;Z�&!,=-]�/�6Ei7����y	�������%$���j	¸��
��H��eczZ�������7��"{�Jx�M�ZX[r".�RYp?K�/7�?���##f�Np�ͣ��.��¡�i��~"Vo��s�g�R�-�54�H(�aK[A���{�ߧ�ELg�80�q�dWl��h�N�H� �_Q�Җ�sB�� ���;}���#Cb:�ח{��F���1��N*�[�#?�9�����Xܒ�fd�bW���٨�cp'�B �_΅�nd,9��*&�3,�|BϽ�J���ʢL�zDl���Y�d�ĸPj�qpR⨚��~��GMݨb�Ass� '-G���4:V2r�d�+�=��5(�$c^������^��{����9t����q)v�j�����q	=N�$YRÊ�Vi�s�]c��_���Ee�:l�T�٤�(�b=��j���&�ձp���S� #a��g�QJi��'\<�]e��P���=�a�~t��4��LM+FܙS0G~[��G�*iȐ'�ҹ�t��Y��;�R�/�MH"�!ѩ����nJb!�'���B,���de��h��T�W�7���||���(A�b�7Afx�´G�������'Q�8 >U��Nj����iK��	�r��3��2ɔ�)�1��yl�U��o�0|���	)�����#�$�c}��-YFi�={W�p
;��8��ծC<57�{5�$��ٽ�)��ʴƛ?��u^����y�C g�G��/ֲs9�S�~_���Ϫ1��!�c��>�`��G)��;��=�b�ަ��BV�e�U0����m�y��n���4�9m�"򅾘nfc�	Dٷ�e<grBl����,j�X�K�{p?���v7 cG�R-д\
�� u�U9;L&ne^�;ɽ<�Yɗ��1��fL�͉	Ȫ!�\�SX�#�ؕ5~���ʄNܥ��͉=�\X~T���J� n��Жksv�E^�pW��=B/�xu?n�k�.3��l|�
�H�󴡌��Et\æ�QG?v����Zoe���p� b�̋�k�����ǇMe�;[~�-@h��#m;�e� ��b�ͳ�GEF��%֜��X�}T�������i#`�� ��v��,�ȳ��I��+��U��OاM�|����<%_G���z��8f��^{m�M��6�OM�K�]B8�KI��	<}w��#H'hN�j��]QE�p���4�Y�⾵�ʩ���N�� ��T��c��5��-�Y��c��I���������6�Z�&�Q�9��	^8�?�'nˮ?!h�x�3���y��1�o#|�uJ�҃�^3$�pGVcT�Mk���X{��3a����}�z��7Z�����9�]n{��S@�B��!�0*(�
�j�kx�j�E�)X�O��O�wj?r�:��c��״�e(��r�����p���4��󗰢� :Z�������^��p�ň�O�,5�л��7Aj�k��/�׵���&U��w�����_=���T���~��|��T~Lq�A�H�W��,∷3��#�e�e��]����c�b����Q�(ܒ:�V>��3�;j���LM.'s�@�����N�](gZO�KXI�y��*<��+��r �ͭ��1��D�n�l-�o�$�rh<c�(�J�gI���b�|�G�I����"��^�>���Q�!���Z�*z�����[� !��J;Uu*]�[��)Z�gW������|�v���呾�D�47�o�wT8`��F3j�P�a��x?��bĉjp��<�
R)�&�������M��l�o����������,G��qĥ՘G���X7���&ߋ��={�s�"[y�^����,���%6��74�_�����H��gS �T��ԁ�m�h�FW|~���ר�Sb9��H.�A�+��<��T��;�$!�\=b�(b8!��h�6 [Kժ\6r�Oo��K>1O4b#��p���fj��
�'.�X�/,T��J����10��� oM�f���� ��dѾ)�j��n��� ���3�#�2{�#�	$� ������j�� �M$u�<s���f~kߟ�aߪףl����+R��a�5E?3����ȫd��l�=i��:����*��ܶ����� �N�C��56��d��%���
�rW�rW�kh\+ 4�j~�ƪz�ˣ�v��x�R9�4����0��P�0x3Hy�j�t�2hN�a_Y�>�ۇVPՅ���3d4��Ef4�dt���P${�=�����4��}!�� ��T�^C��{\��R��.�z��a��d��^��"K���G���`O���*��V�n�M4�$M��Rl�$�M�K^�=�Ւ�|�=q�>���N���E%�0 Eq�T�c��B�P�ddp��Qi#���y�1�Sӫ���%7@��\��$8W �*̬4c��,�h���"#4�T`���.6i=��L��E.	����\�N%�}�]cL��U�V��<�; ���fg�-�����jI]F6�?qq��U{�����N�FC�/�M7b�uY$�1b�"K�g�j�pHtc�U����s�RdbhP�|�x%'!B�m��&�H�@I�:������f�c�X��C&�?����rS��\��/'�/��@21���ǩ�32���LC��0ӹ2�{*�Č$��g�r�S8�/���6.�R4����1�X�=
������n�1����m����LE�c�R���Z'?ɟ�$q&�\��:B�-з���E���C��ź�?w���y�dZY.�ܨ!#Q2���q77ky�4���@��к��D�U�=t�T�z�<�V��` >�ҭ�E�"z,u�͌
��3��O� ��N�h~W�͠�zt�HK�D�V/' 	"/��re�yX����D��3~,�6W�} '�ss�X}Lc�@��(��b�9�~0�l�E�8��@�O�F�<�]l9��)U�P���IPX�GS��y�CJ�l%�����K���R]}�lwL1d&���JM�8v�C/�~2SV`�C�ZM취�����#�� ?eC�PBA�9hu��S�����d{���Xӑ����B��3[W�o��N�O�C��bq@�
O�d�z�t�m2r�@�u�"v[��[$�$�@Y��(~b�G��o��� �6B��e���-<ʐ?���|�zDn?����>�-�G1�aˆ7�f'��qzr�FRԡs�������A���s���mP� ���Q=Dq�4[L!��I���9�AF�;�[���@|c.�;?<5Bu��lw!���������n�Q��Rғ#M��)䭝��.��5���z8�H� ��	��M2;�
TGM�����c'�85`���2�3��'�Ն#R��f���E�9o̞��#(K��8}�x�a+�����jo���g�;ђC��O�"����X�06Q7��#I�:��3��t�td�eA��N�=�"����
P��1f�5�r�
��ݯ�$��%����M�$`����cj�i���W�>
\�=���b���Ax�4�<���F�7��i�2P�� b��Ti����M7wo;@���s�͔O
��K/��BCuta+�;���U,�lk�4X_�,�`X;�,{����;{�(3�y/�W��m��!9��ǡ�z�0�(�(S/�I;�P(� �0���0�9���S^�uڪ�K��N��vЃh?��n��O��3�,",��$(k�K3K�]_!�R�]S�����u����ƴ�Q�2�GU��t^Y9e�g�r	q �C�!����qL�.��*��T���(��Pޤ�e�DE�9�;�|���Ȼ'S|���%ѝ�7%Xϴ �0�1�c���0ѱ�^�F t�i!|���?��@�%����b��`7� �Et|�1��p3&�����(Wf�ϕf�D��zEE͎A��x��w^��;��H��n����Ѝ/z�{Y�dMia�	����J��M2"������8�����{U�XPo���I
B[���.�Ġ�R����Vj'�#����E�������Mؓo�ݜ�U_��s��^f�.��8��nmq7~�nt<\�F�8Z8|���o55Y\���$�u�MyIό���Bݱ�j���#u�ALO�ڞíH�ԣ�{���.�P^[�:�a�3��S ҟ��Δ1I4-��o�h��c�	�!��,ý�� O|�k�	�C j�/W�X�*"�U@�K�)"2�H
�sxq%��J��l�������^���q �	��zX���-ٰ_�q*;�Ek��Re�u>qr&��J��P�	6�� Β��N۠gBj��~:�H��SR���ϥ��Y"�a�>�� �2�0�:ׯ�� ��_%�56�w�kPDJ^��[C7�}2���6���B q�`�?�C�Zg��LJ$�7�[9�T+�f��������-J=��=��c����b��<)ox2�g���o߳����*���]��c|��D1�=i�1\z��p-Y�<��]�)�NI�7�:!�*��>:/)�] X�|��Lb�OhP���W|�ؓ�F�y�9L�*�^��i�fk�k�ȸ�6�L���+N9��H�aT�o�Pr ȋ������vPG��~�2�%�	�nsv %$��}�/"�B/���W�gu��:ѽ�ڿ�*v��$׊�$5,�8�r3��X ^�˺��`uޗ{��k���_�hJ��.��R-��eG�{�!��UH@I��=n��X(����}�B̚���E�mC{vTN�o��
(�ϯ#E;��/S:� H;������4$D�߼ﲊR����ٳ����	g��s<  ����oc�𩈋pҥ"cJ}mR+mͮVC�����~qH��9	��ܥ�s���!*�&���7E��k������,����A��S���jb�c���h�>I -�*E�twŏY��(^Anv�X�.�~@7�W~��M�������~�>�|�"=�3G�G9z��$u���9W�@��SJ���=M���U���f����Y����U�[�F\���g���c�<3=@���3Q}�J�V��;[g�����8�Mo�{��0���4��11��c�z�!(�������Z�R��$ol6�-�-� <2s���1­�R����@�{�z�i��\�vs�=|�su�l/~����U_U~ܖd�J8j;>�r��Ȕ��]���_X��w�bvJ��c�;I�@��z	��S���/�9�4i��>�j�y�!���z�#����(E�?����zusr��i'�)�&�(oI ����d�-�W�d�o���`��|��N��O������Ӕ�Т�R������=[-�uH�m�+U����-T��B���נ
�R|zD���?k?�M�#J��$}P�Q[���o�6��{D@\����/��V��_V/�2�����@J��E��t�}#C�]w��1���GI��bT�+�B(T~���H�2Q2l*�s��������o`2�\�kE�t\;>�_[�#j��3��P���M�������8�i���i5�`g )[��_���*ݚ>�?>f>��q�e��y�s�2Lԡ]A�<�9!T϶`�B��SQiS<X��r4�q�dج�����Yx:��B���ߚH�Z��Z�Q� f����鑎~�g��Naq�z����p�u��:I��q�0��E]Ӎ ���;�,0�ӝÁܝ��z5-�����N��Q�Vs���3g-�y�h%ǝ��O
b��M�(��sR%�)��5P�<-�8���3�_9Ϭ�D@*��y�Kp�x��j�^��H�"��h��ޘvu�m��Z�����5�<d�VA��!;��>�?CPԉ�/ GM� ҿ��B�p����?Ѱ�aY���|OΖ:l�C�|�����O|Ҟ�)��C�Ѷ�߸	v*,��4s��i!� ��u���"_�H[�x���s]�+5࠾_����:��P"���5vԘ 	��-�{|�4����Dɧ'�y��+�Zp�Q:��<�m!I��.%�8�L/f5|&���E�*�� 8.G�J��,�4ge/u��o�����������}�O�{"Ch�'��H����{և�M�}o�>oC��Qóp�X����f(,z���p3�}�T�z+T1f!���_o������*.]��ӭ��� Z���Ibu�,=ӣ"W*�[y+�FZ��0�抓d�"�'�!
�]��o�K������@<*T�]x�];j���/aA��l:�wq�ֈ}��>+�d3�&q�gtF �2@~��eX"�w�ѓ�C�@�~�D!X��8�t �ne���D�?�P�Z���*���r�۷>�1�]N��5���*vc�1�U���3��`oj�p�J�s��J��j��K�u
.�]<��oYN��S���i��uǊ���A��b� tFY�7ԭh�BF��J "�4_�nxS� #b�^ z{Ҷ_��Zs2 �!B�%�{�Y��(mq\�'^.�/�Ԭ>n�F_�>1#����nXj�<f�gZ�[輅lta����P���|�C�n%�aME�U-�MoO�&v����~\m���"�h?Rrt��Г����Rmc<@UT���m�y!II�-��'w�`:��p4ҟ�%�ۯ�A�-�>]�n�j���w�g�J`�-��<r�M+�κ+f��ă�9܅u�n����9@�~��D���Nbg�;��ZV�6���������9���E��֯h�O�f]w$��Vdy���j��g��[���h�iΘ1YŤ�׷%g��]��`���sĿ�\K�gZ�V�VsS[�r���#��t���`*��B�
p�SԴ��al��*�NW_�r�Pܞ $�`��;1x�s{a�u�B����y��ڌ��h�<"�~ف���=�k �Hfɮ��6��CE��s�4\��Sm��ӓ|˫CY��H��oJ�l�c0mО��/Oz��h��f<F��am�����)}�A��������� ��E%E�aKV������ϝ���	[����߶�mS�����sE�$�v74�#�AH����	!���+��##�	wAx�tɁZ�'����nh���5��d��zlݜ���n3H�o��1�\�v�N�q���t�8���X�4��OҶ�bC`���O)�Ĵ&3�E��<�M�|����D�1�'������Z�F;���:Oq\��>/`�L��>���^�������5nAXM���k�����;�'�����j�EU
\ )֮�Z���uB�_Ϊ��"�x�t���x��B�Ld���]p�a��v�3G��#�\���1��^�v}a�+�;�3��]5�>�
��>�לN�t��X>��K��zFl�����pڿh�itrf��}�L��sX�J��Y�t6A�疺���k|e�^륟��Ty�驩!����^���\;��Ι������p,�ǔ���9�V�>WB��*���]�����]9fE:}��n��^�"�9�j�\�lŎ�w:�a��3N�}e�FBB�rӴ�~lĦL����5���w8뵄����GPڇ�*L(~�tm^��� ���&a~�9Z�	K�Ո��5S7�Z���LU��56�&PRcˣc�=8!�K��İ�Ƞ�Y�ሔ���47�0��b4�|�(VO93�� ��`�[����B���ή���r
N����r��P�}ʟ=��6�B��Ѻf>.�.l�}x:�@f�Gi���ZL	�DO_�|O�VO�I�XR\��q��{�۳��1ƅ�=���i�D0����f�.��H=^1�3��a%L���W��,f�,�l�.`��H�y�1p=�}�,g�HЁ���_��uy'^��>�5h��Y��$���I�[#%sh�,��t��wK��]/@�!��ګ�h����'�E�F+�?����#2 l��&`կ�@-7ql˖�S/6''َ�	���]9qy<���D���1�U�m�P�U����8|�
����O5�ALȶ����>V+I�&C	o^�fU��C�Y�}��оz������U�����F�y��/�,���^����@U�*�
��w��n���Y�*M�U�J���y
� �O�#�ʳfb���&4h�i�ޤI0�f���N���ҡ:��V:��Bk�>�q.�/{��8'BK�˥6*C����B}�G���|�L�v:)Ӫ� �H���J�?c1.�������q�f�m�����fs�y;�Z�`p�7
x�A[���� �vHS ����_�P�ȭ�m��8�������q�Tq��t�@V���}a{��dn��&�a� ��=HJ��ޚ��M䍧�D6���&gg]l�Ie1����wQ��Eo���c�[�+��a\��_$7a���Û�X�5��@���m�C��=�&����̀���lΊ�QF���Q��.Ǻ��_��Ǜ��	f��-�-غ��YH�H`�p�o�G�_�T��`+���(g���Ꞻ���&��F�����le{&��z9�e�>~tz��7c���{����6[�ˈ"}����}�`޲�t���㛾�qX#(�χu�����r���j��E�A�V`V+���G=n	�Mcø>f�i̼�4��Qb�7������vVv��Δ�Z2̫#�j�F�YЛ�KDɔ��5*�Y����b�|�=�2��q$�=wUS���E	��)f �a ~�rP�����7O�l�bj1��pw�k�z�E��'�DU���Ks�������6P}����L�jpb�����+4�ܖ3g|d�K0�I�r��ӁРz�^	�:c�$���0��¤;Wہ�+l�4�<X g���Y2�&+R�pH�K�"���9 p+o��,Z	��_̠�~dx�-�ϩ/z�ͶO�+����6��-�t@���h�\��e~���k;�2��m�5��ONκ��ˊ]*Ru���'�Xf"�^Ju`��RkD�|�*��7��{}�hDM%��s%P�:��p�f�`�Yg��I=X���_�,�L"�:ڗ�$���.^�|'S�����R�?9P'��NǁQ�He��IN�G�@�ѵ����.���w��H�����g�I]��y�x����R��`T*$���xM�7.��&��!�/X>�D|34��S�Wi~m<
-�JU����9MJ�7T_��.��ۉA�ս��;
��_\�Tu�7�|��0?/4��e��P�_���\��Efq��֜8߶}I�hٚ�eO�J�!l\�%�.�
��7�%��w�j��h/X�l�w��@���� 8gnJX_q.��v)�`'5p%�n�����Pr�^͔Y��V��y)#]V����95�-����H�%�:?�z�,�l�(���;�WT?ˆ����$��A�nt�,	u�����xp=��� uw3�Y��ID��A�t���ڙ�!�$��z���Bw�7��hܯ�^��ʂ^�Iʲ���J���3{ʡk���/��g˧��k;����{ѵ��V��e���-�z���]�Q\��1�vdbo)����j�����E�a�@�"W������M�!��m�OL�l���)f��Nu�6L�6�+��zN?��lD:m�-�p�[m� ��f�W�v�#��y��������	s�,��'�&����D�/u�	c	E3�p)kZa%B�}evL�D/d79Ć������C��.i>�^кԏ��]x0:Χ��7���	/,|֎�$F�ɧ܂>��Z��V�pʗ]�ϖ@nm[�i�=Z.�̰�����B�
$����2�5k�X�Q G2ك��\�Vv���=�6�����{S�5����ZX��}���0>�6+�Qi(�\��<b},HО����'�шZ�t���>=�,[��8��b�Uk<4�ݫ׽2�� �C���N�z�6h�pJ�a2��æ��8R��D���A��Q�CSoU4��,�H�77��"�3^<�E�wYi�Ƣ���q'�9`pL�4�X~��
Ә'��32(&d�w��j�շ�W��tƑ=�/�ĳ
��F]�>J_��u�f�<U"ǰch�_�~�=�H&f���[0����Kocqv����̦\2�-���)_i��έf��^V�]�<a�[+T�(X�d
g!̺�/,k5��e�=�Q��xiOU�Y�'&�����hX�;k�lJ�%%�3JO#4�#|����������_�AK���v���a��`����{����*c�L4J��\u�8�y$yz���1��|�r
�SX;o�AofK�h?"8۞\9U`��Jo��ĝ�Mv��a�1O�[B֜?zK���A��c�l��vw'k�/������p�A�Z>S����&Nm�e��+�ӝ�.;���K̪�oct�P3W�+�߭�Yn�5�ք7�Z��[�3��,w��2=Vd݁�hϴ
�RRd^i.�a�t�zM�?��T�O�J�!>$GL>�I�L;q����Xћ�B���
m�V���pH��D��u䱾ҍH�OOb��	<�u1���e�!�Pp�Fr>���_��}<��(ɿ9d�@j	�n�]���g�M�@)�5A���p� ���+���A=��%�7i��{�^+����scD�Je�B�&�No�L��Xr�#��(����Z��~�A~��r�J2Y�>$Nd��L�
�%��I	��>��|0�R�2�G�F�]����=����Z/G@QH&b�0�z3�N�E
�?�kO�^�U-�����܃���^{�7'��"\r�d��{�p� ���N̳}e�cA[TTƆ'���0�U���#�x��|%�J,��'�D��q�3 �l��XM1*kd���A, �*�}�����i\���I�%�^t�r��.	�v���O%4�rL9,�4u�s�ц�M�_f�%gv������kۥΊw�i1�U>����)m�ό��g��t�u�[�KS�Q�hz �Bj|u���y�l���)Ŀ��,Q�{�6j�lb�����a_�崄̅sRu�:�=� �d�oND|�����>嘛��h���m�yAu��~0}��=o�L�!9�V��w�jD��n��g���_T�#m�l9�ܹC�Э1,0me������Çrb�R���5Ӽ2	��3�	(*��@1��)!���ȣ'�
3�c��|.���XV/�Z��Ԏ2�Y8VS��U�M��.�f0D��k�C�c
�յH���i�I �9	��j7��~�硕�Σ�/�u �+{|Z��w�� �_7�'�\��l�
w�����A��秵[�BG�o��8��Ʊ�#����\[܊�ECg��->��\�[�.4y�K%,���y�gwj{��u�۾B/�X�kƩ��C�(	v�"E|���:0���6�����1{�}���c���t��+�Q(Y�	&�yF?l��Ӗsxzj�*q�P������@KMR�g<[��#��Z.���g��9DJr_�8��q�1ݡ2���b�o�R뎾0���$f_.�f��+��2AbjL�l�R}*+��eU�qF�4(_�;�}|ä9=~=&�;+G�7�����lP|x�������Ձ��+���)4M@���;v��F������9p�f�2���l�H�^�����a�d�)3�Έ����h:	ɡ���̄���1s�HA��>�/Э�$A����d��	�:f'`���e<��"��,k�=0�P�kxqhJ��Q��.�+���k>: AP��5�H�,@�5�W�+꿳���>���
��ط��Fuha��N�R�lD��Z&6���.�!Q���#m�{ف@���A�'H?L����1��ܻ�Mb��R����劷�m���1�ם�[\릒m3��G5+N�m���ڜ�S�E�&����N4��i5�����ީ8I�]�d��$��PgXr�s�)� �%����D'j��)J���� �-���b��Lw�Z��_�qč���8[�ix��3�;�#��L�>37B�A������Ey��ژ:Q�.�;8 �	W��x��&��=��p��»z�i�1i-�XG���mlo���.E[�Y'��6E�W.Au�h�Д����1�ʲ������j_
��Z:DG�jx�fy�ԅr���+u�l������eKtHP^84���^%`�Џ�A]'v��ⵊ�*�����#:��yDA
�̦j�w�о�����e�]��K��n!?3�8�իp�B~��ӇU+�QU~���c`������e��V1�7�0���^�j�l�<T;��Hq+M�m�����d��"E���*.t%�͒,S�m�������0�|މ*���^w�!��1\t�_��K��p�{=�� ���6�(�5��
�i���eV��X�]�=��-�L��r
�u�d{¢`���?��YN�a^:J=$$�Ă_ڧ��L�������jAx���� ��@�ri,]M9��B�%k���u�� �;Xjo a\�$���������X��n�Ɣ>η�F�p�Dվ�ճǝ���'GO��))��	[�'�w*Ɯ�<e��5Gt����/%���c��3��v�=�&�P�^��;ZhկH���۽'�f�٣������ �����AA�g�����Er~����M�Z#dJT5w�xl����A*���2��Oe8}����(J�,SI����S)M�k��	�����|�v!�3��h�aL��)�~��ߏ��jo���+^�f
�8)�5��ʽ��ڤ���KU�7�Ղϥ;����(l���U ��7�g�t��fǴW{��{��' NM�z��A$��́���K&ԍ9�B�Թ�u�<��hCWΤ��Wi�
&�-ڭd\HփH&"�{��}�Pӣ��#��%�1�w���\~t���q�����z7b�	��b��^���|�*&��W���[��w�KPk�#Af x=)_��)�3��ڵ�Yc��^2��'�_x��!�|�l5'��@zz��-�jtbi�*e����r���E��j��N��(��JҵT�n�Jn&;5�1�����&R�`�0�@
=F$w�}E�:��@�O{�fY����R��p���Ñ͌F�Sm0�<6��ϖ�0�#4�s	r+���rŔ��rgx
bE[qJ4T�L�З-hQ�cq��!ۤ��|uA�H����{1H�!J �-��k]|���o����5���W�	�/
U�
o�k��3	L�@t�,`��ĭSTNskƿx���}��v��f<6�X�Sj"]�2g����P���V �����c�+i�y<�س>,c�r��$�f���b:p���K�i���B+��T�����驊6��3#�=��W�;vz�Q�����Ի���'f]�aXý�=���x���!Y툇1�ڽȁ�\f�q����@]�~Ob�F�ǒ=�_��N0s�EO�J�fFw]\��k9r��2��l�/�4�9�nֶ�*.�d)�~⪃�S$��k�YBB����g�
v,Ɨo��l��\��Ԑ[ ����*���d�w׏u�Q���� ò�w�-���KMM�>��QA�o	�&�_ȈƆ8~�2Əg���v�~l/�v/H��n"�8�H�J�$�k數���P=uׇp�)'m��hX;���u̓(��<Z��i����\���o�k�+�M�A�@BƋ��JJ�hO��k#)���Uu]瓍k��Ѣ���M�$B�wV�Z����)���.A�t�R�i�wP}���"�Q)q�6��q]���>{� �>*V���\Z͜�om4Q�ռ���rx>�sS�-@�����IZ�c��s%�v��j��B<�v�S:9-�g�.���&��,�G6�`�v�_�I���EC�|�;��d�7� ܺ��՘����S�PlHM��{"ҋ��@W�{���y��(��=.Dx�G��}����)h��јҨ��\���6�����^e��B�#8��-m�Z�&�zq�ӎ:�~Q��n)��J����o�Ĩ��h]����������ȣ{,����(�2HcC�(o�3`�0�FEr���X�.�q��JC��Ls�Ҕ��>b¢���_d/��� m���쑘SS�(�~�p�;���=��ܹ֮n	�Wj�I+Ю�9s�6���U��'n+���0�:��l�֋څ�O ��'oW���; 7@ӻ�Ml̍�.�	x�l�n(��yk7�պB��;C�v�n��*���y�Gc�ۛ|2����ÛEsŝ���G-��1��3H�gw���C���n�=@{P���xb$.vr�Ψ�i�5�҄�`��ײ�Q�<ʢ�Ļb�^Q�&��"#�M_ɿ�f[\y:��F�د�x� �t��C�JJ�@>���mB�eBS�f��A߳�܏X ��_��b����aN�.�0k�Χ+�M���B@� �P� �Ӡ@�i���~������W0�/��25@??���W����O����D�{q�q�Ai\�?��4�-��b�5Y��s[�X���g��b� 1�J��U(>?��d�F2�	��OV �M�����_ϒ��	�b��ԓ�[���РBUXׄ�=Y}�ʩ9Z���)�� ��.�)�y�޺�+Y~����LH��2ၼ� �����~��:��Cgb���5x�M���
�uk�K ��n(��N8�t��֢�@�bBt�}�_�3n�e�2��M.�-�ۏ�<x�4�'uF]�Cɚ��<�8�����܅}���Z/�P��CE\@_��|>д`�Ѿ�`z'�q�r$曨S[�9���<|N��$^K''�c��J$: ~�ǟ�H���_HeҶ�PfS����q{�##HOΤYJ�ul�J+�H����m�Ԥ
�f��x~�rOl��T�Wp��1��Xk��^}�¸��:�e��r5p7IPΡ��z=[�8��E2D��3�hz� �5����n�l�U��Pď��Jg�O���_*�%�,+��S(����H�G���G�\�*(���<�H��a;�� ���a
9 �vZ��)�I\��[�#0#r~ ���2k	�'��Y�̗���X��1�U02`M2� ��>o�f����0���-�E͋�������}2��k�@�#��g�
���M�������t�1�m����0�N���'T?k���6��d,~1�T��������$�-���&Y�EZn�h}��i��ޜ ���El���W����V��kHZY�qɚ�^M�����P���px.�M�O#C=�W0�O�������|#��u�Ht�I���<s��} �J�?¹q}_�]O�(=Ȃ�X;LڝHn��Z��^��m�k��=*i[_�N�Tzl��;��>�#Q��C������ �E����9d vP-��4�P�8�؏.q+�7q)�ރ��n�	G�^�ɞ�.'!�v5��ga��	���rԹ�F����*۸4���E3�8�ZP����x�Z�U�9�\�f�p�JFs>�a���*�Ou��t�����G��<= CI4i�#b/Tl�_�m�pAW94]ğ�J?���W�t{\�NwD���}��	�����l��5G�#���J�0@��K[?��
W���m�~	��(�c�k�z}@)�4�N�Y�~TV1�c��bzHEi1��7OGz�ao��Q�S�+1�k �M��V����T��V�-�����l�w�����R]`Ϊ6�E��(��n]O2~~���z�����[��S�M��V�c
Q`t/��J���	��uo���^>�<��P�0���w1d�a�쩗GŪ����h
$Y���#7sg�/����\.v��hi�W+�P�ɂPр��/���6���ݱ����o�Ǐ��G���R{N�d��`����0��q̏G�B��1ޖ;�L��a_��v/�疙6��Yak�E6�w����w#,֣���+`�0�^��8j{i%��.俖��dK �3���1�}��Ю��1q���-��JR�u�m�Å�Jֱ��[kMy�v? ��fK�x���E`f[9[�������z�x�<�Z�L~aZ��@ "��9Gr6���G�p�Q���ņ���'K
�v��+=VZG������0W� C�E	M�������.娟l�3l��Ɛ �c�<���yJ��]��+.qI'.����-<'>�>$$q�/����7< F)�?�@�u��UF'=�y��O��3M�	�j4���9��2;RwE����uq�����`Qڝz���#!^�̡Cr�6��{j���뚳N��<u���hĪ �ԕ��<��6�*سR;5�#�0ur\fQ�L�F�+<7�yJF�j�?|�շw����D|P�N��U��9�h�GV/�yJWx�������)B�\ލ$a���ǟ]��^q|`�w�������(�o��.1Wm ��jvFL��`�[pEn�f���[�<�f%�Z
�P̚h��P���!� j,��J�)%���~͢d*O��F^���)r{�_�V r9GQ���ǐ�<ߔ�45���A��?�\�y0<�
�/	Ѧ�x!���1p�@L���C˞����5ڂ��k�ZE��RZA��vwc,��P��s2�&��<[A}�8����.n��N��p�&�Wf�T�*�&��0���i��a%����^���{ߐ����>�0�G��8���7"-�ϲ�"V�Fбo���!ź�:��/�S̕���� -Y}ZB���NW�e-���g��\ �����+��$��0
"�1G��}5�?�[�O��<>���1�9���3�x˯��H�(�8*|b��=�QP{��QWޡ�Q����0���������P-�@'����.]q�����L��NާSu�44v퓍�Q�z��"�I�,��|U�8V�H�[g�X�(΂c��*�8`��c��g�����o��T�I�nŏ��D��j��w�7��Җ-B+?�2�h]yz�2|������B�D�d��8ӉJyM��OxlA���ғ�����Q��Y��DXVJQ���"tONX���O�,��|�;��q�F2��^�*%L|�}^���t.�|A��	��J����TX"\6A���iN>��P��ya��.AYGY��(�|&��z�l���@��@�%��<�;H�C2���O&!�V�xmO��J��e�Z}�����+Ӆ8��^1���'7C�k��	�`��j�b!Yf��W�X+�ƨ*)���"��Q��
&��ѭh^��o3�]t d6qф�xb���n ����.�|��`�r������c�,�R�Fp>F�����D��wo��C_Mz�؂�M�4`���'r���}��>O|�FHV;�c%	@��C��&��=�UF���A^3��c��qj;�0�)������W|�oQ�e ~��w^NE�( �?�6u���@m�.L2<g��a�!��:@�Oj	�3>9r]=:-ӛk�tڲld��ɑ8���p�m�����>�j^1���]�Hw��k`��h����I⠐ӎY����F�$x���L��w
�T�ʹ��W�k�K�a�d*�&.�¸�w��,4ʒ���8�@C�-�� ݘ����1o���)@Q˅��AW���-5.K��ݲ�Zː7���Jy������ć�<;�dyn�h���S��m����� ���|�-�,�R-U�vǥ�����_���[pO����.������ί�˘7��Vh�V,�KT�p���ul&N��,y������|��>p�� �1��z���q;y~,�L��z�E�_���Z̘Zz����������>��<m:i�q���N�1�z���G1P���5#�w�:7`���zͿ�սfZ!�2�i���3���kzY��٪�6�UD��u(fC+�0��0��,��[��1/�2��sK����£�~��b�>e��Rr�Ԥ�xb����g0A�~��j���-�+9`m\2�yIx��w)˶9i��}8N��0;5�ݶ4q���c!��)��Dw<J�z�����3[�CIWKCg�D�J�d���Q[�e ��� Gy=.�$�P�*x^�Gp�a��:X�W�~R��aak��r10RWa(l�9m�49N�u�@����>L���TaL>�� �\ҭ/gό��t4��#�<w@*#x6�� Q��~ՕD9��@�2Q��pPx�`=(���_yz	=���2���d�m���,�t�S�㼙�k��o'��Eѓ;t�Ȁh�.��?d�X+*_nD8���ħi O�=5<�S���H�7c�]���6��W�#�֧\X�5�Qr�����������a�.ĕ���[��Id�ɦJB#FI j\#��e����-���f�9Y%����O��?����d�Y�fH�&��BRD�GP��������c�G�����V=�B2׿�f=�y��9�q�������>���W�ĝ�ܝ�vЧ�H�pVP99�0N�m֧��n3m^hΝ�v���C/ؔt��!�H�����[�dedp�?���qO���`.ކ]�"����R"����}f�˯���B�7!������jaf��,�Nw��J6�"+����RuM�)r^���[id#i��G�;	�fI��UQ��tQ5m�e<{����P�;1XK!uv
�1�j�$L. �q	�s���B����0�=�,��'E�'�����½��5��@�Ĺ�Uz	R��h,�"11�s����8���r��l����j��0��suF99���������[f�^X���ϓ�-�$@�x�g��a6F��Õ3J�`eh[�FU��7P�r�qS<�����2y�R'�l�1b~)%
�3�HJpb�K�e'�7:P��L�LY胔i��
Rm]ŧE˺��a�Z�.�����ڼS��v��g�J���A����>�h�3��2��>ޑ�Z�*EqQPo�w�H������He��2�K]{��P��<V������g�F�b%��2Ԏ+�*Z����o������GN�r8k�N���Ys�.k�w���m��1y�p�6vp�`V���gS�/�\����5��l+(��R�@���3s}�_qri_Z� MH~ýz�8s�̾���1��S"v��=g�qT��9��?�7�7j<L��L2�'ƶ���S���a�ʠ��dA��̃������ag��ĉ�54��{�x���W�8�|W��XJf�C\β+����u�6Gqj�p<c��2)��G���k�BX9���ܝ$T��CL���)�!��Gj/߰s��m�02�;R��@����m~0�$)K�'w� �dY_zE�݋$�`���	^�Ik�B<9�ڶ>^�� Km�5�W����u��eC8t�g��H.8�H��>�%jW��5��Aݐ�R~&n�s��(�28.��j�C����B��Z^?'t�Q�6.D�j]ZH�ɠeiŰ}d��B�fY����pDx��%�)���� ?��K�{ ϽN�n�-�BɃHv��4Kҏ�CѴ���g8sLs����-�,����c!*��/�ν x
�)T��7�P._.`D1 ,M��\����	��$ -�,3�1Cq7���Ǽ���mog�sc�x���J���,��ֿ͡����/:�*�n����>9pl�
�U[I�J묈�$��O�'�n���U���?h[QI���_$�X�4^����B�6������s�(���&J�]�;�g)��b�߂c�-�u`�p���ޒ�Iʍn�����ba�!fү�>iAެ�F��`}}��I36O��|�3WDxF�u�E��[ߋO���bt��¬�[dn�
�Tv�x X���)t4|�ـ����Ji�&�P��%�9� ��`����>އ
c�h�bĶ�N�Vl����ie#��ոh{�Y�]4������"l��T��vB����&[�3
����W��b� j`��J� ��\KI�9��O<ER�Ѫ6 ksg8���j����!��o���t�d�N�. �O�:�$��X�q��E�"`�K
�
+:��!����1\�կ��_�a��&sސ9Ҕ�p�eZ�i�F�Y�~+K��&��0ɯ)�=�֨�H�������.� �����^&��3��ڟ�v�M[�x�mi�X��\���U��r&@Hf�1��.{�s�E�=�7fxt���A"Cڮ���T��������1?�����FB�|�Q����x��)����q"�d�����J�O{�y~�3w�JHZ;.��1a.	$�$���Զ��c�s�a���h3 ��O�a�0���HR0NN�ph�?�i-��/8w�#�g�}����A��$����j��.���YIY��X���rہH��T>m�0�S��Ե��ȭ���J�㱨uzh��Z��sA�k�!,�s?�X�V)��_a��L}wl	o�5'���%W����5��W�:�L�D��yAD+����+m�XٔX�-7��N
�ng,���<T�1eVa=�K�xN���\�Ԇ���/�4�C�O쀗��C�T)䒧$�q�O������ ���GTT�Ir��OpX��gF��H����D�����d�(�ay1��_�IbT�mպwG�˃��fY�_��6��¨,�&�"�c�>{�p@Z��:�o����z���$���`��_��p�Å��^	�ק�J�y����f�[�L.�`r,�y��Ē\i��q������1�����O�s��ź�
W6�-$�ÅC<X&hRG�n��ԥ�,1��y�f�us����?"B���e����
��rDv=����ѝs䐈��dP���]]�-|��]��g�k��v�F����@U���-'d��½� �:xk��GR�9�z\xm]n�ۖP!�c���DA���h�$��F�"nꖛ���vt8���6>�~��y����x��'o�%���h�dh��� �y-��fyOAf�B��9�2yy/�`F����(�-�u� ��I��Ox��-�����:�H��C�B�ch�H!��8Ip�n�i�h z*��������Y���6ڽ��
j5���ϔh�䞭�3T�"X��]�D���V�9�:�<�GV
�{�BE7��U�
�>I��6+*��ʩ��g�#'�b�3:�_�4xi�@]@��XǞ����V��8�a4��)��/"��m�:�G�2�Pi��!^Ƒ�J�T���f~��_r��UBF** ���^��z,J��1}�����s[�@�O��և�-���z�2eё� ��~�����,ǰ$?�{8�A�V��Z���$_���oE0�H(�!� L���k�4ǆ� �Eq��:�I�QSPI���+0=j �[�� ��V�Q����]Ƚ�D��5C�q��#�R��,�m�`HD�"����h�1j.c��!~�ٮ6L�~��n�Q�'i�r��*��}O%�t'`���<#�R����
�L�	�LB�RL{��Y���V8�niQ+��I.��9G��7'H5����5�'?���!�U��gfg�D?�V�)�� ����f�������Q���g�����t`�&�<�_�J�p-mvu�Q��93�r���z�4`޵�19&7�Zآ��+Ar�ؠA�W�7�HF%�*���&�}{�>ɺJFv������O�66���af������^�r⨽U`���^*��cs?-�"��<B���!�u�N4M�~��Kb @���:2��k ��&2=^�z���ot�͋���%'�SA��L�S"b�014 �����_*���|���͓�?K:Tc;2�{~|��� �r��@��$���s�g$rM:���zfE���@�;Z�N�i���F@���	.WCa�8����N,�]��ny^i���j�<�p� >eA	ձ�\�#8x�M(}z1�r��=�8�}��I�~_��$<��:��r�,@��N4�G�n�Xz���`�jz%F���<\t��~d����Ǵ,h�7ϝ����Ն9rf�^3_	����4#W:���b%V��{��2�D<l����ҡ��&2/�"��;{`�io���?2��)"��u��i����|���%���^��1n��ψ}��na�y�Ο������2*1o1����\-%�\LU_jk���vnyg��)�6�]���Y
�����y��p�ײ�e�F��k��iAB*�j����&FLG��bm��3v�1蒫y�K��x�j=��sX�?m6o$��*��<X
ptH9��?���������6^�L���3�ͺ&�T�Rz��-�cb��>(#|pjb t�tѯ#�F���OV'�-Z�PuJ!���p[�v-q����y=��|��(������=w�h��'b��u �_R3%%�j)�<=�,�e��� 6�
��s2Tq/�����`#�Gy�7?T�Tv�~�bĠ$.�@�"��+���]��ڒ�k�m�­�����>O������u'���}�N<6@Zb�}F� �����9�"ް$."}Z܉�If�n�զ�z�|�w.=a�ʓ���B"�޺_>�wz�
	�BC�~��8�߷��]8^|����i��Y$��ׇ&3~lP��\=oN�僭�t�z�˧|O��C��u�X`0Ipf�x�xk��z˝��o���賈�!MK����n���v��(l/�d��_%���P�mD�'A!� �m3,�L�S��|�,NT+d���l�{&�h}ր�Z������x�p�VeD5�x��@!����J2�#�\����+�kK�f�Ǭt��(���Q�t(zj^ .E�u�q��c.X{K�n��.#����t��c��'$I�i?�a���`���T��@^J!
�����6��c�e.�+�~٥n��!�MYҔ�6$��YQVׇ,[N�q��6��*�~}����u3)H��p�_�X�7��n\1������I�:���w�ʤ�V���o
��[��p˟��D%��%D�o�ȳ�H��e�C��*����2�vS��)ҕ�ϥ����M	%!'�Gڷ�T?g�U��d�P�B\��)��SD�F��\Am<�f/���[+�J�K��eBYbn�{���cH����	Oa�=:��uH�g{������(�{��J5fGI$9ĺo�}�\�W!}�y�O�q5J���i[���$�%o�N|~D�1M�t�������?4��M�͖�}���K&�
�ɪ^4V|�9&�`�&&*��O��%���N��e6y�I�+]��d��e;T�����F�`4` �S g�C�߰������W�-}1w+�ZA�x=_ƛ8���sj�˓[����#����n�n�=Z��A�3��Xrj�K9� �l��O���i}F/^Y���B9v���-ҎY��Wx+�sC5��˳���lh��m"�r*@G�d�Z40���%�f�ܒY'��KB���gei�+�Rn�8�z��X���2<�;<os����8�5L��6~�U,RO����-����9����U�8�3�#=�������\y����{hu�Q�o�]i)�~}"� U�i�*Rc�{�w�g�(��I0�j���������#������-�1-je�8ER�v�-Zk$��{y��ƒ�گ>!vO6���'T���S��;H(t��/+�[��x8g�P��^F���a�F{8oiB�B鬣�X��R|Ef�)Q���5�а�$�8�"��$��D�{��?��;%u���<�;؅嚪��"��^�9;��r��>��L����m|�RyS�N�O����k
����=ξFH��Q7�ﮂ2�H���P��M�d_���_~���Q1K5�ϋ�}	S{
,i��n���1W��M���lௌ_�$����"F�`���V�ŋ�,�Ƹ(�a�iZ�@���(�3�G�|n��)�Lm����c��=/�B�_��'lI�K��y?Q���%�hx�ߨ,�W��ٍ��� �3�o�Z�y�ol+gTm�Ew�~Z��<���|��v
�U�Ro���=?gEӄ�.���'�ʥ��j�o�n��}a�A�0�՞s���'�gl�E0�f��]���r�R���eDe�#�$E>�g0��&� zg�߯�O�͝�y�����:gQ|\uP.��v�c���k�`�?V��p�(�3�I��8t q�hu6^�����=��U��xM���¸�BBN�ð�y��>r=s�e̼K��r6��}~&�V�^���i�-c4x������·�Of�	sTj>�=kƖN=pӘ�U+{��[g߆p$۟��I���qT/���N �Ѵ�(L�	2�b��Z�4�9�/��]rL��#6C�;�qc�^�_0w�zD��=OiF0�e���ݤ�aj��c�
�!�F��T5�\.�|� ؙk�S1]�g3ΪG�Y+����;�#Ǳ�?�E��2Os���AfH1��quiy���M�m*0����(Cf+UE���%]�~���=K� �R]����V�x譀�ĕk��"��yŇ����%Ƕt|�>�MhŁ�Ix~mE^�Dq�(��t��B�(NF�"��3�g����M������
�����B�+ɱ�)й 	�e��Is3T������
x�M�����M׎�CUK�0Z�i�fl&`��[���*�v�1��z��ծ��[��<Y�Q��w����O��y�k[|��1z�?�]�B.ڴ��I�k� �����C��',��[�c� [����I�w*d������O���@�k|����|��׷	��휴O3D+�>ck^������]�$4�K�< f�lNlq�1�n�|+�sډ:����D����Gm��r�a�ET�a�����Bw�}pG���Gꄅ.jS�]�e����q�ќ�Ec;TS:�+�i��7�`�D��-'���e�dw�Ա���IhRB��08z����2���uҏ�ڠ6,ysn�!6O��^WW>�ӛ�� ��9g|���{�{>'�\	kϿ�fP�,��8���ꘜ�z@d��	��BG��Uf�ux����*�e�QH9X* -�C:��6�Q� g^�F̷7�m@���GI�_�`%���a��v1�!��������3~�ln���-��+�b���V6���:����n[�x8 #����'㑡��=Qh6?�a%�&�dÆ =u>[��6�֬�IY(�y/�W���i�r1�v%�T����>P?���I�x�[�O�d�i�Rn\7�v/�5�"aE+֙/��Rc��d�zI�)ر���q��+9�����0E���;�D+_��4!p,f+[�����/c7/�9�כٽ��Ѹ{D������$��b-K��g�+�^�b�m��Rj} t��ޫ�*߅Ǹ~���qɕo�D�ܢj#���J^��<'�F	�������{�Eh�9
���(X�8x�Pڇ"����N�V�RM���1��Y�ݜNj���ׅ�/��vksF�FH�z5>?���n�~�}�LZT�Kl� g��\ZO���Y�����Q:�EvP�;t,����Z�b��#\i���z�>n�f�>����\������i��}���W?֥�G�?���m�T��F9,줹#_���^�
LR�B;�1tK�t�"tV�e��S�+�Gʂ.�����a�d^�Jep$���*��I�	��ﭢ����q����w��P*��,\��QUk�@䒾����5�?�Rh� 	Ȧ�23��i��(qy���2����OV���o*xuw �f���[�A�k��P��B Y��ƻ;���U�+���՚�l:7���*dp��������dN~������?�N�̐���u҆j��*��ۄ@`��e.��eI�֢�,���*��L��+�~�Ybg�Ez�L����5<��{��^��p��(�ޢ\�p�m!�Jr����.�r�'k�7 (�n8XB�Uu�Bad�\3��p<�ڼC[��	����1�z��/��۾֢]؆�%�s)u�y�a�s�g��J���M��վf ����]l��	7�Y;�)!�I�7�7�VF<9q{�~c�ׯ�p}����λ����X-��L�J
���1
(CTOo���3�n��?ո�ٹ�;~NM�k�]��e�]�s�����&�+HGS`xtdz����fu@�BYpvuB���t-����G��tO��ۮ���nq�(�Z%i)@�K����N���U��#/㫻���%�+k�I����eb�]5�۶A�8�����zq��q.7RؘL{�/�K�tb�j��ON�r�f��&,֌�{���0�7�� �.��s�Q��f�?�s�iyE{�!ɡ�>1���1���e:h��d����%J�iM'���¡�V���UM���V�,��P���b�QᲙz�����h�͂�¦aDi�Pc����Q͊��K�&��&Q)��┪�O����4��C	5�8,l�q�#0S�]�	���u4�Ǘ�K�b���I�=�;<�����z|��ԛl��@��v�Il�0$��4�u�q��ۚkb��h��{�u=A���>bR�@.?����/3|�$%��|��{3��n�_�=���#؍&�Y��sR�Տ�D�C߼�vd}�j`��^Lghh��x)@e&T !�u+5t[kO��+�z��Q���h�d4�fda�2!t���� �6Z��ڒOk�i�,�0xʏ�>�{�3��rt$�>0$��r|�W��q�Vf�ճ~mߤ�k@B�����;���ܝ7�e������1�ڤ��ǉ^�0���D�F�<G-T��(�P�����yc
���f̄�Ħgg�ˉ�x� =g�h5;��ۚ��h��~X�z'S=U���Z��K�#��\�����}U�ޢ�"-���^��|G�8(>�u.��G�L��`W��q�3̥=ʮ��qۧ�n5R�6l�g�$���}a�l��;=kP�q���c�(^-�84�A�,�L�����߇��˞������n�."t�pt*4$��{f�W�K{>P��O>�~:>?ҿ�D�ٜ+���8X�q��j2!�����q�M�K�#=߭F�R�k�ۄhT��1+�*i#�}x"L���H���L��~1>�w�١�cS�|��ʒ�:�s��A#�i���ң�9�Z���5�M�ʆ����X�!���{����� �d��ZB�A�(h:�؅�`�u���:9\�>�w��}��\o��}w;�%�=��sJ_l���ߺ�xppHG뛼B���0����A�r�{x����# �l����/�	�<le�s/�v(�o�tYJ� ����\L���9�g&le)/��;�X���)�wQ�p�:~�gJ"��diDܕf�+s���[�q���O����Y��r�� �q$OG�8�!)¯8-���y�g��0`#�=�!�@�;�Q��Y����{B��睴�����d���[�bo�;��;��f��zS�%�|�r�y�J�./0��>�� ���L�� m�jA(��
�Q�t�BK������9o���
�@����:��,ܔȎ��)S��
3\��[.Z�;�(]�q ��
\�<V��� �ŝ 9FŅAf����3}份�Յ��!������h
�����eb�f�a�*��R/KVB/ʄ�G�7�дi�R��������	5VR�mcK�6)��-�/$�O��o{@���Tg���6��E2���)�rMS(᯸c Yt&�to\B�~ߘ$�v��l���I��)O��|�6��3
FZK��;��M���z�m>����=d�:n%Ъc�������]�I���~�hh�pU�c~$}K��2�Ѽ��ooU�ǆMf��p�ʿ��1��GW�>4��w)7L�R���m�N�-ܝ�8�3�U]�iKG�-���������|6�f�����f�l?SO�@#�JJ�����ո�8]/:�$o�<�B�u�
~В�n̅�V+vfˀ���?$�2��-�Y���.˸��a@cc�a�Qh�Owk�h�����|6�roP&��J�$D�47t��j�b�H4j�,Vѩ���3Rl�K�����N�ҏ���L��ߟ.r��(WN���\�M��k�d�x>a����j��!�ƣxf`ՊJ^?����w�e�b�En�괂�~�R8F��\��_ں2�}𦘖��]
[e�>i'�[�fޚ���T�-�S��1��ۖ�Y��.��E=]
&�Ŵ�6�{ء	0͓M�����(����sb��~��ZOI�c�w�8�-66�����V�Rϫ��AAym�����e0u���}Sx��m�#�R�� lp��!;-a����TE�h����`~纐4�3N�uR����Bc�[Y��7����8�C[���U��?�ug��=VL\�rh��]Ʌ�N�L�M1j�}~�n�@��B�(�)^��G&@�6�c��u�fV�W�����AF���^d�^!G�z��5LX�3˸��y���c�����`j1{�B�z^ ��nW�`#P������2�C������ �����Iw&J\�U���P��0�5�+���\O�
����R�5pT���=X�%���ev3���� ;Ԗjk �=��U���c�`�YI�~��%��(����Þ0(�"�����&���~�D/x�iZ�oUa���l��L�| ��´� �*'z�E-:_��N^��j�{���o����Nd@:��+�eru@���J��M� �&�8Zmj_��-��Qd�.˪7��X1�,q�� ��������:�ί2/�?؏����q���a2���wFW�?	w��E�����fe]�#���gu:FH�UM6ѹ-��s2)e�Ԓ�\���Ϝ�f'V��`PO8�SA�B`gh����Hno�B~��ͤ`	���
�����$$�`����7�눙@�Ԛ�������u#��`IB�X6_K�� �f��WT󗻥�_�Y�Ћ�.�m��N�i�g�c+�$�Z��t���%��l�A� _ypB��a
�6P#�Y��𺣱������hI�����e�7�-�&��28�S�>����(�˧��Ar�/�"u��ۿ������$p�;��'���Bz�L/+8%�l�KM���DQH1����(&+����v(�{�šሃ�T�#���UGO�?`��s���B��Ԃ�
v4o�ֲ�TL�"���h�~�-^xJ���Z3�-��`���3�#YU:���0���~�Ͻ Tb�b���綢`G�����k���jT ؘ��;[)�٤=�-/��`*(��Y_�_�/�&h�O0�#��K�*�~�Q�a����f����5�E�l�~��Ӆ��(����I���TP�F'=������
.�L�ssO�
����H�Q�����b.`�n�<��/�X��f���-��mS���s䃓/� ��?�bZXf�B��I� ���W��6�A�*��+?���H�(���
Ȗ��*�(����?����i*"Q�9� ��~X[������3�ț�B�[��!�p���7���26Ua#����/�Y�ڝ��&��jh����H��5U��j8Z�ӬDK�v_�?�p�"ᯖ�r$�Ek�q���)�;�x8�Z��M/+�$�bYͧ{������H75�~�9X[�24�c^R&�����c3΀�Xݒ;����"���h�r�d�� @���'�/�Q!��B3ng�oE�N�<�l�Gs��;�S�� ��;��{f�HY�Ej�GLMpk��������Ƭw�D0��.=�6;�.U2�H;�(?TZl���X�|G�u�ɟ�c2�H����u.������%ʀ��hP�,�V��AU���(�(l?9vW�Xǰ�__�VXm�' ��� \"�������}���6qZ�_c������C%+�8�l-.���&��VU۴2]T>d��:%o�-9�4��Ƚ�V�}3�X�>w�^�(OF3P��L���:�-�0d���m{8�M�
��.��"��t�齋+�b�A�d��`Ѥk{�6%K��)�[D�2��]P�*X��n)�*��P��\�q�l�ZN�ا���k*�?�6����$����AdGT`|�z�("�+�@�䤲���ٟk�ߊ�'\P��	�|�cF卵S�G�*���	�д����/n�F�c�Z�y�;; �k���9q'�	��FTP���$Rs���H�r�����@G��OI|�����.�?J|�dj�}�a�mN5a�{E%�^�kd��hw�:z�G=�O�[�T�[�U����hZ�fѷ%��--� x@����Q�$���ikO3�TU�M�A���$˱(��K�ɹ�Ԣ��_I�pW�J*��ґS�<�3fN��$����W�9�BN��F6����]��U��T6��ݕ�i cum�37t�K6�$�Iu��5_�3�*��U qٶɹ��j�B�qV?K�Ο�wU.���Ѷ��]O54��A �˕�{�?�u=����\ց٤�Q����CX�MV�� J�EÖ��>:�S(K��?����F����y���=Y��x��93�U��@'�0�f܅����.�U�a���A�X�E9"��Iib�y����z����������C���3���G��ڪ��I�aM�B�6�j�rs�߰�{+TM�������ZbqDo�YW1C��3'j^����t+,𨸇��L1$"ڃŚ�E��L����J�q��Rv��?&��4����j��ȷ/�ZI��us���`)���ٌ7�HyUG˲�寲r���b�ܺڤx
m@k�H������\	(���h9���4㳇���O�s�J�z�s=�oTw��]�$k����8���<z�^Ѯ1���ȹ�C�ybOZZ�l�e��!��1inϜZm�:{,���m��O[$jhg%7ؼ����5�)_E�_�WvΔB8���+�B�S�h��rϹ�K��hq,�	dC�;1��/�o�_)G?x��:��"�A����Mi���!�Ÿ�z�;���}�	�zf���Ȣ0&܈\��hi�4#�T0��/Ј����8ė�rѷ���-�G2�w�%��͇�T��O��(^���Ƚ�U���CPp�M�%��<r�2���H)�M[��z��R�P=y.g��qU��:�6tl˷n���D۴x,0��͡7$,�i���������gQ��
g%ڕY>~������������=8�".%
C��U#$"�lj�k� lݱG����#�h�\��#f�w��;V����Zs���ߔ��<�9������8�+v	������ݾ�b]�~�����^���E��sL�c�p�7*zו�e�@d�6�t㐰�u���A�.��S_8��we�_l����G�T��P����UZ)m;�z�4��!ÇO}��*�?s�"�_�f��~�I�i�kWH˨��MZP�:҈��Q:��&P�/H|6�4[k-�� (j��^�0M�t;z}���7!���F�D\�)H����j9,�=�����t�M]�%���m8[��r� �01��xH�{�-��r4Ae�I��L��dSN����΢��"@A���*!�6��ZQɐ��s,�0߲e����A?��9��=f�x��3,0k�|�L7_��1j���Hh��[x&�(�0�dMI+�*3jcyx�k�O��@,�JȬ�MnM�t� ���zW�o�	��}ͷ�0�����uޡO��7+*hI�l���o��l'h�r����^�"IcpV���2x>�l�6A0��d����u��2� j��k�5��(`����&��Ife�u��D�YL�%u�vb�����E��@�}i147��N��DJ� �^���E�o�%�-���S�љfh�~��p�W�X1Tm�ĳ
=�!.:����0�.Mg���Q�c�OI2��KY4����*~U���M)���&n�/X9����E�E
��i��/,��J.��Kc��Ć0���rL1�V�!ʦ�Ǯ�;D��-4�����,C�&((/���/����\b�� 뗠�O��m�Rt�!��XI�eV��\�2F!C��C]��J�Ud>3�<�~)�HxZ�J��5 y71f"��,l��My�ލW�Xv��=ڊ�ѥ����*�`���wWZ�v�>�S���8�� �� 	~�qr%>���������6Ov��\��J��C��$cdGM{ww����A��}��j�}OӊB��-��X�s���sYr����"9"Q�F#$�xZ"8#c�ae��zC|�.N*��2���Z�Uǅy�����~��w#��u��e;Q�����j\l��p��2rƋ8�rxW+-���:EZ��^�V>֏����E*�g�E��\��,�(�;��r�"��n2J�G�R"k����q�!n
���s�EM�:��p��{63aMza|jD
�O<
�X3��:q��9R<e�[W����,���6���/��&*X�P��)�N���h���Ř�p��E4����E&m��Z��@O�?JH�����bHm���as6B��B�]�h���O�<�_ށ��x�'��V��gg:A�A����6N�$�M�C(�������gκ��2�{��7��z!w��#LA�=�Hg���U1>nv3�<k���{����BP���6�#8l��K�}ڎ��{aq�JV��`|���G�����Ӥ��nT�s�D�;Wԭ_X@ ��	(D��m�#�i��~�Eq���{g3H�y��-�,N��et�����D�5і�)4������d��u�V?z�:-�T��e�Ó��4&)��ϒ4�1ܙ*홚P� �#c���H��E͎P���#v-��>�7Nr����}5R��	���LF�HD�8�`�-hzMԑ��Aj.1���*�`�L���_��7D@}�zfR�ph���МK(Z6:3a���`��Gc�j$N-��$������z_K\pU��#b�$�K�
��R�梜�Ӣ8��%��?���Ц����ޭE���O��ݦ�^	༄�j𙧴��	�͉��L�q��D��#I�Uz <ا,z8[kruT�\�$�:��	�cH<���
7Fi���-Ujt.�������DwO� ��6�18��3- IT-���5�ּ|I#@|��)#s�,̙�������l�=���O����Vo�M bM��>�������;��y����i��Ԥ�1��^hKd�w���<F�����?�z�������C�w�����H�CeUq�\N#�! �6=vj�<$C�����|O7-HFw�~���C�w4,�夋�u�&H�ڄ0fThirԷ@d޺������h�Sv�d06������>N\ά<�Ԋ5�� ;4g���R�\��*�-9x�x��ȴ�J��A-Z�?��籲+���~@�6H��FMuhqg�8��k��w��d�o%/��E�C��S1���4�(L>r���*$�[�b�o��1��Z��?���hn0H��t�� Qb��Sb�~�gr?+��ƚ��.�hDx
B��)�ؐ���:4�uȥz��dŗO���nŇ� �+r�8�Eň}�}ٿ���� ��_�������1���F�^��Q2��R�g��Y������� >�"n������⎛��Uk�ʶ�u�L�*�SL[�/}8Q|BST�$�����i����[b]~���Ix$5x���Ec��� ��5XƗ)�<@G�Y�m��i�떴r�+�E�~\!G��3S���4k�������Pf{�?dX��Z%��ȣB9'j_����S}������TJLT)� �ؓ�/���ջ�@B[�J΢\�r(��)�gS�L(JȽ1,Bq��~��Ά&� �������GvGՈ[@x��~^�?�F�;`N�f�鈬׻�)�ś��w�\
�B&<�NcQ��y[�c�vx֮�4V��?���bc��Oss�pmA�q4��v����e-��ÚN�>�8�j��VZ+۞F{����9V��BwKkUgO���v�����nS�6?;Qեj#`��^#�u���v3	�X�)��cZ]Ż^�Q�cw(��
m�:�?�:�\\ݡ��G{\�ٝc�)ݶ�p��@�� 9����@��R���4ɍ[wy�%[�N^~��ծJ���4���t΂��O5x��U�l��A���:�j�������_�O'��P�C��Fz�$��0�zt��zm�+�ْ�W����{��Zf8̥��V�w�|��]�k�K{�5��0_}}W��7���Y)��3� �:���EjA�n��y�?�Ω55�¢�;��41x��,����G��z��c>_8��#k9	�?	�L}t�2�Ka�A�ʲ��������V<u��c���X�Q�钉����C�T{q/W�th�P�	�Z��7'����ͭ���b'푕���Hő�����3����v�_�:�+�+Ւ\'���=�gqEa�"�#C���ZW�*�i�#n���ԕ+1nh�\ͳ�gX��Q8S�S��g ��k��T���C]tJw�v���n�T�%_�R�MU��hX��4ew���Z��Gx\�?槤z�L�x��*k��~���ۻ&|�e�}���j���������G1�
XU\TcR&��(��A@<�F�?��CĢi%�I��n�9����*c�`A	�>����c�$v��y��u���R>������d�ܲg�l��/+.I P����*��+�Fti�MdcV+QO���Z�7�2��^�(�.p'w���#S����k�*����xk������9��n�S-�
��̤��Eq	1�hA���*��ǹ
tG"��QF��b�!�N}s,�j�x��8XN�X.c|(�S-�C Uu7*�f�!9kd���z�+f[+00�@�%�3�H˽���P�kkƞ!�������\�Z�9o�1Ħcw=g+�������	E��X �������m�cs_iZ[,���t�	u�|)��(0���A[�M͕�������w�������߇֣,M��h����iĵ�6f}���_�p����ykPw?A�V�AE4��yÑ���,5����|ac���KN��>��L9ɖq����ޝ���h��i�A[�,�vr��Y�Ґ��m��S��z5R�P�AGhP%	D5y�}��׼�R[��b
��ȅO��]J��a1E:�����ۺ����d���c�&j�N!�؟^dA�:L�/A�1n�5�,`�KB����1�Jdƺ붂	M'	�!ɧ�9)>�no��T;�!	�lW\������0Gg*a�)��|��P�`�8���T�*N,�0�� ^+�nӿQ��[G��!�U+�j�#<q��;�M�x����K`�)�/h�WP�����t�� 8�CZ�ֿ%+��F�B�Wǲ}sҊ<#3���H�?NGª�Aq��a��إ�8�S�����6/�j��͈-T�체'�석!ڗ�����B��b2��.Fv8[5�$2߂f�s��J8���䬈z	���<&C�I$�m�'6nGkS��I^[y��
�Xt�+�^(�MÝHO|n��f!I@h��;���"�d�<���X��6�;��5WͰ�����<��3�p�E���g��l,���k�u�j�:>ݓ��!DY����+EX�\�׌��wih��@r��� (�Ɲ��M?�,�/?�2ځ��;	�_O��0
4S7�$zv�s�i�w��dw3����j����P��U+���'{f�2����vOP�xC#GU����g@X]	�e����cO������m!�֧�@k?��S߅��"��|S(�|���)�
�	>'A�mDSG��q]�)�����U��\ɬ^ ��>�ȻS��xS���vM�)�'��.\��QV�۹[���pf��U�z�A�!2ʂ�O�o�C�[��	�It���4�i:1"���u2�	�ө�u
n�)� �|,;r�����u��X[�#�;Wq�Ίc�ˉ�@�<3ù�e��iӝ*f�;1�I6v~���n�vs+��ӑb{�+��b��ی�����I0�'�s'`�uHh�౴�*q\�*ni��ß���"�L�ÂdHw�6NΤ��uא��y� t$�iNV�O�ϥP�"��/���x����z�?9�gT�x�p�5o|
y)�t�z�u1|����5�F��}x�&#-�I��f6�ԃ*7�{���R�e9ԛ�pqr~l�gҖ�e]�I�ZB�#^��n+�a�>|Y��"�O��&ŧiu:ۦ�&%#P����2���`�k�����T��כ����uڏ�!���H2$�GPw	3x�`�v�Wh2�E{Px���܇��i^���YESJ� ���p�+�F�:b
%��Wwm��9�����s�>:S	�`b�cYL \����X"�d7k��R���$j�b�>z�TԼ8�:\^��V�~����֤AL��)����N�v�H�n���s���R|_H��@�)�_|�,Ac	V������G���8a�Z$A�H~����}�k�js�JH-a$��2�{�!�o�x�|�㿇n�"7���wW�޹Uv{��G����ܱK��> x��>M�@���ɘl<�|X{���C�P�v��+�#gvYf��	�/ڃ�]��-;-Ɍn��U�x�Z�Xݧ�hG��qUA�v-��������E����:կљ=�p�+����f(�B�4ELK
�D��?��TtR��ֱ^[J���<��so�9��4��]�Fq�ҝQ7�������=8X ����'w8{vC�ڿ�z�d2(��Ed����,F2�7��Ƙ�����F�<�5��k��}���I��f�6I�.���&�4� ����� c��u���)�|�v~���e�ҲI���ޓ԰�i-6m�-��6��S��>gj�����R_�d��W�+���ܞ]ydq�l饗��<�"�l��(K�{>� s�tAq��A[��1GH�t5�ʺBЌ�1E��@�w;M��"ke�����@�F`�0�"��S��wdk���t���}��pA"��O51x��L%�Cc��&�T)�2[���]S�-�'��[�G���"���j��=P��i�KO�ǃ�`�~ W���~Fyc�bx�[RR��T� e�3�3m����_>�Ou����.I�4��%lCG�����{�"����IuIࡒogZ�K*x�_2�L�b�dߒ�\ w����,T�@A���2�]�8�S���ԋ���_o ����?���-�>�`ҾiƠhy!��g-�v�� ��ף��J�[#�O���,~C�*�2>4^Y����T�N�۬�h,���Oj���?I�Q��~�{�S�^E��Pa����*Tlsy2}����4�e�H~��w�{7��"��2]���Tͭ$*<ۍ��Hu�-	<�K�rJV�aq�L1�$r%ۀ�X< O�C]��W%�n���́�Ļ1��Ei���w��nt"��\��^�`u���jǉ�����܇k�Ty'�m�]����d��nOE��@쮲&��f���MV���?֔'�3������`�#u�����[3�ܬEL%�3�����ѢQ]j�O�����p�;�=��Y���%%F��KMy�jU���:����Nl��R��=��r�aiͬ\a`��⻘S��o;��@�t��1iڑ ��t0�T�jl�XV��4�
��NK��	���/�3�8���c�0��&�¯s����F��K��Xxl "�
�bݪ�eK;�l@��X��U��LJ���@M��,��['T�|���B�Fc �]�)�1�Na,�e���B�~�)��y�U����n�Md|iI�dނ@��@RS��qb6B���E�+@�d-�kyh-�2��l�8�{�]�ץy}!pP�vPE�O��L�/�� �6�w�c3�f,�h��LE�4a��Em�ǳ�p�x�N�hY+��]b�Ə�5q3���ˉ�fp�/1�Mz��ȱy�pI�Z�#��r���]#��e��$v$�"��4Q�=I!�$��U"$İ	��[)��24'tڤ�t�&���Vp[1���J� @"��Ȇ2s%V!Z�L��6d|�����tP��AE����U����&X�!���3���-�C��S��iH��x�n�0.�#�fb��J�3ٹ����7|������:�̾����w�|���!�#��G��z���M��UI����qO�K�[W��'}�R����"c��b�e^qD�`c��C�ع��a�[2ӛ�f')�����XN�ȑ�g�TE4RT9�s�w�y-�+o���M&��؞Y�sTw%�?\���}x�w���|�]�(yO�ق�����8~H�B���`��/Ue0WQm�,a&}h��a�oA/˾@]�q
:&%��-��;�T
�ǂ�̍;���<,H_��h��v&ѕ���Ф��yA�S�CƳ@b��=�{*�;z)-��/��V0S�J��[���é]�0ꆮ�%�2�v�6O����C���.0ex�Xh�D���
���`F���r���|uX漁��|�	q���A|���R�|- W䖈��<�L����r<�������������r�Ԗ���¨w�D��b��{�a�S��A]vo:�X��ƟI9����˟�J��z"f^��_�;�'7w=��?Pڽ�:)�=2fg��.�r�!�c�2�i�s�3|s1U �8��g/&^�Ӫ�J��g����o=�"��w�)�C��h��)B�1=�������6����3�;6�5�Y��Ɇn��u��+�Gp��+S^fu`����Tt:�Y�%�)���q�U�
�LcBfh��,������C� ��Q�j���Lz�5�p����l���ϊ�A���l.�L�U��e+��5�Q�E}L,n�)��Kt�����5W����Z��>��u�j�σ$<d����II�L����=,��@��D\�DWQ�5�`~�0�U�H��f]�7���=��n,ψ�ir3����1�T����Q"7�Ő�O���W ���
H3����W�Y�������^����ضO)lr��<�tG�I'����O�9���5ٽ�L��J��;Hׄ�R��<���2�n�����2c��PrџIr��.�g�a ��o���L|���zw��B|��3�Q��F�p��RÃ��=_X}	��BR��?�uG���[�md�k�ȝ��ӰZ�fk5P��j�)Q�]O���<�N�*�`�	��1�N!��|�C%��	�b�X//�s��e�#�3�&oб�C��f���J9���x���-~�;b VWe��:鎪L;B���]�+R�x3�݉B�Q�I�+����FR&���� �M�u8=2_p^�?r]�g�7(��˹�/��u.�u�������z�j٣��mh�A@��5����4����E2eâ,@��Ngd��}s�k�Z���o1�5G�~-����4�)�}е*�ފ&�+Ꝟ�}�2]�%d���n�\?�����/��+��<C���O��d�7��٪�P�� �N	]]%���rY��ke��3�ҥ��E���ik��,�O�Q[�Z�P��c��.�YC����e�q�0�Ycx�CJJ�0��_ c�_�B��5�:��,��_�;�Ers؄��U����
��m�N�M:����W�=�hz��(>1���h�>?.�_�і�}P*�jԪg�&Q�p��P�v����l!O-;��(� _hbLǠ��h������T�v�x�ڊꐦ����CI�3|'���ݟ��m����?z%-W��)���Q�=�<jJ�h� Ԕu��L ��t	0��M����� ��� fZ�mh���˜���Fl[�O����)�뇾�����
�;���ow ���^Z�Q)#��1��-\��#��A��XD����s:�$��
�~/�y�Ϳ��S|�j�td�o*�bto�ʧTlb�4�IA�g���`�lC<1'ӎC�H��\�J���0���v(��n$�&��x�~!�I�D�+�Y��-�.X�p�B�'�+��_�ws�� �z�1�f�X��X�m$4:+g�/
�YZUC8�Ⲷ2�.$� �>�����cu�e�����A� k�]-��o@��y��XO�H-Ydk��xV�ِ�z����]�:@2�iz�����ܛGA�ֿZ3��rQ�M�^_�t,��K�sq~m��%������y�EDPl��$��'�q37;��v��a�z�&h�����5/ߔɹ�U��*D��J*	�\֤�ii�R�3��������~4��*��/�Iπ�r������Qf��h��+�pr�jWPQ�u��D�S����r�h��t�an����n�^	Q�ʹzX_�T<�Oƞ�: ��;�_R���4g�JNh�����HY8U(��8wx`���t95�B��\g!��]J��Y���$��-'c؃�4a�t�ڡZ7!�Sp.dEFg����}�h�Dm=��'ɤ�DH�w�Ef��Q�77��.�96|=C^Q��W�Is�<5��Ӡ��9h}b�*�UlEL���ɲ�*����0�B���m1n7=k�9����E�D��e��M	
w�%�Wn��/���:(��� /-���J�-��s+�A<uP0������r�5�#���:q�~h��nJ�6c�*vv���D�`y�t骗gi_H��[!������ڊ��GgS�O�٠T���_sz��ڠjES\���$���r}�|iH�m�+��P���_Q) 4��G�`H�5�M��R��uK��p`e�B�T��w��l�Sxf���R�a�*q�����١2���ϓuw����!"j��ED�_�)�����^�� �wMܿB�/�K̠�R�O���`�,�����7�^�CMV5��HV(VH¾��cc�=��[��X�Q^�����@�k1��Y��a��Lf��[��<G�'�z���	/�F��9:�Ck�X�� Q�w�<]>2��l�`����(��B���U���d3�}��7��
9�%L��aW��lP~��V��Y��?&�i��p8="�;ˑ`m._�\xw �z���Qcs���(��j���+�P�����Ց�H���>����^�Wǡ�x;%�e�Uǩ�OA�9\�V�C����*R߿/ݶ�(�x�)�DJSq�G-�6lm��"o"VR�gf0�'u�8(�����w�K��Y�?�T��"��sݥ�U<�Z�W7����?��#J�=7��T�G���v��Box�ub�K����.E�t�H���h���O*{�7Z��#1;�<"��-}߸�T�#'��,���4�h��B.�~r�֓^p�m����9(��iB١
ϔ��6�-�G�Y��T�b��o���պ�D�.P�1K��=H� tb��#}��F��G �b5�h�1�i!}ď�S:Si8�
���Q;��;�7�/F/����"mW�]V@��H���<(���I�Q\�P�,�i^���)C,E	ms�6�p-H&� �m��x�tֲ�˛)�Mw�Av���#�sv�*��z1�M��h=z�����	b�b��l4�ï�����g d=�b$ti��߮�4�uw�Gph~	�Ӧ�G%tj�d%�!���k`o�cIm��q�gr_@}x�hw�[r֔��d7;���-��ܹBs_������0 </���c�N"��A9��7V]	@&q�JvUg���� y��h2�E�9|Iᖾ���HUM�V�f}<�5�Vn;lN�9v,���zC�Y�*5�F�C�$�p�C� �Z�8�Jx�X1�T�L2�aU>f[}�s��������d�P��̚wt� 亳م�]-��; �'��X����:����� �Rn�MM��r��`�|�
0��Iג�{�q�L��6[�tU�.�7xIk8�"�vj�l�Ӄ�5.���n��k�M��ݹŜ� KH�W�C�u��7o����|JG�K�c���+�(��;(�\��.���n���a�G�>\%�H��;�D���6ӽ�ޡ�j+4"��{�Х��M�x׃٫�;Ћ]�
�*����*�u��j3�Y�/��!Yg�ui��b��I�	y�N ?J�뽯�;0Cy������z��[^�㗰�5�L��m85�j�2��ҵ�9.�mj�|��`r8�r��K�׍&�l�F ���)w�ݥ&�F��F��5ջ��Ǆ�P��^c�ōw���y�\��mZ�s��~	f���U�ߐlG���林��r�a��{=�n�����O���}5�������_Ņ�+e8���6+{�W��d��°u�9����6d��YH8Lˎ���m?�6op�g +^�?�V�6pG��<t |d�e0��/��N�ɞe/��*�e3�t��������Dr@���%����~�QT� �r�P�P��
�zu\��Vt�+�r��0Q�T�`��?Ǚ
���".��X�j��G.m��߆?V���[�IR;Q�w���u���4��dQ���n1���O� L�G��j�Z�^�dlD�r��0#L,���f,}@�h�a�sk���NQ�=�����~׈Ǥ梋S
��X�R/�v��Z�k��U�n�P��А̍���0�UKB��3��?����y)�M'�Υ�
o�Nm�݅������)?��s����n�\Bp;�ov!���F��'��@�&�yߚ�)�;���54W���J
X;���ɘ<�[�#��!�t�{kd>�-BOy�����O�!�����*;�Ƶ�A�!9+�=�͡UWL�f~" �%M�Ԗ��%W+[���YBl�76q����Y�IԎuH�lWW���Q�v�8�|Z���ߞ�{�$��9ȝ֙UB��┏���"sC�5�<����3j3>%IBj����o���L:5Wm������t5���#�.���3�E޻	uB¡�5� '+Y�9�v�&j�B�]�1��]F`|�t�?T)is���4�,#�f�NHC1] N5��?�B��To)m�z���֪o[��Q���C=r��/f���k�Ae�A� #�
;gWc�!�n��e�Ifx�3��Ctٓ��$��㗠��<���w=zl,mQ����C6�E��
R�|�"P�T�����'Y+k{8n��Sj��L8�އ+䢋{�v�$Jܮ���pQ����L�wt�j������pk�UZ�F������=łO�_k	uA�*���B�=Q��o4�2���憯&�]����ka<�j��А�kʽ&��"�w<�Hu=��U
n�iA�%�*�){'Az�\S�	��	ϝwVs�>��9כY�������{�7Rm���ZO2�s3|�@�� �z�"�z�~1��� A��I�L��%q�_SR�zp�99ƾ�}��g%Ǳ?�������sG���Zr����������@�rc�)$TF�ݯ�E[XA�E�����4�+�c��V��sfؔ�HZ�U�[_u���Ku�s/�+�SK��Ju��,�+0��C;-�b_�R[e���̮
tT���  =r8�s��\��Mn��%!gpgX�=��A$J�)N��rU̱���"#�J�aǄ5=�w�2IHc_�.V����+��y�x�X�r��G����䩮w7h�8$��xNπ�����<���{������S�x��o��uf	��oc�0OIG��Z��r��y%���X^-v���D�e��n`�l]���!o�� U���F���׷`9s���(�ߒ�F�Y=� !�v�>,w`E]�v��;;өgkȋ8>!�d�j=a3:��"�ft��~��M��J�e�$�Δ�O�LR�9r_��D�	��,M02,t)��#У����$�ƝlEC 
m�0��ޖ3	V"|/Z�Y�b��w��w����&X�Y�ّ��'u��pm�;�s}hm?��吜�����e�I�9�S�<��0R~c��U$�K���+~g�����3�4
�X���M�QM��	���z�ocDf��3�渹T�M!�}���lAQ�@@u��ҶX:��O�		��a�=����bb�a���j�)�s��<uT��od�k�SJ�7��O۫BWʽ���I�3F+��
�-Q �%%ɍ��(�l��"�y�ǩ�e1�B���(w.`m�׀�T!�pμރI�\��_��=��Z O�+T[����0\�V ��`2�B����'ԏ�?��{*��Џ�y-y0�s5hV�ͱ����/����0ˀ�	BnoA2�n�a(�U)$�*�Z�.Z�ʓqa@��,�b�*K��;�5t_a�|��S_�R�c�57���-�Ќ�׫J=��?�V���ܽ���DCv;�w�M4�]��?Х�4�+�s�sw�,�S�DZ��-(�MH%���{_j:��~��l�kϖ�C�a�薏��r�b;8��}4�Cֱ�w�)��a�����:̥�K�H���j`���M�=ܝ�S?f�ֳ]��!�
�Ɇ��w.CX?S~�9��)�Z�:�芟���lC�X��q'k���@H�Z��w�zb	�d�鈲;�v�s�I����>����YA&���U��3"'d��Q�>��$+�0��nC��/n���(fU25��p`�b�����y`g��ش�� Hy�o;��� �Š����ם�&��G���#Nd�3��=���J��׎6>�w�}�B	����@=���e�=�l��u����N�%$ͤ��H0��ǭ	�I������4�ܺ��=�xD��v����7S{�(�	dV�kZcq[������٭3�<�~��$e��!���km��:O,^���q�(:p�#�<h�~�{���tԱk9p��D,���Ye�<	I�LځD�ɝ�ٟ��J#��)}�u-`JˣA���
V�t���]���,�����έ��yt�?#a3� (�+V����8	M�Ri��{vǮ����1z��S�4q�cm4�aC5���p�_�#6��he\�d��$��Bn�1�T��H����rJ9j���3�b)�c�ØKF�+��渴��w)3#�]X���K
�>� ���
����Zݸ��hM��h]��a��(�����߀�5ek<��ٟx�-�3jE# {୉���O�ؐу7��B9�4~�����9)�~~�[��L��~��=���4(F�i�n�*v����������A~�9V��ٙ�w�@�ur1�bF��4�ĪK��~ckOJ_[^�H��k~&��R<�z#7����P�
���y��H�̠�bQQ�J�����󳏋|�:T?��m ��3��e��D���ͳAZE��r�ëΦ�_�>'�nS|��t�Gѐoۏ\��D�&)��R��J�s��`Zh�U˩5?��Al���Ӂ���S�fa)=���ڇ8$�o[?��x��� �u*dE�����m�u�F���5I0L?g[80�;H��&��tPt�!�&��%(����������Lo�܈AJ��KZe�r|��]�kw�����#m�i�ʺL�=ZO��p��2�ธ~<-�
 �	��M�!��Ӱ5(�?pQf�K�	3�"��/�b�6k�(�I��ȿı�A�wF�c�B���{Wd�h�V�5�;z�dk��i~��C<��)G��qm�3�96F!v,��jV>��}�#�>G�]
�9��g��������k�$8�!V�h�G�3j���wl��\��x<��Z5F�7X�����'�(!�l���'un�/C�4�{qx5�m�l*U�O�p��K=��E�C4%�8���^��������G��q1LVHgw��p�L�o���2���Pˌ�2L��!6��5_��K��?�;*��?�k��H��o������V��z�&�/zw��Fe�Dm�p?0-���-�h��`h�-p����'��;x,!L
�2�_�¹��4F�ʴ~1��"E��cP�ȣ)BBϦ�h��p��.m���۫��"1�D��i�nն���.{w����7�6i�'����Q$@Du��+��Kr
��� �	��c���E�9���D8�$�k<JT�6`a����"�4{�ꎦ!┐�-��jr,ru��В7`,3�"�0���8<���I�|��-�F?aFBT�`�V?a�t撮�4C{�|}�nJJ����F��Wh��g��S^P�Nd`VP�Q������59|<1��D�\���??ֻ2j0��xoi���^%�� 8[��ݪ\V�*���������I(ۨD��Ӳ-k�v���~���Kq1g?m*�}[��D.qT��#��଼/;3jX�c��
$�>a7��9�L��>�^����Ꚁ�W����^��R�.�����Z���e�l����	��r�]5�����Ĝ��D[$�k!�p��@�, ��Ʌ0�9��$O9�����I�W���q�#��ڴ�~�y7�=���1A�� �e�ՊnO�aj��4ib�����0���}�G�<��.�y�v��������r1!����tC�w(?�q�WO��]�E͘h-�?M���C*MB��{������z�h���QkG�p��-�v��
5��a/L$��m`~,m���v�]��	���dL�B�����d�U���fX����}�YG����a6	C�aLso���)����Y����od�[MJ��R#��-Ʋȏ@���,4*Ut�=���T�N��X����O�9���w!f��R��k��@��6R��k���6���,��3�
�w,ƞ��l�C�)�V�4��R�]8��)	!�MC5�����,�+o�&˺p������B�*=|���c�Lf3�}ypl+�!�Vw��lr�ctG?r(�I��q��b�jD 7������4��&������$�� �D&�Y3&c$��tA=�j@��A�ο���s�L2Zs�l�TU��B���vn�]c?Ԕ_���ij��8)f�"ӭb�G��y�>b���U�Vi(�/S�<���*	����e.�v�O�����*x�!��_H�x)2��E�V�QjN6�1H�Խ�f��#G�fC�/GN`�aݒV7!.���Ȅ2.��ml,�AC�!S��%f�m	��!�|���AhB��=y:��?eF�;a� ��O����Z�K��/�e?�3�� �c����s��o|RI0�j�B��b�9'�~�F.�2��]]t��ly��
Et.��u9��I��j�u��$��c�]lq��'��z��akpS���+��~�Ke��nhbN�Q����l�#��8����m$q�DC��A���J����N��6���Y�\��el�=�(�����e`�ףS'T�PF��ӗ�R�3Mf��	uF�m�T��#E�w2d�!ݍ�!���h��`7�8����C���j�n�~��_j{�����x�cЩ���r�>����!4Ү�~D8q$�����Kӹ�O��ފV���37��H-&`�4xɃ0�~����.ȉ%M"���S��,	&d��ػb�Iå��T1����V�-��k���a�<���٫�<a�C3����!N�)�]n��>�D��Q�9@/��	��ٯ�O=�-�:o�<z)_!��L� ��i��+UU����p^� ������O����3�W�Y��&�H�n�J���������r�(zI�z�C6���0��o���na����auƱC�c���.�tU�b�r�/�n�bS�~/�2�ї<]@K�z_;`���{�jQ�����V	�2�@���i����M*�z�����>F�=2�����O����Y�9��7�{~XOH�mG��	�N3�^��v���������S�}�cv�-��_�o��4���S�^J�7K��kh��'_����8n�7�ԋ|�ѽ5^TB����;�\lQ��Pyt:ʺ�G���U�(����e��<I���tc;V�r�c隖a�f�i�*?xɢ-')������*S;�}���Z'W�y��JN��7>s��y��n�O>h�J��`���h(�[m�>�cce�}NZ�m�g���^~��>��$ c���x�XE(z����La78��"c�~�e������=	I�y,��9��L�/����o�-�����+	�1��Ja���+z߱�k�!�!�`\�R7+��8��Ȳ�m&lriN b�#^m�}Z����;N��ʜ���! z �U�� ���V��s:��n%$��Y��+(j�}诲6��[|��k�(k�9���7�~F/D����ܔ���5�b�V��PK߬�"�`)��J0��'��gK5J�0�q}F�S ���ۇt������zB�b8����Β(�� j@K�EԿ�� ��qКg�#�E��^��M5�BOp��;$��;A���ȖO�m���\����L~�٪% �H�6�v=�� ~��f$����#y3��]�:_�]?٩�x�I�����X}/M�8J�(#�9�R����'xz,0"�{�G��8�3<���~�1x��qt��f�$H���lN��';U���9�ѷ'eI��>`%��>��DA	�����%�L��A>�W�_J���mǲ	��f̉M��a$� �}<D�Xb�ʑj�����4�>	$�� '�Q�XV"d�����1%�*0��oZZ�B�b�̓��g0�[pV*Fƚ��]���e�]�Ψ��t�]B���K�wv6n~z|��w�������vU��u����3�p�!$��f��Z>�T��� �8��ݙ��h���Z/$-�μ�sJK�����M�Dn��'��U��!�J�Kc+/�n�Rm+4q��Yx�Z�r�D�[x��H���f�O��4�����H�}�ln�����<�f������w�Qe&���#�_����QS���S��,*��XGX���b�e�Q�-���el���z����)f%�pc;���y"��&���eE��&V����u�5����Q��[�aG��Ƣf����)l�xa�Ӏ���)�����?p���j%��฾ׇ�SוVF�YY1U�� �K�M�qTy��Q��U-���vK@P=���F��ڵ9��U�/��L�S��.6kC�9i���$��wNld^Wݾ��w9�D�?�Ŀ�i�f:W8f�-�jYu/e�aʢ+��o#)|�������Q5��1���6��U7A���v�6$�geh���>�1�AϞ�n�g�}H*�	:��-I^�i���x��=��7�
��t�,M�����~��Ѱ�&��@~���L0���U3����ӁjõE�*���ꯅk��̯�ݱ	�3�]��\�+��=MH�����y�lceM��2B��X���{/"�z
��D;9�j+�J�c�5��"�<p�6�C�l�1`2~��Js"�S��c�e>�թ�p��2M���m����|�%��2�5�M�!�r Cn�jo3e�c� �>�c���o�:�C�"n��̭�x{�ADsW��n�Iť��!%a�j��Y��*kjMsT�������$@$ �3��X�ፚ�z��5�O
^�����@�[eN�[�~��H�������
O��uڗ�|U|�V6?;h�n���}o��e@]2�3V��f��Rv>�2rQ��L;���"�N׭sҞ@�������K�N3<V�m��*�pa��ug�k��,�����!��۲՝�����1�<�Ȭ���g�\D�]O�p�\D�eA�A�+%�ڻ#4o�]XA������rc<f��!��ϵ |���	���.=n�A?����j�u�j�NkT��5� 5�p��
��U�G������O�l�;ջ�wQ��&�rˁY{��aU,"QloU��n�(Z���!�S �$X���� <����"oӳ��?����ð%3� ��؞�<�i!(�յZR�9��1���Ӂ��[�g�K�]ԩmbR�yS}�ï��`��I���pŔ�ۇ���i5�M&4�g�n���	�Ծ!z5t����2qMA�f�F'K�l�4!|0��m(LC 8�(���������ͼ���[�\r`P*"?{rW��A�I�6�x�`���IN&�ǷOL8�q���ܞ[%�9m[ߡ���5�+$`+:�Y�|(�g�'EA8�ݔ^20���Q��$6.�O?��W]�}���a��{8�{���^��5��X_8��v�8�DΦ-��?�J�
��Sѷ��N&i���	����ANK��R8H����wh&[�MG���%6?���ն9+��m���@������˅�1�N�����ȽkfB~��VS��\�D/�X�s]�z\�D�$��u��Dj7��sUX~cd�R�w��X|y��n1��z��3�֣�)�3� �g�#3��:#I��ɮ#�f-�ȩ pJ�jߑ���m���0B�P^be�5��g�m��V,�T�EXz��]<jbT��ϴu��h`8W�,���p�
?��v���|�
�p��w��s"d9���'�ρx�j�o������pE��@Jg�6`#.	Y-?���7���{�Vy-���И��N���B�����lPl�B����MU�U��������8���B7ѠȰ�tn��Ң����o�/i`~RAp'8�fx"�A8�� �L@0+�PCr��H����k�	�#���nH �rޞS8o#Qm��bz�'�G���X�@n������/Dh���dkA�rݡ�AMU�<�'����'Z��Ӂmꟑu\���z����&�&������[���9�C�W��R��4�Y9�N����ޖ��-��E�xJ~D�X%�+�s�˥���
:J��	���x�0�S/�$x̰A0������kN�o�&�
,� \�WR��^� �R��ڈ�s�m�uM�KQP��>�����Qw�F���E�����W:������F3�mw]������Q8m�.1�L�M3mS���q��� ��|!�����}��?�����,��ϫw�J�y�/�f�M_�#�B>��O�kRi+с���ϷbG+�k�a��J�i���m���a��\��AAANL1�3�ur��Y��d6y�0��d�뙿oLj��R�6��IY	 �঳�H}�@~�c�E�/"�&P�F�%'�.�+�(q��}Z#(�;���Ǉ�-��J�`AXd	i3���S���M��_��RH|�&�E���ĤOMC38���	�m�LI���oZź�P��o�H1&0$��ڬ�rN#����݇��{x�q�lk�EB.Uꪒ��sB��S���I<yS%l3�8�����K����/�����U'��E����iS�`����5�W.�p��/ ?�EzG҅����Xm(o÷\8��W^���V?����lZ>�{C%+-Q��VgA�-l�@�F�s��<��,]؅`E��+�3q�jf���nh6��)8�]�eY��syS~A��$�����p����7,Tg��>u6����k�'T�+߿�v���x����27�X���tA��o�c Ip��ѥ����<�4of���x[�C�0�Qe��!� 0GȰ���\�bO���@��(��?E��|�׋�6}�/�h(�����in���{ �y�t��r���@Nd�
�ga7N-���;{Pgxˁ�������� B��Q�g>�ʹ�[�^$�r���Q5Ӷ����T�{?"ڽ��E�D��$��l�[}a�(Ƒ��i+�HJ-Ξ:QoN�9	��)�b���9m�[��u=i�o�ys�ى�Nk�u��І![q�E7y}�U��dY?�"� ���� ���En&�pAU�$��D���^J��/�7�
��/m}�f<t�Z�%uC�^�Q�H�#BD{vU⼖mP��5��"ɖ�E3�߄��V�X o(?Ǥ��+�F2	6�w�JT�
%/�LB�$Ɩwy��2���=o��<����E���@خ&�x��T��w>Ix\��P�������Fy����3���Օg�͸����� �b�4�z�"q��ܢne��'?&Z<�V��r����u Ř��*:��}��w'�2���;I5kd;+����
�����z߀�6��/����'�.G���{ ��g۳�B9K��l�;��y��q����w����6`r���E��2Q0�Q�'��JC;08D-�tJ<���&�����C��	hD*��fN���Z�˨�0�� ��f�mX[/���W��l��,	��~�^�A<I$f�����xYG�*����Jv^4r���/�^Ҳ'Cy�J��砜R��fQ՛xX��y"��xc�)V����J�|[@�K�<]&�@�wDJ�R��.[wsEܹ�楝��rn����j�V� k�s\��:y�'@���q5W�pϻ�!1U������9�w�M{�IV���i�݂M
u�}��v����f�zwA@���&C|P�������7)��qY�jg=6���XT����,��	v`?���v���1�VG�};��L	4�uD�N�K��H8���Q�R/9xN���jU���'d�oo�N(���"�+0m���o��+�}����O.����|7�h��YB��ǁڮ�`��h׍�M�b�KN�� t)�����.�JPbR�����E+N�y$O���FK��L^��>��@�0���52o<�Y�1VpD�zE�Đ!�kb-��	 p����!�	Y$S��)h��[s��m}Uc�y�3F�R���� J����[������Lif������z�,
~�t�O&��t��&�A�9�����֮�G��9�
����t��M5�Rڗ	����8�^��[j8�&fe櫳�"���AY�9���ft]L�~p�Ӡ|TK� ��u�n9�\h��ٱ4m��/�3Jd2i�&��?�����.k�r�P#W��)�2k�����4�/�Ql憊�7#D��X�Q~��J�n�f��m\��aus���YP"�TL����fSA!���w�
c��+���p�E��Bky\P2K��[$�4�Ƹj�j�=�ЍZO{M�/�-�H[z;����7�\�i�d0�0��N@�U��_�q"�ݽQ�
O#����P�,]!�+�7Po%_ؔ��v 3Z:�8�P�"PZ���yBzt�� 8U���*��qa�p�գue��E:�!siA��$awn��m�v��WݟG�L���ة��]��׀'�|_euҋ��׸6ڣ�!g��Q���IQ����-�I��� �q�('NB�7.�(&��@�$Z�5�T4`�+�fB����ס֯'W��~��(#s6�����am�8�$[aܖ���q�*eWLЯX���E󀒔��WF�cD+"�,[x�-٨��F������/�PCj��+�m��E���I�ph�A�J��~Uk#;]?�nf�SW�`"+���ךd��%��<�WO��C�[ɂ�Z�Oּ�IbI.�ntq�pn~��&2j^<xj���!��,NuC����>���������ooX��L+�
!�8�0���Hokǡ�����o`����'� �kO�d-���-n�&J�)t�'��v&R� ��m�����p^�n�=]�<S�^�~kF�L������8ŉ!u�)�0�v�O;�ں��4����#/H�<��R�)�s�����jg9:�oIֽa�کsM�#�f	POJ{�6��Sk�cl��ss��vųQq���o>O�X������l�TC_�Ϸ�e��'8�1� ��쉠0`�x��Z�C�U��Pǭ��E���0x�����;�Ӓ�y+K�"`�G�'���Ɖn�s���L��p1�x�D�)���#�h{%Y�������r�G����jy�+F؇��Y���A��	o��nvh���0�=qF%�y.~d��t�j�w��y��C��GMTPyԲ�y�M�F��'	WR�G��u�> L�5W�$2@�����"b�,"��N"	�6="�������K~�ڛ("���k����R�Pl�%?�����A�j�Bf�i�K�+v�̐�W#����=����_<~����o#�����߽9Ϩ� ������Z�6������H�t���M�9��,�?y"N��m��*.��Q���=�T�����Ls�.%$^�� rwz��
�Q좻�a��%ΨD�e���],l�Q���9������	-�lT�^î����-R*K���RD"�Ӫ,�"�$�S&�*i��)d��ш�O��<3�i���Yk^�m��R��A�����Uq�$�d���~��5?�V�/�rMENE1�^�+R�_ V�e����\����=~� H��~��-�w�O8=� ���
+���M5f�k"�E��o���o|';�B�]�@閔A,�}D�#U�}`��\�	$��f0��_B��[
jp䉮S6�5I�|�1ٴ9!��T.�s�8�M��UNt�)�_=�6��Fs�랱cr{��k�\D*�o1��@'��>�~��3��Ύ�O�>��j�Jƛ[&��#d��E�󺑲n4�<
�&�⾟~+ 
&��4V�/v�N�}�dT�I��WWj�,���O/·Y�;�/=�+�dB~-� J�ZO�/�VWz
OrH�<�/J���M��v��u�P�!�?g��Ǭ��M�O��������Z�-�ޕ6``>��{ck���~�<���ȡ�Rj�F�cOa!0|]��}>-A�*���4
�f~�D�<��^��!�Lu'��K�p͎g�s���Ɖ$}�L��VD�ƥ[�Co�����#z *�i�׉b�ntSBu7*�p���Fj'I�I��&ݦY!J�D����ֱ���5�S� I�'�Q��o��ѧ_{J���,b2;0˱��k[߄�&�f�̄�?�zk�J���0��R�d��r�U�����}.tG�<$������ЂHi]����8�/�� �#P��9v.��	תm��� ��p��m��X�8�5v�$7��]�c�֝�D~�%Hr
�\Y/�B혈�w���I��PH��q����P+�W>�.�  �R�r���Oʩ؁5�Y,�!�r�#��l�'�:xa��y{$_=�Q�*2a'���C�ܑ��?E��j�LһV�cǋɚ�NMI�H��5�5�	0ÙU}���Jn��%���%��5'=�@��䣃�k[��KF��\�v#�����A�:�k�oؤ�6����0Y��b����ۇ��H<��C ��i;O�Ja����?3Zy43�H�&��F�Wx.��ߥ�YrVsz2[�Z2�
�|�F9pw�l���څR��ڞ<c��Cq��kjz�F����|��c�̻ ��� �*�J���\nA7꒯+�`�����հd�S�0����+`�$g��ߑ��{�I��ݫd<��s��x!L��Q���<��ԝ�>�r0O��B/���]#na�����T�ǖ�y	y��`��0��>	G�L�	�[��i5�� �,��%d/���Vp;�i�q�'}�"��N��Owg��+uɭ�����(RS�o_�V�yCԄʥ;����Ԑ���� j<&�t�����J��n��3G���:iAGV*�ђI ���ֈn+���Һ�Z<�h��O�1u��I+y8|ܤ��䣤F�p�A]�SGb ����bP��O�!��
���	����6^_eeq�?8{�K�
 �n�':��ŷ��dy�Y�����~�c}\����e$���k�>J̊��w�u��0�pٺX`V-t��W��P+��d�ruC�z�x��ߌh��~_z�D �L��,�OM�%ϯ��3������L�Fp	�&�����<����3uDHC�����|a<)� �%e�M*.��-=>!��n��7��54�V��V�Í��A%\&I*����_g����!�w|�d�� �2��H���q��������|a�?2,����2s��ʦ!L��P��k"�p_��
2��>���e�V�v�؄g��s
˘�qڙ����Eq(�8�WRW�af8ql���t�Q6�!��^�2��c�����7�������S��f�A�ul4Wk�Y�O���!��p����ZֈՔ�JV�,��B(��
N��+36��j@�.BJ�"ԝA���V�2�e�)�*���LW�=�uj��1�vCz�(�������G����|���;IcLK	�4�����Ћn��jЊ����{\��'YZb�05�Y;������#���� q ���/�fD'����o��(�O����}:���
��Z-1&
�s$�UW�sk�tn�j��/�0�Cf�u�`?ss�S�)���O���Np�J5S��ӽ>ģ�����T����d���*�.�Ppd!��#n.<,E���;��C`D�4m�Cq�6[��6~�$147�U�X*��'��TB�aB�{��K�Ҡg��2g@�1׼�J2�$c2v{���Z�)���8C>{bo�ZLС��ɊN/Ή�)�o�Uj�l��C8P�vȸWČ&�Y?F�����G�ySU�NS�g�f �Yx���SjL�?�d���GQ����2����9�i�{:����9�E�;u�΀{%�L��C��Q\��#ɯ{�*�;84��)2.wK1r�F�����K��{��d�*�2-�f���D���+�Wv�	l�>{�����8�~�9��W�X�� ש��C	9���+�0�j�Ə�>c��]ׂ쀤�v�
*U*�{����+����#�J����O�&��
@i4,&G�?e��惵;>9�3"�g�:�������1mt)���Eůs�<qg\ak][�^���@kç���~M-���{��G�o@����w�v�!�;x���&WBK���{ɴ#U�sw?�E���l5[p�hE�����
A���)d2�W!�?��Ȼ����r��W���x���oⲗ�"x]V����ә��J�X-�,^�=LS�.��we�v�Q$a�7hT�4_�+˦n$Ӡ���d����LVx7�I&zEfBD�Q�l�o$F2�E7�J>E��tT�)4$��FL���v�ټ��=�&$'�w�u�S���6g{�F��X�f�{��'�wU��=�RR���qLr�y�OV�U](t��{�\�[�Ξutmq�㧱�9,�+w��5��AO�Y�
�9B������'1� ��p��5*��X?�QX.O�lP�B53[ >Q�t^hq����ON�M.�_���W���`�<���3;r������8��2��mg�jn~l��-�������%�� !{�	1�>��͇�E	�x�a���>6Gr�gPH7�����:/��W������,�a����0�6�\Zp)�tdG܋�h9Z�;�p��Ŷe@�܅�p��7�G.ۇg��rDz����+R;|�)4E%�iˑ���R�d�׎K� ;���~h�|�m�!�cw�Q�J=4���,ЖM��Z+u׶~�!���XU��.ּ	.�q�i�x�K#L����?V�^qz�>����vU�w�q���̤�e&1#�3� ��!��3�uq��ݯ����eE��#�X]�wh"0��:\�t�������,O`���kL���p
�3��F��(mO��A-;�^�e�S��%M�D0�h���'�%��
�ⶳx�X �v�Ep�EN�����,tc �x��W����>@G�ʯ���6nz!�r��)�*2<=�ے�O���^��`;j�������\D�]��_*Yhp���l&�^F�Y��F�,H!����_x��'��$Lڐ�z�n>�^}��I�ʂ.��B�p�����)�v]����N���	��xt?��u�m"#�샳FW/�OW1�����uHK��$߫���}�T��!-�\aD��'��Ͻ�������m���9��\���2�k"ʜ��ܱ�;����$�Í����I>
��6c�a�E8��i�V�)�����FvW�Yo!����Q����o�;��ҍ�z������v��ߓ�'��+ |��q��0�$�)�����(�?Ȅט�F�_���9���bN5�[��T-��7x�E���Z��*%����%N�JڭS�ts?��>�4e��\�+�(M�:��6�e�bv��9E-�����GxȰ���w�\����8�̸����@�O��(�WRP��{��ڝ�To�uc��`�)Vu�������e�EE�
"V��U�Y����~����z�HxyQ�Ͷk7����ub�]
�����[��!�-���cK(�'�~I)1v)�
0� ��75?s��;x5<m�#�����o�U��������F�[
��v�U�Iy�i�\/Qj>���zñ���s:*+q�♏w"�Zf�-�={�Z;b<as��s_TϷ�����?�b3��KM��o���Χjs䫱x���5���Vp_�M*�y �_��3+��ҳ4]�<o[�%I*!�D���(�j��$�O�-��(��S�R�\E �?1�!,9����'D`�[���[��YU�doo[�Q ��҄[���qz�^%�Dke���M2�ّ#V�����N��%(�)��H�H�fndB}�n�K���b�Re�����6NXq,������I����돂�
�TZ&1��?"��B�S�������d��0�����υə����8��Z�-�;��D�yo?�3xT��@��Q�\����Hl�ۆe���w�"�g��^r��nX�ݻ�|f�ŷ��z�;�#���ˤjF�PLFo<h5�����KV���s�2p��iy��z:�UF=���j#��Y���
���QJ3C�̈�jVY���;���貉�	C���y����GH�-��n����T?q����쁇�>��h��sN��K�x��	�DR�:I�y����Z��tk�Z���D�qA��:5.��\�=|?*l�Q�6�PUqV�; vAaήF����]Vγ��_DUl�n;&�GX�8��R���[Y(g�Җ���f�h��@$�����f6�fG��A���&��,�GX�ݲ��@�ogq-�J�-Cy˧��(���~��fn�L���P����T�I�q�j[Ȧ�n�n�;�X��{8�wRD��aL��c�0�Ѡ�.��(]��S�9�m��'�jxj�Lc�$N���?G�/e+��7b	��jye[ͬ��el?>����W�mA�s�l���������H�� #8����@Uq	l����K:�+p��]i���DEI��3���+�n^���T,}r�G�
?��oŗ��E6b8]�Zbh�j8�8nqWe��y�F�I�*-<����hT��q@5��)�/%#Õ�V
�a� ���KS��iC	e���!=Ѩ��������.P�d�=��̶�C˸�œbv�`~�Х b�����f.0��u�R鬝B���H������a���:
�����)�W��w0{��zhѷƾY��ә"����+��Z�=l�.�K[�%'TLD��.�j&����@-�<^�������[t��߶������S��E���^��.(�)��a|$O;4�T��Y�O�%�'&(<Eo#S�&�Pn⼸�E|��|���~^=��T�هL6*��Klo�ڄ�T�ܚ���rߵ%�IwҰ���8�ZA���h:�O�ȁ�j�bpV���J:U8<���4��B�3f0V�	��h��,�U���Fx��K�'q����w����%f�Y2�<⎊���Gy�3w/����ի�5d��z6S�w�r�u=A�����F�)M�s�K+8)��:=Q��	�[\��:Q&9I�V[.7%*	���%�Q�>U��!�����7�-+��$�������������9G3���"C�J�,1Ĳ�d���v�&|���1�E'2:��������vՔf�;]g�X�S[.�Fu�Bp�Y��'8��u��"��Vc�P��Ȩd�)���|�`�qt��ԣ�A�S:0��';BV悿��*�a����Մu�PԴ��0��IS;�"`�����rZ�F��T��'�R��N!a�σ���h:/�pYŇ�u�5�:�jw�Հ���Y�˩���4�|��OD�0 � ;&�ɀ(�{/�]���o��;3����E6������6��j��j�Tpq�V�ϕ����7�gsNm%�\j��a��l�wQ��PD�3�l��=)K� 
ބ�x����e�)�6��	�0JG�V_�?��𐙈��"����L�'������e(8#5��A����RȆ��U]�z�Q�P@�6�-�����`gn�>�d7��@$�(�ոL76�5�œ�c�rj�\,���.!W�-�F嗺ϊ+�ׯko����t�-a2��ؘ�(�7T�­@���5��g��
VÅ�ΑB����M�*���7��KE�'8ch����Oڃ�	��n]I��^$oO�&�
`��X�FL��(��ڲ4�1Y�sSWM�^Ҡ����%s��jyk���'m�aJ��9:�"�@���G�����*�����Ɗ��i�q"��J_��`x8[�ytSK����R���/��B(�0W�`H���7R؜��%��_���`fL��S��,��%�{t�Q��NuL�M|J0'�[2lX翷61 �� ���}K֥�X7� 硐�7��
4o���)h���]cH��u����1}�l*�dh�uSY��9��	mb�y��� ��&�ż�)rhm���_z!?��b�WB�Q9�vZ�� ��=?-�z��J����_���`�(N`[��^�.b�؋��0��K��4?����4M��U�����6#��zj�
��d����;EI�絹��5�0gI{S��G�)���9�Q�vS�z��cR�Q��G�O��%掮�$"�4]>}�ީBg��"���x�=ʚ�d?K%�ԓ��/<f�%��\  ����.47C���6L�=C7�n�,�$������aC7�iV�4���j/��YѰT��ѱ���w��3����GoiŌ��V�^�dsd7C߉!K��\�ǝY�-Z}�?�!����֙Y�ʭ����d�����;*�M�7>S�P��%B�8��Y��Og%�$bZ�AO��t���l-�s�1w, �d���dDt�~�U���Z��#W^�($fU�w����ʯ�,92�?���I�e�7���x�~1?/���C���`�����{LYpBJ�'&۴kj�?A(�n/��B�SkQ�J���Z��wag/F���.����O����W�t/�Y��R�<X�2hn��x �̗9��Iv�`xP�@2�T_��؟���*b�_G�~o��67&T���m���ɗ�]��!�7��y%JJPKP*���І�F����q�x-�
~�V	�4����'CVm��U�w� y�f��a⻍Hu��M?o]����C���V?i�#��T��h+��.�7[lW�;����\����򊴇�]����o}Ÿ�(=|�e��<t��]{��b?���f��8H�[��)�	z唒&�;��~S��;��+��V�h��G�1� ��h����������`*�d0ЏUI⾓��
���Ǵ""�?�!E�}�� R�&�8��BT�vgI<y�UT�p��h�#�o�1q~`N�~���U~�}٪ q�i��
A㶁�c-��6Aی��iLt`{E�5kEj�G���7�H��u-A�������X��i%!Fj�Đ���Y���H�_����Ҭw:'|wk�5F��=�Z%��1��4<����ܬ��dm�a����\��1Y�(D��9����ٜ�9�kX�����l��e����%�ZLlL��xM� �?��6M~f�/ڃp=QJ��C�b�`�o�ɋ�*�Z��}c����p�kj�p�<X]V�5�4%\G2;*��Y�tk���;9pJǮuX)��K���9�� K�c�	�;��q=��q5�/�V���y6���۟2Y�X����}7�a����~b�C��͛x��!�#��x�xX���Λ�����	���W+���G*?F2�|oS�xxUl���㱚r�A+�i�G�-6L�U�MC}_Fk��������
�KL]�@�O��1�����[fv�]3t¬��?��M�K��QF/��}�� �,��j��|l}S.>���?��V������9��������0�ڭ��-�8���s��K?}"�L�d8asFb'�/r�%�A����w��H�u�Ӧ��G!�3���W]��-���{��(���Y�2m������������l�,�,��֤���K�X����8Pu�eȃe� ~j&8���V�T�R��J87d#�~����	���n�H��	�����ߑ`|�c�]��n*���0g9�ci��3�z�ټ�Q��'�;y�)�t�5[3(|T,�)ښ)D�߫N����<��{�nnb��Tf69_���,,^�E�����ޥ%�/Ԍ.a��7n��]�`O���Ǚ����|��M�<S�<��ƈo&�i�0����1@�KX�ɯ��E�s���1���gt�\=�+�7%q����
�#ǭ����ꝯS:���{��t@�8���
�7*$\�߉��K�$���>k��A[/� ̏������K�G�|�R9�G����H��P�9�$J���W�$��.��c
�Y�pų͹�-�Y����>u�Up�'ֺ2���R��RL N޷��ꐉn'����Ĉ���
�� �~���+-�<.h,�>"Op<��#ȡ�7ux� �$#Q�X��a�0D��8SvL ���{r��U��y�(Ug��[cmI� n�ut}��7�X#���O1�������T%f�x|�աȉޚ�{VA�c������q��!�H�<����j5/��@��L��x"�X��y�E�ޣ _l��.\*F����HY$Ő�/��J����P��2�bo-�����>��q���K�6S_�Kh:��X��N|c\��T=a0��|�o����ݐ�`;{�=X���}!'\N���io�X��v(���Ia>-%�u1�E������=�P�#9
=��%�k�#�i�g�o��9}��-T�F҅G��zd���[�6 �θ���<0JB��)A�J�j��tC��*b|$��iy���i��E0�qD�<��'?o���,��#¥O9H&�~R��|]!W��|g�����K�L50��D�����E���æ�Cؔ�K�gKM����yz�b�V)P��t�A��A�4�C+Y ��}n�t�lbߡ�8��~���:
��)-=l�h��ÎCкd�>�V���,�,���E�=Y����{��x�Ti�~�Z���	��K���������.ɞ'q�?�y*'z�U��-j �nE�^��L*7S��ˢp9ۿ��� e�"M;p��)~���L(7�E� �07ȞJ7��?������cGz�-}b1�~g�۶�l�_��qa|
0�;$#7��A���֮���*K�p�JX� ���˛�)h��8��@(�����ۭ[�g�-�.de ֍,�C��=���j=ŷi����|8Q�K���
B�L��I�Vh�����f"�9�^Ce��ſ��������p�i���W��W�
EL�R8�&���h��
��Xl�Q��~?�����t�F-:�z���@�@.z]/�E�߀:�� +�Ƃי�/wF��b�:4�v�Ƕ?���w�K�v�r���]&U������	��W=����U[;��$�Ad�~=����5B���>�٭�B�kxMa}�h��=�c�r��usߎ���,�<LU�}��J|{q3��v������.���kѪ�o�:ʾ!��g<��P��|� L*R6� O����ެ�����q�0Z��Ʀ�ڪ�&w�+����Q0�Vd�.)_�G�	9d3�PX�pۤ�$�`���M��a�W���ֳ7Us�gL�Jm���	W�a �������t��D���s0��Y7`S{m��"�%�k�uNB�u~����q��B�]���R1Y��9��� "erz	dF�)2W�7H���p{��#��@=%`Ow�g�qX�Z��f*�(R��&w,V������Cl�ʽ���e�hz X���)i�:ۂ��DG]=i�nJ7]���ㅊg\gZc�
]�Es%���g�<C8/���u�Ҕ=��,�~�1sJj8/�P��:O�TU�J!�W���w�|�x��K��� ����#�Ʈ��������O�f7m��(}Ǵ�`n5f!�'��&��qǆ������HZGp�1��̐�i$�'�e�^�ʡ���R����,ږ1�KX��5S^��Nyε�Ҍ}r�X���k�+�Ђ�0(��L�����ڰ^�O����(��2���V��m��7_�k�g�)���06²��'�����`X�޻��	�Mqf^ܝ�ঊ�x:�[�-��S��S��Dy��u��
���y�l1Y�z$(���17)�V򄝃��'=����<��./)�LT���]�v��h�hB�O_ǂ8�<��e`!��X�;�:`b�6x����|\�p&�Rۺ	�=б�G���;]&������(:!�E���qӪ����]!�����$p����&��3AΰG�FUIv"�����#�$��E3�� ��i,c�xa�m�yo�7c!SH�"Eڜ�0m��T�������[yP��<X�J��V��S���D���΅�[_����͡:&/"ͥ�����#5U�1]�z�S��7�3����J�PLٴ���Y�r6��wG=+���t��%c?N=D#-R�!=/�7�-�Z/�2Z��/T�,�!IYP��F�8�L��zb���6�V`�G�����$w�;��_�����f��w�&�����ꞕ(.8E�C�ϲ�*������z[DP(��GcJ��8�Z� L�K�L��ڛui���<	�F�>
���pw{z�6�S��ا�u����b�y�K�k:��5�a޳���>ڻCLW+�
�����zu�LR��?W@6;��F��r��}0Z��Q C��?�я��iSwE~Nl��� @�/W᜕���f���LeoFH��ɯ�!�8�	㬡��*K>y�+�)�|���i�;��� r��.����Hq&,3�a��>�wN|��`��n��O{v���=��5���|��u��
�L�uC��~����RHP@V��i��E��Y�*=�HԽ	.�H⣎�Q������)���;���klGӊx�5j���8;�h���b<�7���Z'���YA�S=�{����	�y�yF�ܒ�/�metS�q�CS�E~�y_�H��C���1)@C�� ����L�o�q�.��FI :4_i����Zz,j���vl�UXyUb�=Q�;CF��{��P]o���`�nǷX�I��������$Kx��]��҃}Q��b~
yK�*WHw��Jh�&�=� S��'�� &W�ϿLR�"�z���O{��	�+��&1�m�E'�mQ�/>�6�E�^y pU��$r��v["�a K�U�V���8P &ɑJ��҈w���~��{dɃ�q��P��ų䵛�$�IM��$��[]�?@������B9�E��Zb�T^yUt��W��0F<}+ۛ|�O����`��|�O$QhO)r�1�ݺ�30�m�M���?�(XO[E�-n}��uw�#=6Hx�@�Th��0����ύ@�Urrѯ����~g�@�W���
G_2GU��b�OE����l���T���̞�ժ�U�����vM���8�2�;?�q��9o�ˁ���̗�ó�J}��<�,�	e�Ϲ�ֿ���i����	��؄F�����2v��<�c^P-�^��&x�Ȣʹm �d���{�d3vLb��Yy���9� �l&D���6���������p�{݂�t��Z���brvĹf�cR6/�h���2��I �/-K���f $���}�{����|���&KTљ�∷�i1X���#�B^��=w�|2=5��J�̆s��qcW���V�W����	8�V��������+�Ѥ�`V�	�05,_���A�ui�s�F�	��Ѕ�*�I�sʣ���4���۷9M�����>�|�ξ�5�����MOX���Qϩo��#�1�hI�Z�����*�P���T��<bNĖx�]Q��u��S�$[ ,ddJif�@�sr �"�*���0ܐ<�a=��a��E��Q�m�=�������:�4=��/���5��R�E�m�A�o��ߑ�ӕ�X�����l������n�	A�)��D��=�aiD��3���yvz/�64�ޘ�1�So!<�)T	t�'/Cޭ��a(�b���` �E���\$�[�
��~6ZF��-X"��;?˸�5�I�1��D�j'�74T瀪�t�Q~����^Q��S\{��JL![(g�ϧ��m�P�f�HЍ��{,�ҐOS��49ݭ�>�6ѐÔ��dk��N��G�՚.7K���K.�hԛ�Aן1x�k���&�@�?�c'{}�;Y�j߸G����_y�������;ż��HP�s����ě_�w+d�rtȫ��m�p�]F�SV$��j���-�D�4��4.�$��{�8S$!]4^#7޺ŰG�XT�7B���/nř�����9���|�;����YLB0��^.ۺܸY�����K����x���t��gU.�
b,sx�<@��3��}U#��O�B��t0M�L�Y_F2%K�U�[MQ9ϳB�Ba.�v� _p/Q_<�j�Uxa�89��\5���ՓAJ���Q_�z}P������wh�~@鱋,bKEJ�����S��!�s���Q\�ū�p�`��j-ӿfG�6�{<�����Sܑ�ʩ^�nU�f�6�-��2�0���s�y�(��e\���&�渰6��£L��l%xd޹��˕lX��\M�e4u��.Y���Z�PT�pT��G��A5:Hh4|�)~���������,�����H�toè}�ut��,_)�!+��ﳎn��]��-$C��;R�M@VI�e�%��x����S淗��X?�H�3N)�退=4���I�7k�)V��v���-�=��|�Q$zX�$�3��}���y���e��\�qfN�xCކ����%��$�����_[�$9���X�)ړ�jӵ��MwsZ�&� $�;���:�����鴬tXeUJ*���T����B����5�)�v�Qݹ�O6{�.U��fp�J Gm��ov�q��l��W����L؄5OQ�hW�	(m�),/@�L1�so�hmࠛ�d��)��ec��I�b�"�q�zn	��&.�%֬�<��Yv&ES0�p};m̊������Հ�>U���o�@�mٍ�C}�����;)�-�*,-�0s��+cAh��=�9*<y�b&E���V�H[:oZ�VGj)5�c,�f�Ι��Ui�s�v�O)4�h��z��AAܕw��k��0���ޡO2>Ҝ�`hZ�/&t)������w9dl{�����3�vd�������>�O>����k��k(�l�+<W�;v1�S!%�	+�?z��� N����#�����BS��!�����`[���+b���ŭ���u��X��uI+��>B ����_���6H�v�:��vp�#�1l�M��Z!��1#���B�<�Ļ%r��Nj֞�mЅFl ���02b@�+dHp��ʰ��r�=�
l}en�[F��.T��J�Q9�F̞�]@���9�P�
�gW�C�9��*	I�Ζ�~����N�S�D���r�W@g)Nѡ�Sz�����	�w|��0�mmǁ^YF�C]�p��'ܵ���[.�+MǼ3�9�H��1��9�׺?)8�03=�Q�zsrs��mL�,�W2Ċ�,YP}W%j� }1�u3<�܈�#����:��D���W�{�=��)�y�����~A���) ���=��;WeԵ�#�W� �p������WZ��d�/Ħ|����s�}d�L`�:�Uw��VCS�C>6T��U���ԸF�td�~\9oO�M������N�l��M���w�:w��'-?7.-E_m����քbh��w,�k'ۨ���<�i��d*tr[��c����H�0Kͦ�r��+dS��l��:Q�����~�Ofu.��+�cU!#Bj;\)�C\���m����{(C[�JRzJ�՞�_��'ի��TvJ>"L�~�L�l�D�ϝ(�nz☐t[�ټ��GE"q�Z%3����'��ʻm��w�f���Br�gv���B2���ih�ྥY�����F٘H�gӏ�;�8��`P�\��\�km��3]x�)c%&N���vʒkGd�ۯ�Q[�@|r������b�tZnﳴF����1[ά}g�g�mn|
��^q-�Rj���a�j���A� �'Ig{�F҅+�*~v��hUt����R�Ӫ!:�vAk����4�KC�)j��ɀ�l��;\V��<�kd�l��ƅY�63��s���y��}���-4�u��؈V�T���R;��R�9���Z�`qY����[|�f���h$o;��I�.�d���S��`vUK�M�t���XjT;�a��N��
�R��J� m�K �c~Җ�
K� x�9�:����!�`�fpQy���C8��C�РN6�0|BR1��T(�@��(f����XV+P|Wg3��T�#����/��)?q�̄��ۛ$�j֜'c˶����~/m&n|�
E���~aH&��P�����F�"�s���t�w��q���#W����cȮ$��۳��JS��n�~*����d�%�eSB���jh�:��t����Y��e����/׆��r�ʬR�f�o������nh�Z<����Ic�6��}�73^�y�~�+qĄ}��q0K������S���{
�� ��EQ��)9�CuD�r�x�t���.����:s�.4_jR�O�o���K�ѣ�Y��:��jb^�ۢ�r S�$�J���k:*U�\�_�QpM�:#���"��8(v5�H2�/��ȍc�B@��+9�u�	|Ry�v0� M?b�˅Πf�YOa�b団TA�>?���&����׍��I� M���e��}����<(�.s�
��E��?Z	a!c2zڹPZ_��%D�r����?�d�+�.��ͻ[Q7�A�S1ӥz�3�aJkBT�t7P~�a�� ��7�l�����Zm����1��f��Ve͕h�>9��d�^�J)����}�ف�x^���_��ji`��TwW��O�h���R��Ix/�ϣ=7�nogb���x8��՛𱞫�P
32�fXX�f8���˼c/-���D\����W.?g�tBD�Tp.���S6����hJ�V��';��,6�zc��}�2*��{��ؘ��|%[�������b�e�&ə{@{|;=;�\���0N��B��)�dR*��}Z�1|Ykr�3B.; �,S.���'˃~7��j�'�?}���'�s#՝^5�*�:�ׂ�����Z"3��M�<0�z�Dn���ނǭ�Bz�,���c9����Q3m�)����A~@V�`����cU�*����&y,q���Iu����_��m�
�ڛ��I��ӛ:��jU�sg�3
b26	ؿ����M�CU,��jco�U(N��Kqp�0ߞP�������|��f;32����-����o�Gў�J�).7+4�� �¿~�{hy�vCg�d(���s��F��qfŢJD�n�h�FK��l�:�i�]�U~��a�EaX�Iku�� %�Ek�, �����H[��ny���_�\R�|vS�d���HD������+�#����@���nR��.�(��DW��|��fh��u��Т��@x��'Oѽ�ܤ�ty�������X�o^*I�.�/�|Ǭ,2_�)��~�s+� tOt�]p�_4l��̈z4&�U��}L�w�w�t(��{�+�{(kd�/V�˱gAہ�č�Ll4�b�{٢G��������F��	��N��E_���
h�KPuP#�	 ��U�6u�ǝ|qk�x֟ �-�o!T��I��#������tM�J��[1A0�c'�:�E@w($�rS���\(���	f���"n\���i9�ڍ��6�u� -�6D$��UF���n<	4��Cٱ��h�}�2�$Y�ӏ��|�̻PX�D�!״M"�*�(�"�)���o:�����lQ3~��2�'*â�����p��܋�_9�5�q���Q�1E�X���FZ��v�5F��#�<iҟڱuꭢE`��*���`����H����;���pGQu�V�G�I���R�����4�ac��L1��c�|��
w�E�	�6E�<��	x��:����4�	�X��#V��PТ��Y!2�A�$�=��`r`R$z~^�m�#�8�}���K̷�gc A;�s���e�z������XK6�Q6x'[��ݯC�!��7�=���KN�c� ������U]$t���;?��R�!��$a�EZK��c8���J�I^�oPEۺ����X�޷9�_枛s������*�KNV�P m>���n7Ol�����)�\��MGI<,�L���x�f3�M،��� W8:��ٻ��*�窣�_�:�`nR$6s�-���t��^�K�&-��!����e��"��V�ܖx�+��Ou�t>��o�w,�8����	??z��9�p���r��.�]?c�O���B$�pmn77 ��$��Iԅv����x�����}{���|	#n��, �;����	��n��/�~P5��^1���R�<����
s-�]x�P��8%����;7z!/vSGAS�J�
Q���7�{��w�g�-�J��_e�?bق2�)Z�DK�f7�h�������
�J�(4��~^Н���+��=�낊]�D�f��g ��5���Hh.��i8~G#��_%mE���eM˕�¤�MՠO�2a�t(��Yt�I��ӣ�v)�-����4Q��>y��#���l+Y��4�8-��s�Ok/�� A�fxG�R��Mr��R  ݅�Q̲�~E��{���n���Z&L�{�gQN��tz\=<����m%�"��	���?=Auy2J�;T+�	i<�0�`��Ҹ8�ȁ����B����U>%AE��p�!��9r{��͑��&�lѷȧ���e0ϸ6XU��8�A]���A���p��^-���x��Dv9�֣�* ��ע��ž�.��`_�,~<�]H�"8��g)��dDE&�c�[�ݱ�L��a�󑨗,�:e�j��� �ܖ�6m �������#7�� !K)�*�nf���#�63�oJ��4��fk�]�Fs����� #�=�k88�7�����d��+V6C㲩C1����1;�z����	��q�������éj��9��52��w7"*�L�H;+=F��#x�5=����^c�i]E�-�&@��"hv�������w���W�T:\|͖�;��f�:{��
ݖX���%m�3����n�z�8_YX�}��:p�m$_��=m*����W��<�Zo4u�d��<H���1����}}_��� 3����|�$&+H	�o;��ǳ��?'�g�l:��?�o�%Q;VOST������/��.~�����R��19��'��p�.D�q�����y�Py� 6S�>�;�ד�����H_@��.�u��8���{F$��-��St��Ee�Ǿ�I+K�(?���m�FFP+�-���b5Fy �I���қB^Z?T��y�p{��d��Q{�s��$�i3-ڽR�ͼ#�Ag੩7	wk����^��5C?"�6�ku��@��d&�_)� 2����D9��?xI�5���L��B	 �'�8�ID�7���i]�m��y�Sy�ٽ�p��ڠS��y�!�=����na���*���\�Zqe�O�$~�]�+ �~�u&Q+�z���kP�#��d�_o��G�Ȯxg����.{�����}1�윔+2o���RP����-4�m4lc�&AA��97�#����4�J�ko���2JS�"{�������7(�k��Wv�슄m����:�9\�*K�
+�lZb��2�ļ����lb���M�����~&TĂ��G:��~3��y'U"�;"Ҡ�*����xF��,4����f�_c�ЕCQ7Hq�+H뚈/~�2W���Q�%�`Xp�!�-��Um���ƚj�#�ٖɉ�:m�#昳�y�
�q�X� ���_��đ�"|6���;~cBR�/�	�R%�jS�V_�nt����GL%����ȃ4p����{*�lG� ������fK����D\+��@e��f�-q�����;���v��e�Ó��0z���$