��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f���9�rQ �rb�?��K��]��a��qY@?�9߄�g�� �`d;Y����d��g��{6����	�o�C�)���������l�kOK,�d��VMMC��&=�1za�)G�xF��'Ŭ�;X�8�k�M(�$~_	���q#~|Fr���W��zO�I\�@���j�N#	X����X]��7`��q�0$O�*�f������oy܀����A�%&�����k�i�_�
�w��N�Y���Ǌ�2�h� ��:a����aJ��/���Kv@vh ��*a|�MK#p� ��u�P�lDb��v
�!����At�Il'�AA'r���e_����\.>�j �`�m:�f���Y���/�S���ʚ:y�)K:���ڸEp��Di��
<�1�9<p�f��O��)h%1����]��h�y��@3�dk����b_��DN
�t#u��ǲC39��Æ�xj@=�%�6�	�1̀����ϩ�xD��K̜����O��`J^ó��wD��X������8H/@�^�������)��Ss9*��ɩ�+�eZ�=��}�K�$�t��z-����6���ZF����S��ir�I/��I��f���FUڗ����]C���4�i�[�v��y���4���R���L��
0�\H��F�F�;��n3��~���Y��-݅	����7�Wt��ұ�����3�-��ڣ02�uu����ѝ�GL�[YC�޾!��Eg���rq�Uς�Q~[:��"\%>�׽��]���0O��@$��A�tH���]o�Xޞ�~ ���<p�M�P=C�4�
�ڸN�%E7��om��kH�)ڏ���=u]QD9����5n4���� t�V목C��$��O&��1��!~�8��Yܸ�l?�.\��Ě�J~+�;�<�rc�/��P�,D�\���觲m��2wo�_�kT!L�o����xo�<ff&�'��1��?��^'p(]�gx-ycA�j�YtnӦ�6��):'���HڒO�7� ���/�v����v�͢e�����º���W�q��1/�_Y�V.�7�OK���!��}l>�c�W��R��HD��'�e�W�}��U�c�q�-#�����"�?��ȭ)�p��T���o"�o#���v�Vn���q�+ǶK�c�F\]h�ԁ��g&Q����xd�!k����*�X�_�*3Z�㑫��3�P!H���J�!�:Q� �\i�Pņ� �|�O���"&�D��1�~����l	Fؿ���*��!3Y�0A1��ҒJ�g�ىR��q��1E��tm	���t-;��^��S��8�f�o)���;	�q$��\�e��.�Zj�9�9��#�����S�m�>�0�m$�",�h+7p]�^�ީ(�<�o�&�u��sG�=���]K�\�;gma���8��TW�jT�~ޓ��?��zR�tP���觸0�x(�"/q�+��4��v;�S���ܧ7���D����J��`R�K��}Ĳ��� ��T%��FI�։S�%zp���L�%w�<Hߌ�v����qJ.�W�L,��	�~(yf�����<DUdbE��hV|�Dq���Ø�K�s���pTsQ�A�zg�JzCԯ�̅/��J��N>���|�ʿ����&�ڶ��]L�RW�*E++���� ڦ���菍a���&?b���U}^��9GR�"��%0a9�m���=�CԪ�0� X����m��9{ R%B�����I�5:)�!t<N�Ju�x�/�ڤ�$�n�@Z�s~�k�^"LVe(po�c�yy��kXW�ʋc}��+<M��S�=43<~��m>Ƒ��\���6Sq���]��r�)w�=�h�'Ho����,�P������i��F޼�)Ae �h�'1ڰ�hܾTa�H��X	.��3�Z�'.���15jx#-G�E/��8up��I ��ysYOo���"Z�9�����4�bm\r��o�g�$����ߴ`q��@4X,��[#�ޮ�?��Z�`u�NlI���ր[|ay���C,�p�Ɣ�=}��G�2Y
����d�YE��xC��#`�}"CT��Фb��|�@�2Ĭ��f�~M�ڋz\�Dv���t�κsϵ*ƶ� �!��]�����I�Z�q�P�D����{:��,��g�cE�.!T/;p�%J8����*�_��7j��1�z R1骟�8��g�AM�2������\݄�&�6ֶi	?� Z��Ŕ~�$�ig��Z��� �u$���v�EJ����j?��|l9 G-��`q1v$�v9��麯}�5������ChK���@�vAp�2A�F��x�P1��EC����~�Pm2���/X7yYy`K��-�#�P���}S��q�ۻ�%Ȼ�Mzu�����HfmP^��'K�[���ݤ	.
��DX�0�k��	����<U��Z8$����MCd�s^������!�����|�wM�HδCf��x�C�+4��hNZ���l�I�����%D,_�Ku<�$�R}#�3��˶F p���;���#�1�;����~xᾳ(˄���3��i��'��w�nP��*<��a�6?�g�3�����v�qÃ�S�4a����2�����v)����BʏiC���y#�p������%��7s�9���G���˓`�%��N�,����W]�d��Y�*K���帤Nm��ۖ��ג�S]�d4��`��q�S�\VӖX��։v��N�s�"�Iڢ�[�&��v���?�.<�I�3�2@`�eĺKT�%'f�k(Y�V��W@��#���Md�v��j��Ra����I��i�	e�& �Xf���\H-�5?c�����c����2��#|�J�v��i�M0[��g����s�/�28k���"S��@���c�n/��c�����׳�d�#)�����t�͠2}iZ�∆�(1CB�D��WͲ�en���o��_N��ƅ
fd"�Z��U[}n�o�Ot*Sw@���G%���p�!&{S�j�,�5��ק