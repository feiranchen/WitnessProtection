��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K��mo�G�
����c�LI$��#��%n*�D������2
�<_&A=/ĩ�vT`%�2�@�Ӯ���bR�)��(.C�>�M_؍2,��EA+(����H_(�Jn:2��f�1êPb5��[B��������ʠ}iƭ�Z�k̤p�<�7b��F���� �[���U+7�3��V�����3�j�[I��:"T�;�Sn]w[����ILG|z����
�L�g>���$�z?B����9��F�sLp�2B�ເ'��>���;ME�������8tS�j���p�5v�}so&���@��x�ٴ��@�*
�x���<j���DL�^핳���p�I���� �ә�8a�Mr�'���.�aK\�����Gz��+�Hm޶��D~�XH���_L��i;rV�-���#c��Φ���75TB��52eZ�F"�/�(wG���.��=�!�h�S���Z
���c�ܒx�'���ڞ����������W?��+]��mՕl�>��2��	{ΤfH��g�!��XQ�'�&\�ت� ��kS(�O�+��U����Ӏ��
$��5k��V�&<e����%�'��q�%5lo&��f��5R��ӹ_uPJV�4Y�j��bdׅ�
r�~�Щk�ZG���_�2"zQ�!5ޜ�f)�x�~V��T�2f��oiM6�՝G7�|/R'BKTǲ?]l�ҩ��Ԩ��� Ϛ��n���oqur:9=Z��P���_�Ju�� l���⬸	sz�� PQ_	��!�I�r�9[d-��78�g���zP%7�Fk�L��k�#=��bU�K �r�R'z~-.��,<R��͊�J�JШ"w�|t��8��?�O8\D��?��=�F�;����.+T�������պO7�+!�:x�귖�9v{��"���F��Dyi]}�"͆1�kC�⹆i���\k�c���b�Ʌ��m�>I�	+�gU�?JO�m�F�R�urC��Ə�A)�&ù��z���`�����NS��h�}ݸ$������c�C�˘�Z9��H�V�'ss��NC̼�e�FƱ��,��nC?��HJ�@ٷ�/Ó(L�� ,�Wt�~���(�2���)!M
�]!�m��ThR����ڦ(���t�7B���/4�<���9�a�����ɟ����M^h��cLN�u!ߕc�B������}�r�AI�NIM�+r�n�V􉼸d5��L����%���x�s���C�Q�C�.�f/G�5�֥N$;�L�T��K�7��s荑(�����+S&���F�^2qѶd t�w���σ�DT��2�����Ȏ2H��뢎o´Cx՞z�~��w
���WE���g4F0��o�q��Q�>Q��<�#�9�嶄���
��f�~�(��a��NI�˫zq�����d��y��{-9y�F x>E���4��4W�|���wc��4`��8ĭ"$���Ǧ�H����|���.:@|��X����ӕ��6l���(������%s;I��uUnl������C� Uz���"����y+����^^��14_�$���q���Mg��"�N^gj�~{	ˌ8��ݬC�yB��T3�Ϫd��6Z`��)L��Ssw��-�A�i�s���+N;��9��%=޻[܉��=�����Os<4��&TC|�A8��ɦd�4�� �Z��"��C�Q����j�ky9Q����`J|u8��o�Yt�A�(e�L�-�i?C¸T�2Qt�KW\��-Rk�od��z9�K12U�<�����H��W�[\E�r�5m�ٺߋR��:��� c�v����T:O|�3E	dل?;I����C��mK-���:��*� U�E+�k<�~9d%vSޑ-��6��H F��,��54�=��얞XG������_�F�.���tj
޾A
�u�R��~s�$B��9�b�l,� �_՝�|P��6���,1�l�ύ��L����7i$�\��/�����wA�@�1��o_�0O4\EoJ�~%1��|s���=���X�^����8V��F�
�?pR-�F?Rtv�f���I�aˮ�Ӏ�ݘ�4��7���S���A�����{���2��x��YH<?�3��n+�W��fF1�?���SgW�(��N	zW�r,Q���9Y�5��f����0���=]�Qr�:��Q=`�/e:"ET�0��r*��B�3i!8������7ܮ�zCPa�iA"9�� *��3a��0�&G�`"	���hY`U+5�%G[m��Dl�D0oI����阮͇���*���<�&�JM���.���r�u#�i5'�>0y�����{i�N)��	��FLS�!����[*;<׹�U�&��	b1����|���U���,��"J�XW[���SW�=�?���X��r?w�i�@ă�;F�Jn��eH��C|Z��p>�<�f�%~���߈k����Hw(����'��_w�Wh5�5=�GޥvD`'���&П�"R�?������順�}�B=�B�ٷ�BD"Ȗ��ȷ*-�*�8�����UO�k��hB�t���� 	�F脷����^>��]��Pݣk8Y/{�����#8ViQ�Rc@��{��_`O�i����ǹ�_��Z[pE>8�]ԳIɒ��	\>Š �=k�kS{8t��BZq��rn2�w���yD�$���c�����!SP�66�&��	-4�_�{�� XƢ�r� =�+�$��ЂS�`*����%��+��6�*��]Kv�
=�ֲ�G�.���j���-�_%5�]�0/<���t�.�2�?�ť��6F�u���R.^�s�\�`u(Y��6>v�U3���;�j�~'�p�[�u�ڝҵ�+}��u�u�c�����$����3WLI�B6�w����>��N�HC%7�,~�a��2k��寜h �9)��0�_�����0��q���!��'�3Eǹ�1�bb`wt����!��2 	dV�����Pb�ڡ�!�p�������y�}���ce�^zF�ֹ�5��1-��� Ӳ����(�L���K�=zW���l'?$��˲�,����*�ʳ��f��~��L�te�9_41�$`b�5yMs$��_V�/ɟ�a�>1�,I�3[��JT�973Z�Kj���~e������۽���{�bA��%/2>�J�v���z�]�6�CM3ˮ�>����%�����U�r¹������a���h��j�j[����+r 9*(�+.�^�E3�X�?��a��Q��.09�t�Y���?����5���ᓝƬ.�]f�z=�ص�QQ��OY
��7�y$,U�z*ʴG>��