��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��-��5&I 6��mb7*l�����	��ҭ`K�J!BZ��dn�*4���'�#���Q������k Qk�i}C��
�K�W9��}S�4.7���dR����q����0/��kK$SJ:9�v��P�rqQ�(�97�O�������ҽ��!�V����^���'y!�M�#�;��b�'3i���V��;^��e7��P�
M����ZM�ޥ
�E(�~��EML��n4(��GKU��Č����>�f. ���Tl��CI��xT��vY̪원ذ*�ۺc��{�ϕuP����-:�(<�+з��`ӏ*���4O�PB)�W�}'�J��j�+��+����Q����/ ��H@p� �j!��e���p+2�:���� ��I���2<�g��u�X����N�že=>8�kkN�k�3��S�)���q���^�mR�</9%?�Y�k0aV'IZ���&��5u�U��>��1��<�t?��Q�x�nƗ,���I6�[�"��X��v7j�N�Q�d��l�Dq̝[b���<S��H:q��4v��\��OjI�����ʇ/�h��"t�D�n�8>+$�-���aRf�*�{��K�<>x��~ӟɨ?���A��.�E�;@��(c1`��M{�i���P�
�S�Yw]l���^}:��C�$�����O��s���.�77s�4�A$�K"I͸r�J��z�K[��e�1�+��/m��3�r���=UV��6�i+�J{�A�P'��E`t��y{]�W+�#�1�J[H5Ĉ���e�J�
�X���Mm�9rV�9xT�Z0 �}�Z�F���e���f�j��#������A�9�a�BEq7�Jsg1ƀ��	��G2�P� s�@�$����12����m�<^�����UWLo��Ct�ꚟk�b�k�u��S�R-�#�Z]�QfB!'f��i���H��<xJ�H�o)��Q��U,.��X(P0��1~8RC���i^%�xk��Z�c�Z}L[�)����qd'�3i*��i�N�M�O�0�F��p�@��QE���DC��_f�o�|vh�.�IT������cKSF�v踠4;����s�1�� �������+�ߎ:K���o�+ �=��;��Y�:뚄���}�W�3��,��=���pd��N�xG�B���
t���-iw� ��abòɫS����'n�Q�;YuV%b����Vo�r"G�yç�2џM�X8�.U�+�&#S�&s�)�e��w��{/v
�in�c<�@�R���Z�Xڰ����楂 �T@�h�fn�-��g��)�E'<�^p��h*�y}z1��DL��� 9S�|�&����ֹ�8:����&�fn
"�/��Ac����7�o � �{��K~�\/���cX��*������$w��v<�k�8:��Q���n���G �w��鱁����&��j�fV{b�m��� qT嘽�To��0D���H�z�ō1x@}필�*�\��='`X�K/��'m�~1)�umnx�[������F�j�}"��֊�#��Bx�J�\����#��ʣ8� #�c���ffQ]�
���������-rO�$qN
���qh���G�߀�W�u��6�?�oyKt�����K���I�n`�$ܨ$o*�:˾$�45CB�F�6��n��������Q�q��x�t�_���2�x�͌��a,O*C+ @���*LS����<{}���;�<UѬC�k�����W�]�k6}�fS ���Ȍ�0�x���L�4���ɺ�	�N,`��*$=RA�� �`��^$���1������Do�q��h�������1�F��g�?,<x�P��N����1SK��?O���� �H��[�FGC��������$��z��U�D�Xe��!��&ΌV��oA��ae�ek���8�̐s$�U�K����gF�eh���}�~�=��Z�)3sh��{�F���M���-~-|�1Qf� ��p:\Ԑ�￤���O���T�	�_�w�4KU#���ee��p�R�.��U�\��r�<���H��۳���:�E?Մuz��4Ӂ�w�������̑K���1��Վ�D�+=3�TLP,��z��������;�	�)W���~�Գ	�R�HAB4�ThxQ��i��T��91��'�D�AѥU(�5������l�΂^�e��3��/�]�H;�Q U�r�ғ(��0�Z�+�'e����п�0@P��;Zy�Y�l�wen0}#S�C,��O�9>=U��|�S�{���?��x9�Wr\�M�Z�}�k͢�{���%F���qx�Ӈj2"��m��xա�佋Z�r�<�C~�,F�ߛr�؁ҟ6� $� ���2��T�D.J嬯��0?��VyZ75�,2�S�J����)8xz�|��	at�+'�	eV����Ǒ ��k8&Ǭ�98�1���J�o6�X��*ko��:	�0Hz��S�2n����+�8��[8�Hf&���r	�2��<�����}�X^L]��ȍ�r ��1��<�HZ!naepa���m�`�˃�=�����6
ˍ1�� �?{f)�_����ln�weD�tC����ԛ���m�O�w}�>��8�k_���1�H79>����;�8 �Qh��p}=Sd�c"t�n��J�1���'�����B<�s�"!v���/�۽m����|U=�n���|<L�{ǜ����_8������?s:��0WBu's�f8�85��������~W5�3!�U�&��8ga�Q>T��cmX45����|M��%�?Hx���d���;�x�����]��g	��N~?�2�����s��I��M0W7����o��Z9�|& ��uߔ��G	=#ILf�ı^S���UZ�-�mp�_u!��)Kr�	�`�|:����a:A����݋��)�@��^�ḧ́�iJ������s��nW����o�[u��/��N<Ԥ+�d��Zz���G:�h��fg:~�*��9����1ٓ� ��&R�3���]�mY��t��U�o붷@<��19��2cg�lш��rP���p\���͒逺Y�n�Q�U�_n�GȚ�1�X��wZ,��1��3_Co��^;Z5��{~lG1p�~�8���/��|�Ѳ���;>����rjl�~�@�8*P�Xrt-?x���������O;�>���m
�T�-�W�I��d�l@���dt�z�����"R�c�뽹VE$�5�]rM,����m<��`<�lxId���5����N�Ũ�qw�Vs<W�DM.5�Ȍ��*h�:q��d@��b�J%+��|�Q���-�ۂDV%H�$�����'G��Di���4I�$�"o�36�4-����o�.t��5��8������\L�	4��E������/
oȘ��Ignz��w�h���@R��'�����h�Ё�z:$��KT;38�tg�@޵��'<͕��t����V�!m]|��9� y���c��|�*+ɫ0 L'������b �c�*C�h�S�B�t���ys~l����~���O��_�e��,}�Q��z�{�W�Jd�0hHj]�*�����9�N�JZ���ot\_q���!��F��t��M�P/�Ռo�B���A�k��Zv^��.����[���Qp���t�ͥ���&'���|�Ј�+j	~�.${�1;"XV�j�\ک�N��*d���B��c�r׋�6����ó��*�'mА�#lz|�ʿ������U��=�r�B �MO �^�@X����v3�y�lc�w��N]�l�a*��"�b��(�RL�x�����U��0`#�zF�|;~����}(^�u*����O�SV�g�M��7�I�6���^�o1OK	(}�^�d'���;�V�o0��lì�x9H�M��'g!���F����o�IG9PϷm���%�ZGTc�X�<�1s��\�U	�,@wz�08���d�EDN`�8q`y�X�4~��F�(��u���@��܃��4ϖ�.ۆ�CCxj=P��;�#!]Yi{h	��rX�ɛh���tZ�q�,Na�4s`���96JG��eټ���ƙZ�� ��qX
��[ض�K:pZ���:����%�qb�����K�y���K��W�럸��ik�������