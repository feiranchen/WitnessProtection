��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,����}\G�Tγ����s�rO���x���	���2T�o>�N}��i��Z���ko�W�� ���,ZE����M�a�T��a�Ӭ(� *۵X���fT�С|ja� �2rɷ�}n߳p���ˍ �����Xae X�y�L�I��3֓?�.�R��+ ��H1�u���:�2��9����n�8KRIau�,6�
�U�v��,���wԿws��.�|C:RU��B��8(��<�w�^_�@��S��y6H�>���U���c�p�_|�k��9|1:a�88�">x�O$��5G�Z�� �4J�����b6����&.fe�����g��\�@�-�w�جnv�0��h39��4�h�6�?S���}����a�HH�x���%y6��hZ>I>p�(v����%�#�VXQ;֐�K�^ٽ/���V��#��`×�kt�v�
o���K$a�"���uWW��A��"R����-�1��\�ڰ����k�׿f�dS>H�,�I��W�J �6��6H`L�J :��l�ڦj _v7��9Fz5m�s��jR���T��H�4[ȫL���c>�7� ٛ�˒��}%�ė��2����k��ꏑ`K�<.�90�Mf��q�Q�G��f�`O݅T~�&1e���O�=v��O��s
<]eB���� JH�zL���U�ealN��ߔ �(�%�pM 	�2���av����|��)�c'�˟F�A�O $F~ӧtn��*JM����FO�6*ʮ@�i,�ٔ�|H�kY;�n�.h��� L;6,�?߹I,����f
�D,�
݀�_��DX�����r�ߢ3�H�������*=h�_���7���t��4�����A�:	��l��u�p�,�¼���p�����kR��:HE5��?td�@�Ǣ�r��2����;�
��8+V:)��n��SKC!��j�:�FO�KK�K��	!QPV��o�����7�Z%!��y:��9v�����<�~�@�,c��_��EW&u�*{�H��pW��88�h����K�X�!w�#��k^/"% �ښ�En��w��ovKy}��'D��ʭ�6�. ��XLB�G�)_.��)d%������&4�Ǚq�?�V?��s`B%+�_�9��嫙$ϹCG)��}�a�j�fek-x|���v�m�_�j��ȏv��1$.U36Sƃ���bL�m��[":��\U���h�E�Tڴ9k��"w=@��=�����O�[+C��N�4� \<|���C�;�A�29h_�"$[����o��
�?��~��X� �kV�Q�V�r�PZFՇ�"�?�,�;��fR�N�޳rK�����J<�8q_���]�=X��"��w�<,���u^�K8�D�Un���o�W���0���mt5�nE��uQS�>���ev�N gP8���Xim�4�r����+�#�	C�= �������ߕ�p�@rj�"���ZB��