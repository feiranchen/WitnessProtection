��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�/R�ؙ��a8E?	[��C��|_EM!���MP��� �R.Cw�j-1�,?���Mׄ��E��T��� IZ$\��h��I�d���cL�mG }������3���@T�G*C��'���"t�a�3kM�����p�s��7�Q�0�[0�yS-*e��۞�`4�,u H��{�k�p	O-O���I\��vC&�] �oV�T"f��.�=�-ԙ�v��vd��__)��#� !�z~A�]�=��ւC?��!�*K$�G�kFԪ# `����ȡ�T�����}���Ys�-�|p+�^���SPb����4m�]���$g�O��z�}����.�F��O	���d�C8㿗(Uz���6#��}}s������t σc}��J㇔x��#�kh�u�g- �ƺ��w4Q���p��e��:�@�-^_�W�z<�6p�P�2<_��Q l�yP!`ۖ4ॺn܊'�(��-xl�qH�"X!�r2v}#�v� A�*[�t�T�N=(X[�E�37 ��c�?9���*)/V%"��))�j͓�i�=��M��D�@�h����n����!�/������I������-��\�Ōw-t[����>�E:ؔ1*��7��ҹ*����S�6�̲�D�U��]�|>��9n�p�ycf�|�FB�H0���Qc��@J�{��j�r�~�$�Ԗ�z�D= E�;�gMj{�!T)�5xR7m��Y����>]��`\��m�W��^�'^���*'Ű���)Q�|G
�8�v��}�*�7NY�S
������ ��^�*I{(uٙWN��o�c�rV�Ef X�x������`Yd��D={xk��.Cm�dl����!�	��&��~�F�hE.�����n��"�)���=���[T��ݐ]�Y(�򦭈1���I,�|�"�?h�P4C�_2�E�1���+�ϵ���^R:f@�j��$0��^��x���N-nQ�Hw+�Qh�؞B�U�\�'�>1I�4���_������o��kR}��4mM ��nm0�q8�y�_�6�#N�6��o�L ���0�r���%��Qq����[�E#�9t�?�'���8�¦O󽾐E�˧>��w�a����4>��j��Z���B�*�s_1�dCY��Mm%3w�sQ��>��!�Ԥ�V�v�Y(0 
����wKp��2���R�f�XV�(�͕�1� �I;>�8*:� xf��`p��&d��	�c8g�M�S\��@׬g�`/sӳl�UM<ڕ�װ@�&r��m�@!�|���)	p���:8�2�I)Ȍ�.L�����`);T.�$�'J<��,� ��;_���7َ�5|$2�,p{�y�]�D��
[�����R21�o�����rUd��YN�S�[�������.����{jr��\�=`�K��s1�JGǮ~䙂@y��\V��+{���l��6X0�����J���V��|�}��պ�<�[�{�e1VM��"U����rEs̃hD�����/oO��Q�c�Ͷ��o�Ӛ&q����NG)����`�ӷ������_>�ʅ?����Q9�^S�^.�u]"V#��S�gߘa�O��ϧ=s��f]K��y�(���A~��:��mxRU�U�kg�#q̎#n�;u<����1ak���Ʋd����߹�����]�	���5Тc��
�}��>�Х��m̨MR���	-T��@�"x����ς>'�f�'�<�\u�H*쪏C��$�]�upS����Kk�3�^x(��U���睔*���;9X�6�MB!%�X,�f�+hǬ@��;�:��n'��T��9~�'��[E��ǪA\M|�'�]*`�uM�3�c�e�l���瀕����� ���l�W@��K��m�4�ݏN:k�0��u�}
����$�P�M`��S�È���b�wY=�p�(�e�S�_+O�s��29��LSw��ʽʅ��j�V�~����m��b=ˊ�:$�T4��{�`h�8�R���T�GFC��[�����fT��\���<��z���]�����C��O�l3mwĪs���J��!HQ:x,�)�7�JP��_gs|����Iå#7	u�V6�஺6��>�U$������p�p����g�~H�(Q-��3�G����%D ��t){?���[s����Ⲅ�ū�D�L��p]EB�9��^�G���.99��vg����(�@Cl��S����v�i`hbʴ@�l�Kƺ'3f�L`�:�\0`JÕ|iy2�ۜ���4<�@�4}��1r�r�?=��\d�'��rW����O��� |�Qm��㢃,�<��NBSь�o�� n���� �,�6��Z5����"���`2	�E���K`��b�ށV�r-�K��?.��>��8���-�i�mX�B>V�!�Xzr7����f�_'��j�]&j�RA��%����ie�S�V.D��*l��%̡)F����s(�%��R�a�E~��l���.0��&p�0��S�/Z%�3�d3�{Q�sR���J��NV��O��2/���8b2cjFG�mn1ph�bsV�~��Ge_B:�d�5�g�N���ܯ���F�QΦ�P��hz���ʫx^�Îg���u]���w�ąk��a� ��D.Z�ǿO�p��Z�a(j��bS��0�0�ǰa�jǮ�A�!�P�¹���o׍��8N���z���eE�r �D�;���V6�U拊���p��iEO������9���uhŻ���ȫT%7��ϜӪ��Ơ�eev��1a�!��·Qw�Z>8I�����Y����	c�v�{����|]��y55KSV�\��9m�^?�{�@&w���L�tF@�u���ht��G>��Ɉ����u�k��Ȗ����ޫ3X�.��w����w�H�EV�;�z�:t��}��܅��t�>0�����(/�W���}�̌�Ji̸����7��٘�<�������������,L���x��cX�"�`95�$F���6_�ң\�u���8{s�8NS�E����u�T�)3�H���P�������\�&��l��shkDh3 ��hec�	{7��'���>4��'z��p�:c[/��h����0��yn�fw�I��AW� j=�	����.I�*<X��/ٚǒ#�i�����l����9WYa͉�����Ll5��5�#^ym.�l�'4S,c3%�������t�B@�����Re��6>>#��}$5b����c��U��e��`��b�m�|�ơ�I���WyN���&�7 ���Q����
���e�8t�<�m8#=���QP�� $Y� a����a�UP���;�t5=:~�Z$&}Ķ�;�V�hZ
�f�Dq�n�ڮC�q��E����,ȁx�uC����f���)v���˘c!$"�ܿm���Na�ϐ�%�������}��P�2XQ�%��$)����H}N߱e�������ݡ������2+��ޢ3a�����D�g`�iCN�$��4Ʋd0I����[H�-и�;kS�MS.�\:%���1r�%W`����a����gl��8�$�Hq�<N'K�FC��R�.��k'ߣ2��a^ԟ^�3I�6����ƹE4�#�R���)�b��"�NU|�PhU��1�})��	^0&p�In���j5}�`ޗ��	cf����eY�vN}<��y���k@��b�~G6r�n�4#����+����鴴���z������p��1��2����VF�"�Pq��H�Y{m��f���'�oH(99�;v ~:��H�7�4ts�[�Z�T��-s��@�|�h�Ø��d��b��Q �Dy�p�����p٬��w!#��]]4U�>B��ۤ��q�`H�t��v���W��|S��<��I߇W�<���/ d������I�B������ч(�[�]���2�O��.QZ�o|~�����5!M�fX_�����C�ބ΅qD����]�|�M�TA+d4
��F����Y8��o�^��.DuڴIz��
�V6��C�J�X�i�VX���QS<�����]�H!�-��u�0��o��k'Η3S��b[��JԬ�ӷ�ڡk��|&�@�f�x��4	2��
�;c�ƭe��x���������]�|�ġ�Z��&�;;r�!1�00�������3�\���`���T�UXD�g.��
���d�3ɂ�����0\�s�n���w�c8鞺�T�8�G"�Px��H-�!�L�?8� ׭��:w�vS���.jx����R0���ܒII�� ��8�hZ���V��..Ҽ�Zc�e����@�X���C��٭5������k�W������B�ɢ������IY ��ۚ�\��(����"��2���&w�/��	��J5�D�� P�zZ��,����YL!XepW�'Y�%U��V�ۺ�e1ԓ�8��v���{z��F�R�<k�����������ռ�����	
�~�_u��������<	�MI�����������sy!�n`�V%�����D�1�i!�#u�ͼ*X�/+k2����2����0���O�4Ï��{:�3J��n���g�@���;�U~�Άq�X�M��O�d�m��Gc�7䈆�nsK*F�Zt䈫ݮ�\RaB��
�,XFM��km��@��톀��W�j�������S�O�n�z��~�i����W:�g{W�r�v�>��b yء̓� -y��~��W�'�Zt�C�ڸ�\��(��"���)�D�ډ3���R�\X+&�����a_�	\xe�[A0B ���ujd�JtXYX��s�8��.�l�1�%�hH����xZ�������W�H�F�.��#u�'=�
�X�D��z⢝�ɽXm��C��q9�6?�s;>�Uw��(k�����o�W��w8�$�T�#Sg`���Բ�#�q<:S�}ڶa1w�=\Z��$�̪Jv�4�A�[�1;�G��BT�k1�Y���������cʔ}�H#S��:�
Bgg؎&�@�8@"}����b����^�0�c��t�����E{M��z]@�S𷿛����E�2���p."#�2�z�iFA\���0�p�&y;N�a�I�_`tE�ۖ����D:9}s�M@�T* �*3�&��T��N]��n8��7�~y�Ϲ����&��d*t��G�;zc"0�Β������������w�	���.�F󢪒M����b[�nC�M�N�v<���u;h����>�܅o��V��yKㅯD="-9?�����l�Ot���&�>�}$)�J���/����'=YC�>&m�Ίd/g~*k�n2�"ޯ�֭Usc&C�����ʤ��?=�*���A4M���R�?�����uh:���ѩGJԟ���x�"v7ALk��E `�Z����Ժ�����*4J�~"�"]�>V��l�0�T�}�g58��^2���a��B?��WT;�aa�n�v}���u\ݘ����{�s�za>���;>��+6]�<`�������+�Bً�X��Uq����e0]&����LT�>Z�q�S-�B�����B5�nj� A;���g��ڠ�^FE������9WsY��;��5�8���i�	��/�#�C��(FI=]2�h�b�=�gҭ"�P$�mP��Y�E���j[�DO?�t�&ٞ���
~�Y��6
�U�:�֢�\���U�H'��P�K��ă橪�8E��AZ��;Ւ��/�h5�"����=��.���!?��--8�Y��/�4V�
�2� ��Lv�X�a��t_�������v��L��R ��qւp�I�
�ƶ������Q�IspT�RR@P�aV
wt�~�~��)9M"�u�QE�:�U�ځ����|0����I?`���2ۈ"��դ�x�%��׍��T�ƣV\�)�+��2ki��| ~S��Z%<g-hbu�b*��X��3����!Q�Jx8�'g{�I�z�̫n��x�Mb�$�%�f:9���Oc����_ہ M5��^t���p �8
p��y<��Yt�����ED�`�8	�Q�%) ��ͅgO �(~�=X�%cr�\}{�]�q2r��I7]����9V�f,ZkR_�w��Y����la��^�`�Y ���O�V޼%x#2��4�����4�k��ZΦ�j3������#��q�=����B�@�w�o���!$ѽ"�At@bf_��x��`H�L_�X��p�aNl�Ij
|�0,'�Y/�LfK���e�_K"�^��}p�&��a�Z=o�~�AM��r�EG�2rSߵ�.wy�0��>2�}�f��p��i%7s���Ɵ�8۴[}v��\@�?�M>%.eL�V���l��xf�F�f��'E�6-RDiL� ǖH�m�>�FB�ww0~[�]� ���j�O9*���1��n^��#�MC^$6�l�� �ly����: X%����K|¶����I-��R��I���m	���O5�^N^+���7�+ �l�e�C] ���с��>�_8D�8����<[���Cx�x"ac�^� ޽�.	�\���Έ3c+�����1/J�ɯ�j5��ೇu*�#3I5���_u;�m�I$d�e��}W�w��G���S�::\�b�y�&���_b��G�2��|�ߓT#�����a�"oP��t��"Q-{�����6(�U�N&���[E��%����+R�@��Q�f�H	[�9<z?/<E��Y�h��{ߦ��tE�4g�1N�3��.�0�($����J^ԯ`2��O��c��7��'�Mo G��3C�2l5��!��U�t@)��2E�_��q���3�,�3�����63ʐ��̤��[3P�0��@��G8�v1,j�uwkf�fy�	���o��f�����'#�,Qo��!"+[�=a��zo���4kݔ���{f���a6�*�ɣ=W@�$v2�`�Bh��RyY?�e�,�|�C���&���o��s|K�����%[�%.�������M5��]��A0Y�<���-eN'1��_DJ�)ʺ{)��v�Εm���2?bd1�3����A�qGI���ReSqg�d;Y��!w� �1�9@�־�M�v�o��I!��0��A�\Q��u37�(ī�	��3Ł�~�h�_.�Q���;�,}x���1f�?�8^&�"�T�#t�1��d`F���@0XaR�g�y*͛�����Bn"%�ʠ��MNҰ%��|�o�5��)Ю?ߌ�Ր�rH���S���q��{p��q����-�R��@ �.��f ×��3�� �w30��~�g���;����4C^i�G��b�o,��(��j�+\�hyN$�{�3E֍�W�8"�pd�-U�� �{^U���+HT��/5%fu�1��G��^E�4<�j`���
eT�fz<b3D��f��ݩ��
�j��G��$�L���ofI5B����䮊×����`�1U�G��m�7Vo��`=]�A)��������Dיbϙv����n�e�P����puvvlTpn&% M�w�M�ͣ��O(���J}m�E��sI��$X7XvSu���H���Kr�U��I�*ֈsQY ʈ���O����+S���{��&a�Y���U�����Z���d֋�[R[$���
�XD;=9bl>B@�X�e�]��ݽ^4b>�N�36�����TD�vb�8�M۷ˈڽ  ��	����G���'�X���gTF�8�HU;[f���3��*}T���e0�e�J���z�.A<��1"i���N�0�5��!�&��(�*�k���R\�e�B�9�O�9��3b[��G�N�8�kr~	�Y�k�,�?�KC/$rU{M�h\EA�`�g��4FE�j?�NB�7��a�fY��}�%�H�I�C���������@}��zH��i��V��ǵ��!���Z��ثE���3�\��Tc�V�h�>Y(v�	�6�+��,�HL����B
�$�OB|����
0ge�����1��R]V�;n1��R�� ������ i��?*Uz�j��/x�=^bU݂ �Iu)g[�4	�B8~���&^`;9\���<�ve���z�n;H
kK�u٪7����}k���)4��rƛ'��dΘ�2>��s]��ú��AsԺ)����[ *o��r#��	��M?�>��L���KG�R�7rۉz(�WX�~�� �uj��P:�^{vU�wV\��Ъ.�����.�W�Y����2Y|�9��L�	@OF����j4o�@��,� �"H\%�_`��-k	~k��~�\t����d$h�
���٩:��k�<�hR���T}�v� 6K���N>���֔�T��̝�32�lR[�˘��9[�k�c+�ю�v�Mg�
X�Y1*.��Q#s�]���4yؗ��-����w:W����J�ֲ��}lљ�&�0��{$=?'��.�	*x}O�mN�Ѧ!�bɟnW�{A0�V|/M5� �wx���p��L-�ן��M�P�
�tn4�t�0�N$/wd)��<�0��l�>f�p�AN��</�(@�wv(�]h�|�`����=Q�û��i+&��bc��m�F�?��h���+������E�����sD��=]����>�p���uP\����Ez��K;t/%�a��H��"pL̢����I��;!��������z^F��B�_2T�p��'�D��1s�ׇ�u��^�	�[�.��@eSI��_�?��F�"��qh��¯- +9Y H�
���WPaTܩm��L��R
4�I�#��J@�ӮNʘ�c飾>p�$T�!��|(=��#L����g��1eǫOӏژ��F=�/P�����w,4o�%��@�Ο��I`�K�P�`�8�uU-���E�
��衈��^�a��U��Ho�m�����).��^TN�bl�c��!	��R�h}���� ��du��#������/��kO׉����J=xJf�nj��6�����sG�i5���a|3�%x(�{[���8�=��'�F����ڍ�ˁ�d�t�= ���˫�G)�I���K��F���kP���F�wj���=�+Qk�������+X݁w���}���F;��Y�V���]����W�$I�۔e��Ȯ���XE��o}X�PO�e�k�����N8E����f�9Z������ޥ/���<:A�E���Y\J
t�y��/јEmo 3Ѥ���Y�1��,ˈ���h;���3r���l7����4��p�Qjx�S�AC�?�l2�*�4��P��&�U=#���C����{�q�3~'\���L��_��/��G�o>��DήL�1Mn���7d/�Zr#Z��4��(ܤ[��o!�&tU��#~M(te�
��)�}m���os��iX�2g O��}�Ba�3���8�n�pY��z]�������\��z��y�F��"�&�82J���]�����b�-�{��y���ǩs�?���Ay�;C����x&�N:jN�6��������W�u��S�c���mՄ�K
�WA������I?g����X�E�Zh<_Y<?�����I�}9�5J�7	Y�����r����x!U������里#6.xp1�F^A���������'|�u�x��r#W���j��\�ᤈ�
��6>G�dbN`���G��֖:��;\;M\qf����v��#=CIh��s��bk���Ȱj�������BN��Z��Y�F �C�M��V��t����]-VTM�~fW�{��Y����&�@B� �ɋ �`͑��Ka�/��w�l�Q)x����7���!C��p$�+��Jh֊��1ދ��m�q�C�ƥ1dDa:�jUȏ��"-X��d��}g�xG+�Z���̊�z�u̱G���e�i MQ
�ޗ �i�߷r-���K�m�I�͍�-z����gL�E>x��-� �;�%a��
�z0�nb^��gm6Ě�\hY�1(|������DM��YN�K�;��+<��\X9���>{?H���	�$��}^��wU�1Y-oi�w��Fl�l���c��^sΨ���T�����!T{�2\��4}�D�er��vS�΅��<�W�2فQ9ntCa�y����XH3�Яh����F�	�^>P�^��ͫG�S8p���+a���ng�}�p&�?�io#|���h�c�+l�<�Fl��f�/�G
�' lH��
�v���h�+C�4s�l��Qд��K�G0�3hl�<H�bo�Q����-ٜVW@XA�%�Q���[˞�<l�� ��t�5�5���Q'("z7�x&ͭ�mUO{���p�'8���t��s�й�u��� ��3e��{gM9
�S�-�Hd�_����{"�&��B�v	jꋤs�>=��l!�z��3z�*�.󴜥l4�sK�vqx)��z⃤���%�Ue�5�kC���Cc����%��1Te�|��;����k9y'��ח0��I:�U�f:�٭Cq4���u7+[�rA�f�E��p�Κ���r�)�(܏��wM�DK|	��D�&������R��+�Ug[��Y{���5�Rz1k��!1DP�@7�d�?�'�58BT.�R0���X�))I��ѻ��I���S/�)��J��O������)ZR(l�(�mc���������ES�\�p*��\�����uA�biNu�ˉ�Zл�]0���h�pʫ�4�Ƽ(��3O
J�&��?�O�%�c鑖�m8/���&��7|k�*�YUx��v<�?dB�����!��1��k�|�X�G����Ǚɞ���g�D��u��f�p+E��HD�7��4ߟH�%��xӛА���TCi~�=�#�����`b5,y�eV���Y�8��^���Y$����s�X�T)��m�0?2_]@Z`E�V9�w�H7�}�h4��h�=�t� ���䁍�-f�"��e���x�=<���(�~X����aw�T�Y��XE, ��9?H6"f��<BQ�Ϥ�FBٿ��յfv �[/X;H_o�[VP�z�R��$��bk1��M��ji�f'(6r[tCP&�xٽmԞ�����Ig�A	O@��l�7:.����Av�dxѹ�V|�`w��ƫI���?L��λ$P������=��։�ءΜ[�]�Q
\���*^4	��V�9���F5�N%�u�7ǖ����^oR0�!;I���pBP�;����Ǧl�����h��a)�p��8{��
6�Ij!��e�A
�B���0�������3��R_��+ }?rw聨�m,���;�^�v.{�U"_6��*�і�+���٢��o��.d�x�|yu1}Ϳ�	��o=B�ͨ�Q���r$Z����F�D氞n:͟Q�qz��=馺�����������'r�ԏ9m�z�X��w��윚k����6�.����B;�[W?60�'7��\T�?���Q�.盼�h"�f��mrc/�y6R�J��R�F��T��K_ìGa��>��i�>�������]z�i�eKz��T?V/s�������R�2�}�	9{���R�P&L`�B?;�I kq�����y�z`2i}-�A4p�9�O��p��#�+sW�134�#�h|Q����l�T����PBV-�zN��	��?Ú�f��M�.a�ˮ�U;p����+�4䛿�t���t�Fx��X��F#(�K��@�fӆ�;|I�;�xuOJS��*$���\�E"D��=��g���83��z,RPp�}Kk�\�f^�9��e�Z�]�a�Z���L���Zü˼���bI_��X SɁ66g�@M���v����9cs[,;z�-=��jp�şD�t�X�b���M�]?|y�#C- 4A����]�����s̘��\0��)�U�ΥڙVc���xҾ���:�}Y!;˦��;, e=�V��D@��|��EI�l��Fȩ�x�R�����������~�	���#N�*b������c*hZ��B�ܝ�
�7�x#�d+��=�$ɧ :e�p��w�Fhx�W���xq ���}y)H_=7Qx�ylo��7hB�e�($�V��ǂ�$��L����Zx�i�f���ކ�s�.�
��L��|UeHT�
�;��@0kY��#��UA�X`Ֆ0/L&�!�zE���]F�y���:�Of�^���2��d�$~�(�LPƿً&��;m��\�����2�3i��7X���XYڥ#z8��<�ON���(�c>���[�m�����(�������q���b:U�`m�z��|�k�7�"����Ϲ�V?هv��A�0�p��A"6}���FK��y,��cBc�LhU�D��KqI?O�Ə�AwJ/�
�+^�H��V�.92�",&�R��d=n����j?����L����S !�T�S �L��h��r�賞%�����a_���,� &C|f���=�వ��+	C����JS��r�<nl�F�d$�d��e��j�!N�c��u1���Ԏ�e�s*xL��T�s�D����?<��F���:9�4p����̺�9�}�P��F��#�hd�*<��
���f��L`G�!�Ԃy.�5��F� �^��Ab'�-�K�E9NjY���Z��*n��6�'ǑEB��d�QqI����m	�X.	4<�Y8��)318w�+0\���|/LK��hঔ����(?d
)�H��z��~��N28���z17�c��J.;)�dc����OI�nB�C�f'n�#�V$��%mWKx�ƼyE���9�\0�1:|��4y�L$.d�<Ϲ���w���S��Տ��G�Q�V-}/�L�S�
־MRg�E��N�l�E���yw��[����
�|oK��Z:V	�b<��H��2T~�ɷ&����e�D.��e��Y�}'�"8�j	%�2H"�ր�2,��^���	�n�a��J�Ί�T_���OEX��{,�{��V����P-g��"��72�+� ��s(�Y��G\���,w66]����V1��s����i��:2�c�Ja��4*��w�>e��xm��4pYk�]<�]m'ЋfPT��O~O�B�"J�m�!K�<Q�@��$
Q�j���1�[��e�۱���hX�;Y��`�B�L�t$S����ϳR"�ޤQ�%�2�zя�9�ݶ�'�U�JJ���L�#�.$ LB��ߺÆXM����guF,�<��z����K+�m����\W���]����+�(�����s{x\��!ˌ�fO�i�{�S	m���S��<X�[��Ԇ{Ar��(ůi����z?]��'^@V��O�Ow�C|��[X7���d[X�T�G�C9�.����^o-6�q�D�����/�Em�T�yK�{����"Z��o~���B6 jﯺ��ݞس��"!����,��3̘f�\�]��K��O� �B봴�@u�.�d.nC��7�3�=F���}0,�яb�LQ&��nU�V�2+����5�f��9���qU8q���G���B�n.p�JI�?5M����4�IRѣ2ԇ��	�|��["���Qt�C3���Mܲ"�G�pE���Vj:߆��v��vҾm�8�Ԥ��4{6��@eݶj�3�®� 	;]��~S�*{�S2䵆+%���$,[Rl�V�4Hc�����Xل�k)2�����q!��\�<<\Ƹ�]�^��U�%5̚�hLl[���0cs�n�0�rQo8�#r=f��'�rԳۙ#��	�n���_��H�|2T���9z�u�=̚޲NH��!1���9e�2t*%$��m��;Ty��E/VL�,��B&�*��iŏ_�KQ���6�����S�0\�"O��VNb���<�t�Kq�}OȪ�ڣ�Ʉ浰o+P�1`�����!�&��QV7!��-���	/#���'H�����Nj3�����)q�{ݫ��T�Z�DT��gڳRR#�YQ���+����q68O�S(�lꢱ�=�-�`P}��C�h'��o1�N%��r�P۵BT��y��W|&�3����#FdL�Ǧĭ��_*p2k�4�ZRn4D�c�*�p7�"���{C���D?�)2�{����c��O���E����d����"�d9%�;Vy{�5��(���e��A��V��Y߰��yI(/����P�70����jsxM�9v�*�2��)�.?5}yݾ)eB�E���䅾>bB�V8�F���Z{_e�����A�(��]�W�T���H-zv^pG�Z��g掊V�����]�ɵ{���?ZI�(%��g\2�����*���y��-��)��<j�1��do���w?X��&��#���hD��f�i���u UR�(X����E+�?�D�+L��b�8���\V��%��/�*k^���"3�1�SA9Ի���IQG�_Ee���N��+Go"�G����+4�Q&��ߔ�Of��i��"{ |�+JJ���$��zD�4���h�.�[�rG�,b������H����~3^D:.��x�xq�0��)S��/�P�4Y�4p5)�J�˚σr�W����n�)�ӱ�z4`9fn���n�#X-��]�u��=����<�pY�����Щ�~3����Gt4Y�hC̱`}�Z����U
F� k::`�$�����̀��}���� ���g[�چ�.����G�ɧ(nˀb���D�;����n�%Q�
�������:j�Ў������aE8J1�"�p���K7���$T���T�#%=�'Y@����h���2�� w2����b
���PF|����Zap=�N�t�h|u��y��%j��<H_�V�VBJ&tY�ļ�\���� ��o�^�{$̜b�Uk��\u�wܩ�7�}�bZD�^�g�鏇��6�����Di�1���k%��my��yi�P�,�YQe��Z����g�
J?��ߙ�*/�hL^r�o�7M�v�/k|y� a�LF��@�:�EY2*�|ꁠn�� E�0XGT?��:R�_�sߘ6�	���fXȎf�h�T�}1�kԦ&ԲΏC
)ǋ}^h��S���)�K�qD¼1��{�4�㭱)Q��`���j��'�b�Pxљ	i}�v���~�y��T^���>���l0��O&mJf�7�J9��W�B]ܜz��~�d�}e��mƊ���e���-Bz����mS�zw����i���m�T�COU���ǅ�
�����%���~��j�4�#�*F��EF����%i	1�G��1iYw]�Ske*oE�wB�,��KE4#+�~.�2鬢Z�1��x� '��*We^�i�0,��`` Ƹ.iO�UZ�r����~l�u��"C��o!�����A�W)ȶ�@?�Q�Z�<ͺW�.~� JE@���o�P�#v�2�;7�H=W�k��9��S�w���s�w�&�c<��dP��M/:Z}��Jx%���!��"��p��^(�W���-W��Ĳf�R�����9LH9M�v��ã`�OR����T���������t����a�g��
�ȷ#�{�k@�^�1"I�������9Uɾ �r�K#rϷ����
��ދ?eh�/s~�s�"�a��gw�nS��K�u�j�Vs|��B��C�,��nB�1��V@l:sm�F����.��J�E��t�Bc�*����>=�v))���麮;dם�N���Ҽ|��XB ���5�����臲�W����C-<���h�����~�Ce �8�c5оv�󈌻��~�Kr��U�5bh�p5�7���F�;����{�Ŷ�C��à�@<Vڽ�LQ�Ts�k��l5}��#�MҞI��a������Ҁ���H���'^le�\�aGٸa�:��т�O�dݠ=��_��s���OO/�߃���h-�Zc�a$�m��f9�Dc�7̙��kc�����[@�-i��:dt
&_�nSV�M%�,p/4��h�|��5�_�m��u���Y���-��{
����Y����"�����ou�,���/�eϏP���؞ʓcƗ4|��eQ���}����5)�ތ͡�H���
\|�^7��m��͐��S�'�U� ��'�ȷ:;���L��dvCR�蠏V�
���x	��V�]E�-�:Ri�8��s�9v�vC�XA�lUI�v�.��r����T=��%��������u1�"���HPPF}g��oH]�̀P�~1�%d�t4��ӂ%�a�0v����y{�[K"#���[�az!/ Hx<�~�Dt��PZ9�����ƍ���. "(���Ys����ƭ�n�9�K�X��g������T����%	��we���߫"@K����P5�t�-<�![��\욤�4c)Q1�CUe�q��q���yJ�(���;>��أ�����O���s�Ӎ�X�6��f�f�M�ЍÃ�X���E�Rxk�>�q��f���I�
��_��dj�uH���ʠ�I	AH�pp�U��\zYz0%�U�?�}9G��������|�4�'V<���\��/F_����M���.9��=A���o�{B���Q|}���M���K�l�O�!1�n=[>d�`\e�hHJ�>��hg��� ��\��5� s�l@�] ��Pm�pT��0w���[b`k$e�+���TT��2;�z�T�#<i�&�T`A��bj[�%ӊ������G�����Jw��s��J�} 6.�	IͻQ_4��,#[#����<�Oh;�SU���!q2v��J��ɑ�#
�w�:d��:���U	�)���[W3a�n�����h6�*>�b
�(��h�^�ܘ��
8@Q)!|JB��v�MT���?�
�`�`i&���D0j6���B-���_sy��@���9f���r���;�\�d�և���N� k>Uc���:=R�*��C.�a��ߵU�Xka��:�����廜�[�}��X�c4VS���YT������c���n^˒�"�vF��QBq�� ��^�-�9��d�\�,C��CL����M�|�+�y ��[�+h���lMT��0�K�K|.�v!ڜ40d[hR�3�5 8����c��Ǔ���Qa`:��w8([�G�q�$V����� �^j'�2����O�v�� QG����� Y�x�����3+=�~D�tQnH�*�������qV�<��Ք��E�F�n�l?�xUO<[�]� &�����o��M�v��]1V��0'�MW.+��S"�Ӄ�Q4���^G�'��d���̨n��e2툊�AbZCo|y�0N��V#��K��N:v6_�	�'�";g,������R�y!������v�0��E�QB��ƍ�����0�f��7.�R�k�o�|\Rd"L�[	9;!z�Od��3m#7���1��ݒm���K��
�Ysp��:Q����K̰��0����D�k�q���!و:3���\�(�{�h�Ǟ���r4�ǑL�,̅�s�Vl�^��g.�1!��Rݖ��0�BO��5�6M$.���^�}��:�d�(v��:��E���[���^��T�I��/��J��~1$8�棣	�â��T�,��n
7��J�8w�#��
tU���N��>�V��
su�4]G�'ǥ��g��[�λ�Q6h����w�I���w���i(�j6�.f�#�$�ӢGQ�,�Va>j���-n���c��ψǸ��-!���ff���'� �}�r�}�/�[ì��������r���j�3�zV�����1��HOG�^�������B{���z���BK�E5�T���?Ϋ.?�(�~�����Q�Z}#@?Ρ�.eR��O�t�|~���'[c�b�o��<�e��3��.'"5͗,��[�A�^iխgѕkт�FI�t�QV���}q��&���=߄�C�!Lt&!�Q�4�E�#^����4����cv�k��g@5�Ov�թ�����1BT�0�nw,���҂�]<�6҆����RL��y:<�f����q%w���F��K�mP���k�˚��&{ ;,�H��t���a��8}O�̈́���j����z7��ϥ��� $9�����%b�.�΃�F���ӑ�>b�k��)!1���Wl�x9+ }s�W��xȆ�*_&��C����0��I������[[t�X�P;�J�d$�Z�@��?�4uH?"V�(�r�3�T���|���y�d�Ef�T�"��5��)~
�5��3t�B�� ���u� ������w?L�8fp�L��e^�K7�k�2����/��Ku�7��;�����!���R6�Ά��cy
��w'�W�hQ��4��@��q�5v��v�hy�Nc��ߎ���%��p��f��AW<L�O���~Y��3��z���$��RI@8�7�I����z���7,��e�D��y����گ���9�wOW�7O�躭� N�p�;�h�T���to;_m�-@p�����Q&�epvM7�����~O�5���5o'
*}�T;5�Jj{�f�B�8dE�ܐ!L'Lh,��8����](1��tr�3�~�8H��M`t�I�hF��>':ԇ�����6�Y�ܬN˹RO`���K���NYY����3c��x<5
i�U��w(�4#�M,>xѵkd�|t��K�WY��d,v�*s���shƌ�Ŋ�Zc��f뷘���[�
��-8��Ӵ�Od�4JB6�<�#5��ǽz��A�p�K��Ԃ�6^cDn�8x'?l,W)[l��f�Ʒ���|�,������ߙ�8���D{dG���))E�*�"ik�M�'~�����J��������LN� �s��� Z�g^@&_���EʯJ���N2�Z�Dm�?�a���H������o^��������칞ј����e���M�y���F���D]�d��۪�ᅫ=����<Q���I���:m2�l�
N7�XƜGN}<G�z8�Y�/�����{?�
�1�%��%�������U��k�Oe���5�bӍC�����6��(!��>є�a!O�Ys��슙���$-FB�)B�+��RW	��@)x7��)��G|Ј�AV�f�J&a�F�s�e�X�@2��uP{2�q��M�*|�~���)�9��Ձ^v��l��",���Q�B����ep���A{��H�āE�q�������,+0WC7�#@U��,R��e|����������%��OiZ���
D�����?�6l��t�,����zQ�,��w���Γ�L�W:�S�#C�9C��y���#�h�0�T"��*���7U� On$f�
Q /|��ݹ	i�!�a��>�K{@7,���Y��T����#嬐�_��O��*ee��f��j�EB�Z6�8�m'��?n�	�C.ꃄ;!�8Ϙz�����z.]���uwXc!q!�6���ؚ��?/ R�N�-j)]�ϕ�T�����x|�GA�|2I��*( �+�
���ǲ�{]#�Px�l�~���S�#˟�RV�W\�u��&��v��KaC�E��M��cD�a$�٬p�4~��ށ�u~0`��ޟ��V�yy�"����~J��|h)��S���X�qt@bѲ�}�@�|�S��2�PR���՟-��������.ⳃ��s ��c�&�u���˻Lh��j�N�������$��F{#�s÷^�Qs�Z�*���W��0m��y�M�k��돓��g�,�Ҕy�W�����3ܩ7RFYH�ݿؚ�Xdi���ă2eN�_�U�XYʏ!�6u�*�a�Z.�p_0-���r(j��rr�,�hY*g(��n�ӌO�������(1�H��^]�zY�
xe18�}�խd�fQ�^=Ȳ&���ԥ����d�2�s�0�p\��B�u�Sn)�w���HW���u��/j�4���[[�]��>R<r'�4P���PwA��׮Y��\�r��{3,]�U�^����4[\p��F2B�`�JSP��1�O�hZ��P1H���ν�l�[�t��VgUg�rЪ�61W"�v[��v�hk9~*�}��,���<�b�^*�%�ۇ	���|�������_:;�bY��gf��gh�L4W���[�i�N����b�^(}h%��8��O_�+��(�]77 �Z�C�KSk���3�o�>W�J��E�qy!)_�x��і�&�f�}��!����S��x����{�mzܻpIub6�~�n�n���p��0�<�<�r��?��8e3�f���{���������4��t���c�+�j���A���ܦ�18/�|�d��J�	����$+һ�6piD�~��[~����j9���}�@�ind�|UǔY�L/+컄��� �d��etz%F�w׌, ��}���ީ�1g�]�a.�/�۬VJe����դ'q��*i)?���J��KE�=q�n�%�E��I��÷a�y+��y�����n�؝n� ��V�[��~Z��qE=$��H�2��^#f�M���Tͥ����}[�.)z	!�#�/C`\&�FB�����/�Hz�^��0TfS�@�륿Y�l7��F�$���G\�>�ʠ��8�M1cu�q毸0+<t��U�CUڝg��ډ��ب:�b��x�/�`�;k_�<�rL�O�h�}E	��d��n�B��o!Y�Q��ἧk.���ɭ���|7�L�;��A+}T��R�eJ��v�v�����~�ϊ��+4(��Y��D����]O̾�l�O�5F����-HU:�c�����;Z�p�S���
����Q.������۞AL�����R�q Cy�X~��uf���/˽[vji�2A���@>_����fZ�k]�H6���6��`�Y�@��%�g��d���1$�uS��E�W[��i���j�q��۫o����@���o1ļL�@$f���\�Q�;�����r�S�>�Lv�+�
aā?���i��Zj��DoGWd��'H�>kuY?�7y���	CC��#s�O��1�*�H=��5�Q߂h T�b��� �l�t�pvq�F�Q,H�d��;q�.���g��ƚo�|��H"y��3g�qN�i��~_~X딒��H��C22�B:z�s"N�i�=ku��lw.��,���(T��W �r���8*|��i�K�ۆ'�h\1rd��G�6W f�fn ��Զ�����_o9b��a�՗]b9���qojث��c�OK���ٳqW�J;��wae�o.#�~�T^'F�M����`Y��uҎ�>>)�"�Sze5c����JHA���/���-3OA]��`��3D�b"�����Id �'���vӐ�|����EӔV��!e��RnR��.{#����u3��g�3��%��8qI��L?�G	BA&Q�Y���Ϲߌ��mf�j�}(��	���4��FFp�\g�I;'.t�gv;��r����9���1%��r��CB�����E�`��H�K	@)֧&}HB`0��8XCK菾F����4p`po9�**�0�:�gaG���%B�h��P�*�C�PGB��7չ�Ү��M��t|�P�Dޟ֢��ĩM�@�>(X[�h��IX��津h�P~|ao��(˗D]�h�Mh$,�!�f-��sZ�� ���t�����b~#^��WM�z�ճE�u���+��L�?�gsn5Բ!O�e�E/������r��C6z��2���>�ͮ8�\�����Ij�lt@�q	�̈�^��QKs��m=T���:(��՟~�t�-�<k ����ʡ�
��ɽ�x��v����|��?�v*�>aϹ,{�Ե	�� �A؂����/?!�Fk/���A�B"%�R��
E�20��Rw&����~��N��hn�+�%�c<Y�S�Yf��0�����@l�-$Rt)�,��1�N5��$���O��F^V˝���¾>��c�3�r;o,Uv�Ώ~n����rb]��"�'���@9���?�����!�3'���D~�<����l���
luZ��UK�̶��?�j"j/i|��+�4!��cxϸv�Q�-�[��-P{����靛/|���'s+f�֒F�&�ً�a����t/K� �6~׳��L�Ϙ&;��(��uPLq�-X��q�O1��"� ��?�N���[���!�+�P�Mld�r�A:�Ng�rܺV�Q������f���]'�Ȟ�>���u�я�c�R	;�J�Y���6p��n@1��O돿p�+��=qほ&��`ZKr�Md9>��W#c�h��XV+H	ߏ��t��Q�G���]��b�)�:�a���_;Q(�ig�Kp��η�_%�_@���3�zG����a�s�wa�!�m�= )�-���a��t�)ĐY��j7�чӒ��	^J�$J�.�53��1�ҷ{��^��6߀�8����E}�f�����p�x��wҋ��)S2����PL|tV�n�d������Y�jnK�����Ζ^��q���y?4��	��zQn}+u&������ƺ�!_) �8V=����H�ݫ��L��hm�_;M~��̨&��Wbs~.���Y�N���j�3X��ܲ����G�!l
�/�)D�y����r�1|���{ �ʙ�E�or�߭��gm�����$f�^؛)�k}����	�tF��r��lZ,ĸOT ��{�'@���"�u4n8'I�O�&h�dsI+�j/Zl��z�7_@���0O��Ќ)�|�'������/���Ҭ�T. ���x��yz�=/t/��h�o$k׺�����@�Jg���5'1����3
�T�v�?[�N{�@�;�?ˮf�4�E��0�T�,3��&Qᤥ�`�Ph�w^P:���v��tpV��w���0�-��Tk��T���9M���i.V�K׽����y�s{R�dn6+++p9�� ^��
7�J	.����Zs�n�"�|�en���O�?zq�s�C	�'����)�r��=���l������k	�o��� $͉�*L]��!��m�<��o�}R�T@�څ������U����Uj洢�<8K�kF"��:ݥ�e�(�"���K����˽�˛��q�d�@�ӳ"��w�#�:��ʕ��2��T��U_g�'K��A��IK�ΚSd��7�l�P&���*���2&�n>Rm���%�"�M�D����48���f�	��v1��i��⽻�v��op5�D�l�g�y���g+��
���唞����#�2*�$�G&� dG��+o���|�GI(�u+��"���,Bc�hŲ�����߸ɼ=��3*3�8c��P�����%�Td�ANE�X]���o��p��.%�zTA:��H����7d���]�p"�M��� �]���+3H��5�#��p�X�_}��)׹O����5(S��^�E������-Ⳟj�߳��\��>e����G�1TҷtYB�r�|�J#�T�P*�mva���1-�-�5AG&�1B����Ҥ#{�3���N��Nq(�(mfd��Q�����=��gd�:@��S%Hc�~��o|�Z�j����X"�����4�G������df�B����3j5kÑc�}��h�\pa�Z�mq�W���W���E��ywojWGu�K��_o7zT=8BI5)��`�M������ޫ+
T��2@�l��?�%�
�6��u<Xc�Bh*_juj� 5	���	����:q�����p��iW9~�x����/�:T�qs�ܛ=q9��ܯ� Hf�K� �#f�b�.l����r�I�ͧ!3�>\ �b"m���G�c��L�?؈H��n{��+�-��%�b��ׯ��Ubز�L�a�ѹ)z�G���
d}�p��B"��f�"=0��p�_t����2F��g�)psB���������b��A�N���%�$p����<��E���cɠ�X'1��Q�).�/fVk'�dD)�cv��!����Sx6��| u򈒤,�������G2e��`�|Km �ᰐ�=�+�I@����Jq�>�u��W�TZ��"<�։����:�8UB��B�N2�2i����E�=w�X��{�|�Eu��0������{V9��^���Td��t b�K�3 Ӈ��2;�`e
�PR���[i���(�8(�R�X�B��)ϗ�ߝt�F�p�����(��`���*3�+],Y�;MdljO��k~N	piR�@W'�Q�1�J����m���9��X��]�`27k��)j�xXD���m�{�FPpU"���=,� :b�����p��NRc�^�ʲ�`{d�d�_"�Z��a/�6��J����$(n

j��U���U~���2�|4�e*9��Yh�a��� ����!�nf��o��� 3[
�e�l��j��ws���/�G�ݪ}�6|0����vZ>+�S�	�/09�� �����i���H�� �.�MG��l�h�CԐe�q���}۲��e��@L�����K���qU'��R�k�*��F�I ��	�Lt{�	���ƨz�A�[�Oހ�JS׭���y�,3s�([�q�ɳC�JX�b�kp�\w�B������?�FfȆ�����F�GdBR��ϭ�nvg4�d���]�^��!>Z�-��]OU-V B~�R�L�o�U�1��K�l�o?��#��y�Ȑ���ߟP��A�u^z%��@�hJ��,9>�n_�;m�p��պ�󬑔���ι�4hw&�����]���v����%���t�7�K ���9���nlDF^�or`2uf��N/B�ɉ]jWD����>���]�¾19���,�?p�mϴ�Fĥ��:2NN��s�8�{�ܺ�|  H�B��n�~��w.Bo1�L��6?�=W�e��C���T�T�Se��u:4�����~H��C�����ނ�H�5Ș%"��F.�^�!D#�0{��9�v��`p3Ӽ�ΙrA@���n^�3�ۧ��#T<t�L!0��^΁`�JH�_�Av��q{���ٽ�&!}���$�Hd��{5�i�5�V����g�MD�*��'[b�H���m��j{?�vD(�"�1f-�.�ܡ���G֏ty����̿BƝ�R������6z���_9�H&����l��P���_��������%�l#r�r̕^���R 6�_�}�}�Ҩ��F+�u�q����X{A<���ۇ�B�f�Q�+4�ސ����b]��r�_���Y%���7� /և�}�����1���h�� h9
"̲��/_�S	*Q�vW��P���X��`"�D4�%>��������	Xf���E��&������"�{�O�=�g�5v�&y�Pb��m��(�r�8A������tzh�[�o�qCs�93(�yDn^6JiJ�#�l4�@�`D �X���<�WE�z��[�������Ú	ٓmH�{�S̍��QD��Ě���3G�'8���L�:2)ґ��l�7."�ky�"آ]�~��q���ZI�[��ow����]Z<&���T�E�A�g����z�]O�b�����.���*5��F�L�>�5.�������l�n�&i�!�'�Q1g��f 6���dR���2�
�}�5mg�xE,�Y����Xv�J��6#`��m!�$��:��X�[G7S�5�[|��/�J��bGJ���E�)XнӸ����`g.E�x>�<�`~gɪ�����p�)�i{��3/Ȉ�n���s5r��d���=W��kWD�_��q�sӭ�> �v�a��<�ڨ�����)!�"Z�h\.t8�Q�jfco�.!M|SyK(l���'Cs����cfG���u�`�{�{�.�0L�ML^�G����!I8���IX�r{�A*�Z���N �1ʠ�.JM0���39M�����48W��F5�BX���|F�lS��:P`�.��ied�p�;���k�H7'OϥH�Lq�`D El��#�+@J�͚#7E���̻(� ���l��L�K]O���	~��i P�F!,�7�q��>��a.�7��k��e$�y�N�-�MX�z��z���C'� �x��EF��x�ܥP=k�=tj�de���	E�`B�!A\ٴ܏i�^d�\ �����p�$;�t+*.;�(8h��\ZZ�Fv7�7x��iz��n�Z[,`����`��@��y�=N�39�q�E�͚F��<�t��>�˅T�lOȗA6���9I៼�8�x w�����ic_�s�J�޿�4�D�{���(5�1�r����j*����g���#�������v?��D��,#韯���	E���y��>�U�AbHm	�7�'˃�h��J<�a��'5�����B;��gRvռ���6�D^�8)�m�1�K�����P���%��+1�I.�	�p���p��HGv�Mν���ft��r�t+&�89�V����@��4J��i��{�rS&-:���0��E��@	�C9
\m�� ��}��վ�i�:�|���k�oW�����7G1� �ax��,�<�;qKR ����ݘ�Z��)�)Y
5��
�X�L�c	�eŘ[�+�I5l{��x� ����*��Q�9tZL����uŘ�9Vu��j�eN����"ӗ=R���l����(�,Mt�}s�����i��̰�]�!�2:U�6v�Ϳ�4e�x�Z���]X��ĵ�e��a5�S��u��ir�H��Z6��c���(!D�A�`x�s]j��aU_�>���׾����Ik���s�ɄΞ�}k6�
u�W�Q�Y@ە�n����W��r��va �}D2k�)r`Y����<�D1����VT��҈�*�i+(ݬ��/]"̣{r�Xd�����P���猊�;b���X��T�&���ftà-i5'��{�-��e��[�G��Ou}��g����>/j�P:��+RV/��!��0���.h�Vvc	�|C^޹�.񻠕�~J�;��|n0�f�fpЕaEs\�eL�xF�c����]�װU+�}-�ha��� ��ͰV��Q�]Gz�Ow��;,���٬�ރ�}����;.`��V��f�y.�v��07�,�������;��8�}>rD�����{�z�*������r���a{��d�^_���Wi`����!I4���o��}Hl����@�����~T40ٯռw�>:��. `{�F�ay"�O�pp�E<�v<d�|m�c��\�":��'��������E��+�� �+a�p$�+��W���[��ٙ���g#EFG0���˓�` �r3pb8�e�x�i~Ӟ\F�_o�/��o��@L�D�>d0����_Kʮk���^��=�?ą����~n�����w? 9	�!���z�����K���)>�:'�B�I�󡧧�P�V� :<ʕ�5��O��.� �ch�v�lGH�;�����1����S�@�C�5l��z�D+��璃���¾
�O%��]��l�����-/J���,����y>)�1B�D��׿�$��Ft� ���vm{������޼��>�T6\�5���ݫ�lDW���*d��v��:���F�
����ҕ����B佤7�F��<�oꁎ����_1l�c��00EP�w������ӆ��� U͠9j�<��kK	�(���9��[��~�+�2b���L�4@Z����H�ܵX#M�6��/7M Y���FG#���i{����{��g�)�	ƸNGׅ6qpYd�Q,a24O&<���a�_�<Km�8X��ɉ�S�������m�2���ֳ����M�R��I<���D��Dgh'�]�@�M�Rdkz�E3{� �2�[0?n�/����� ۅf:<0���^Ԑi"�Ѫ���� wО����=�I:J�-���^�2�97������{�s��U�Wk�)G"��$1��.3�5���C�H]��lK�న��?dIw�J����U�"��:k���`
�0IKQE+�U,��5vӷ��y/
�b-�&�)�C^g�ȁ�x����k��naI)9F�M���U�iwb�5:\7�6b�_ �fpy��TX�c;���F|�Z�n���xߝ5�5�Ϣ�'�-��`��bh#��74t妠PѠ�5UQ��d5r���ŵ���Ӽ3�k�fF������W�Ր�C&�U@�.�☄ܜ�=T���Ű��E���t�����r�dk�©��H��80��+1l�7s�|2�]����a6-|�]��h�d���`��v�u��&��a�l�