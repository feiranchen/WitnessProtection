��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�Eݹ+@%$ѝbNs>�%���%c�M��e���Չ8Q�;��0A)֟ &ȩ�I��=�N�q??G�s��ˬ�}[���Qα���1�-G:!6U��c܁e�O�#���P~H���n�G�O�C���3��>��:��Gҁ�>"@�9��x���C����՚��ɛʱvvH��3}�ID0�
s���z|v��c�>��0H������v�ާ�S���vҹz��W��R�;�m�0�����3��,�D#��i<7ׄ�Q����\͒�qQL�޽	�hJ�s%�Fck��kJ��Hb����s�}�B+�|ޗ$�S�-ϖ'H;E����l/���1�E;�ɱ���B-E�� �$k{��h�lz��Ǝ�� #ʀ;+���9���AE�!l�OuYQ4q�P� ]�eV嘛�R�1�N��5M�����go�뽝 R��`��e-q5�;5둠��:q,��$=6�6�2�����%�d�r������S�Ԧ��~|����3�D�}�o��lb����m~V?��B�ﮐG�`/���E������2#�L���a�$:��bw��]������7���v�cǘ�Mn#��*��6�u�h �U��[r�c๢��.��CQ���V@�1SW�_���0�}N�"�������L<2��U���X�2�p.F+���+�kpOK���,k:5�z��ݨ�G�b��G�E��ў��7��=����:7P�S0[� ��ۿ����/�&�7p2�jm���.:L��C�͇|�<��'��3���)ߴ�狼��b?%{��L�C���,Ϊ�ק��՜땞O���;5��������Rb�C�+�WR��U�Dt�,語X����L`ob���J�Ȳ�r��<��\�{��{�nqN���a&������8��H❠�<`FK�A	�x�~x'D�ś�Qx������Ddq	.F��W�����~����"/�TIK��%.~E�ΎT�R^��.��A�$-")y�&��j+,�MwY�Ϫ��a��^�i����������j�;<����?�t�o�h�{���9E˙�3~�o�۩�fM�Un|Ͷ�Ȕ����/�AEA�������Ǣ�Fm2��+�س����l'P�^[��Kݮh��b�PĚ�l���%�
��[A�|=E:�w,UB1t��:_޳c��J��)��HFؤ�{ڣ�Ҭ�P�G��g�����=�:���ʖ�B�.�ҋ L�/��bF=s����� u �n���(��w��۞nSO:�N���0C?H�kV�l,(C@c#��`�����n �^��%j����x�編H7A�iң9r�/��@�,e
*A��0��͒�V$ͧ����6�T�w�������� e��J�����r̴�A��ض�J;޾��w�w�{p�ޏ�r墢&B�s�'�+z'e�n�@�RhZ��q̼_����.Ͱ��ԫ���f�(ϭ�=Va���(6�q4�,^�v��]�=��R&t㓐G|��ť�N��v������>�^
@��cC�7$@ȇ5��FE�YA\·�&`Q����+&[)�TU���}E��>� ��{���a�]!�~��G E�ƾ8i�(�d�%QDr��� ���x�^q��ꆚ�d��%�Z��^�;k���̌0��a)H��-��d�_��u����?������čd�UQ�gS�t1����7��3�2-��1�����v��
��tr�����?�F�ȕy�@��fi�MT�Լ���Ol֨�:o���3!��J �g�|��t��/�^��bc?��5�+�N%��ߘ����Y"���(�ʘ��NyfG�b�ApUm_!�á�0��^�F)W7+�f���r1j�7��>�b���'��4�ń�x1��c\�Bb�L��B����67���-$��Е���"M��;���^���;���5ig����s�W��|[/�(��&,"��sc.�S��.n�-��?U�����סa����*<���@c���mb��@ʍ�}I���"�N��P��"J�z'JIb�Z���\j|�.�8eTTm`0u'�}QJ�Π��{�QD���$��)=�ˏɽ��x�$ܺΚ��u��b�!`�u�(�OJ��[�>�6�~�U4����&<tyc� N��.����Pe�l`H^8��[�o�ōa�tl�R�����xT�,T�@�ֹ�WU �/5�E"4.-���)Z��7�����keT=�*�	���t��w��A�dӚ��gaﲳ(��\kn�W�\�_��+�󞂳A�s��F�`�+i���̉N�e�g�>�7�v"��H�V���B���{�,���O&�2�m��p�e�� ^�gl3�5��I�fw�y�]PZT̳ԎY;M%�}+W��va<��F�D�,�}2j��
2{H���ꔦ 	�K�����p��pDݧ Y(��Ȓ?yv�{�5��ݛ ���'��q�H>��y'�&|C�Y#s��_���@��23��p����$��A?S ��u��
��HI���%�+�Ek�5b�(+�f��o�e��z�P����D��28t�i��:)�m��b.�y�iy��rGc�5Qs�	�M���V~R#6$��e�C�d�����5��
��G�HMʅN�Ӊ��+�b��&����S��x�S��>�뿘M��e��uMw���ӛ~�_��_��D�?]���̋�"�P���X�e)�o�V%j��'�pϞ'���,�����5��ø���Շ�B�5�)k�}�("t��3s]�T�A�=���ܢa(��Yy��s-I>]�^����2n�z�VT�(q����(����C���,;]7o����r�>+�˔� ��SO�]Z��]�cX�2�M6��M�R�|�����<����Lig�OfÐ]�%��w��c�B*I~O�ᰯлx�ɻ��>}�Vi|<h^��y��,��!���}�G6@������hmD�x kԀ�M�M��$��dMӺ	��q�o2+xǾ�J,�Z�禼Ez���z�c�Zjƀ�>J �r:vm����Py��|vXܟ�f����x���Wl&�؟�Q(E��)b����}x)u�s=�DW�H	�uT
YA�WUe7<��n������>�fӵ$�P�6���q����_�\�bY�8��L"?��U�:��m��l���B�t�0'��oA>�G�o�*l�ILx_�w�UMF脒7��<d�6�np�� ��,���˃d�R�K2�Xf�cZo%5�Q+�uH�!{�d��	��I*��/>��q@TV0�󥢁�牽^\C �2�K��ñ�VrInu?�q�	P�<s�)���G<x$}k�8#��ߴx���7���'K���P��Ӑ��p9o+z TT�:&��兣�Ad?����[��_���H�ͱ�
�5u0�!��Y�#s ~�hΫ����.��ُ��0��Ȧn�wZ��f���LMë�`��U���c�3y�]��-�S��ﴈ�r�A�����0�e��u����f��}ŕ��̷�`#��T��^� v`m����m������Fݓ5Y�;:ܨc lߪ�my�{H�
5(55���#�񏘕M?h����Xpz�o���9��c�內�l��ta��<���`'�m�g�Mװ����7�T5(�9��%0Q_aJ��?<j���ksKG�P˱�=ŶJҦ�*���y�����8�3�x��	��(���M���� �"����,��� RX���<:�H4�VbK��#�mZ�J��v�+��$����c0Mk����ô����Q�s���4:��o��R��8	�B�l�'�kS�@�B���� ��2��ɿ�Og+�:��e�N��O��}�*Z&5�v'�֏������w9;�wJ����}"�IUtLL��c��$S�I�/�0,��0lKl�����L�tF�UWIV���<%-�D0���)~>��	2g%���h����q)g6ZL�q��)���?"ً�.(>��q�is�Z�����S���������J�&��q�&��[l��`n�<�W}"����ֶT���t��q�sK����̜Ɖ�d"�õ��)�\~�;&R��J��S�.�)SH�~����g�-7�t�P׺U򅑨X�Ս��.-1�Wd�Ŧz����#4���� |�~�[��{�����R��v���R�*X5l��?_֔���LYU��5_lBR[_��}]���Q���5�B�(�j	�=������N��Ke�+��M���<�o�f��D��;3�bDŎ�x��*+�z�5�eWW���!U�6���Ƭ.������L�U�A��LIρIH�sY�SWׂ̓��P?�#T�.��͇i��f0~%�V�q��P�m��}B�2@��VCq/��P%���yML�9Z +Bj4yA}q�Ӽh���!�&����B�v�h��������]u�yF�	D��f��	���\���=�Z?������~�6�����29�W�tw�;�n�q�L��;E��� ���4�$�Xr��ھq]u'�V�&3w��s)~�<ƶ�YyJ��E��������e���E�xt<n����3��b��>�!'>��ӛ�`�����|V�3�ַr�s��P�i�
EL��x(�ta��<H�H�z+Â{W3x�V�������աF������}�`��׀�5	�qX��0��YQ���'·�&�xWc>a�����9��q�շ�Ǆ	%��4��_H=]���K��Sx��+��z�-����@�H8s,!�#�`a��O�C���YN�-�e��S���M^ְ�gn�,�ox����qظ̯,=u�aܦ���"��;�F�P�PLfMPz*p�?���jKSV;�\LH,��T�WB���H�,���y��A �(D�%J���B�e�`����~�kF��R�8���G�O�E�s�q[ �w=�yv������Ʒ��i��% 褒�:ҹ9$�=�H	RIr����{��?��<��$%�?�qGl[�m�L|�O�ɏi\ʪ��f�����~ꃲσ3�����P��+���{���v��:��K1�I�f'��ixR1�:��TS���Kz�h�D�2  �͙c�b�ѢD����4�@���8^v���.@�Z�"1\\��Ipr��6�"=�$8��΀�9���Ԑi�'�{D'!
��T65 �#BMT���`���Y�O8��g�t
��7D��/�ڛ�}g����3 ���-�^,�A!_e.�M�8L�l��e�7��On�B�cp4R�8[%� A���̲��(�8`c�M���}�d2��)n�a�F�/� :h��_�y_鮟�v��I�`��5�^>���hy��m'Y	����~��4-�ylQ(}.����6�[&�ߗ��v������x?�=�y��|t�k�X�=Iw2^ei��Bk��m�\e*�C�j
�=i}<l�l��#���O{Y�ޝIg�g�d4`=V~ΛE��K�c�q�mH��U��c���M�@9���`����!R0�Kh�����t/><�,�N���� �^G�lҌ�9�6�����Yɧƌ_�cOX���ǉ������/���f�x�)�����b�ˆJm�J��m�
ߤ�U/
�z��@�����,����BA�G�n~�w��]��Z@Q~Uڱ�,���e�{Du��78�o��Lmӣ�#���;�6jU#�N�g�0d*{$�q>�9�+�_�*��%��P�{��+)��	�U6g�s���-`N�+�>��4�z�(}�u�
:T#�t0OR�8ҙ�Θ��Sr&� �V(��Z(a��B�iN�+��;D����ՙ!�[QP�(՜a�  Q�8��v����i �o�ug���D�
�������j+�<���a\ iY^��V[=�����}�h`�[���Z~Tiao�Q���д��3�� Н�e�s*V�/	񰆪7j�tbfB�NvG��=!m:�;L�I�и�Z�ַ�������w��O�И1>����Y��i\K�P���#OdkOZC�n�m��V7H���|N���4�$~։'��b�/W�y�KNj(��^Ox�<q�U����h<��X������e[l@�ux$IvҎ+>)V�@����W���x��SX�O�h�h"�P'l]���ekgo>��fb>c��Dƌi�`	�؛Ѡ�g�V�k����P4����jTJ&݈a�-��w�F?~�\T{{��,�V^�1)	�
��L,�^�a������ȅ�vz��"��V����0x~xg���n�z<��<&x�(�WoR,*|���}�H���]}�c�$�2�`i)����|(�!�ҽʆ'ik�&)^��z���/�Ux,a�C�P��]�ִ�z��@<��]m!4�d�8���Acx^}���"g|�S�yT�E����HVG�� ��}n
�##^��Lq!8�e� ��B��B���4k��?_`8��6<���� �A8c$ʹ�c���ֱ���U-G�s���f��V]x��PX�q�6�e����l
oX�@��L64Sު��􇉋P:0�S�C3<t���
,CgvA���CO���i��k���M�f44?%�.��Ґ�ߙ�PU�b 󛂼g�4@$��VáiCo�N,��&�t��+`�����z[ń��4	E���	J�]j�2<;�*���?f�Z��c��������+1�	x������ЈT+q�b��.���^����;�@�@��W���bD��i_ژK"�	Z
�g�@\B��f_$n�.5�����p�HI�}�d�n����dp�[������1.?)��!��#��s�I�kH�,O�����M�0��ZJst�9��
 �+���.�>oZh�.�d��{�|J�V�ȭ�\Xh/ٝZvV��3�YY��?��놳m��ޣw����l���'�ڈӢ.��=�"X4�%sÏ�$�G����&����^��Y��Y���;�I��=�yn�[h�2������6 �=�RN�ݷ;��*c�fj_��]Ŗcv6��W��Ӆ|g�C���[-%�?���_�6ٽ��ֺ;� ���A��gAK�^��&6�Ȇmf}����>�
���I#B�i�c�n
���7�ܞ��{X�1�ɘ�q�����hM�P���у���%>����j�eMO�M�O�j�Q�rȉ���|uY�4��G(J�JO�����e��R�����j"8�a'6���(�����z|���៵�9�qɟFG7�rj�ɗ��/������(�t�Qs�נ`~|�w�������<�.�B�C�dc�In�P��S�
୻��oa�9���"���ۭG=�z�yx&<@ۀI�<�F��Z]),˺��ƶ��c�8;ґ�c ˪���&=5ѹ�%ՏY&}�a�.�9vݫ�28���t~0����~:`<��p��6���Z��7L�إ�s�vܛ����m($��(��5�\2�lvM�%�,��J��//�]��*ǈ�h�Ks����ށ���Q��-�=2ms��=���
�lKAR�e�N���LHp)��������5� �͟��c��[� ϧ�꿿��.�8��tYٚ-���G���U�\�m�W+�&�WF�i��Kܩ)�lA5�;��/}g��!k�Cw/��C䋓�R�i�P� ͪ��J���s>Ի�.�O��9���}9���P+Y�� %샵�`'W|ψ�rs��:ڴj�5��y�ii�� +��샍�1ey�l��%��Y��Q(�f �~BPq����̪m�]l{�[�Z�U\l�\k�O�LI~�)'!���g��W�i}(z�m?\��gƭ���#Ť�aQv�i�C ���~�c��yV���.9v�@�m?Wp]��4le�ײ	�A�qE���5$B%���r�U9#��2W��%�6]\��}pl�P����~�^�K� �֬j���9A@�7�A��q/��ޞ���6�?��,]�Z���u����2&��ɿ��2��\ �ķ�D{���_���V�.yV5Oif��)k�7z!uY|Fqi��FUo����I)9��Z������ I�0*]L�WRY���.j���+��_$��`�L	���M7.� fN���T��d�8�Y2W[x�1�{����R�w�,Ԩ��0-�tB�yF�%Y��-itz�n��i�p��8E#��Eb��N�>Y�a�m`��m�����3|0�Dck�Y�]���P	Zyy�z�\
%��A˻���h���S��K�ԧ�V3"�ڌP2"O�ܻ�'b[Li޿$��FP�E�"+�����[P0������A�>jkߓ�2H�'��2�Dor�Bzؘ���u�6?�����w׿Ы�2w-�c~���p�/��2[�o����8
\�g��g�4��D��r��o�$�@�lRn��쿁pv�=*閇
m>�x�B.��BƓ~��>NC?�O�/!9-6���9>R�j>J���H5��#��)�Hk�����9:����ųy]w>mX1�!J �?��l�<���X���\+�ukB�I����7�,�_������8i0�Z=e�룗J����|���ƭ^K@��,�؛���3r��7�=��C��8LF�^�x�}T���0W7�o0�G�5O�&��{��xlkD"j���(�Ն��\m9ˬ�PlEV:�5刽P&C�f�%���οW��$���"��Y51"��lM�%	��?T^[���3|�Tt�.U��Ѥ�����$����ǳ]e`U\I
�{��&�?��4�C��Q��F��r�!�뷂�!�b�L�4�!�xF<Xi���`���V�p�!�j�X�ҳED�ش������N��r�� �NbyM�I�Ђ�*�Ϩ(Օ��b���5T��\#�w��D^q�]�}�w']�c
��qd:�}�2(��N���/ع�X[��'Y̮Ï��whg�@��щ~�3�C�rٶ���k�[d���Q7pI9�eCtig�}�0�u��(_K(Y�h5�f��0J���a�B4`
J��C@�zC�:%/z�I'Ÿv\�e}�s��C3�q��*�^��&c�{&+�Cr�*�0Yq��Q�S�q�=��jc�6��w+��x»�3qu��*\w'��S�O;"�ʟu�ы���W_��Ro���!�͑�ߑ+r�NQ�&ݿ��Yfp+K4�x>�U����c�&z|Raf>�K�o~dL#7>ۚ�
�	H�S��^���j߇�\l<�����LQ��l/�0I��SW�Y;`�.V�L���p��M
����@�n�vl��w"VQ�1����GR{]���S�����q#�'7��'����)!ulI��?R9̴�o.�Tƾ�^���� �'Zr^酏����aŃj�kw���O��h�;V<�r��-T�n`��3��ZF��4<56̈���b�S�Y��e���w��U�<=�e⍹>Ko���DiI\�����p�pFMA��SbҊ����'���>��T�9��j#�f�arq`#�@�@��U�(��A�meJ٢*xG�)��25�v<��g7�UA��a�/`�~��(_�b���Y���$��q�mKio^�g�b��uH�+1�h�\��mk[Js�����ǫD۩/�N�X��N3��oW�/�M�&� �W(��ߠ��#�X�_�r�ݔ��|��� ��iQ��������{��e����@�B�[Fβ�_�y�mo�B��$u�d>��oYׇ�֔�`=�L��`.'XU�׈�fԢ�`����9�� �T/n�9�.8��LP�9���5��.6�w��Ed�d�}�	�ޡ��}U̔� ���Jw>ԥq�ƍ�D`���.p�U�%[E#T���:�w5(�W�'Ϭ�&�ŗtS�d<Q�S^���<Y�?\��~�"i�2�v���n}���$*��/CO�W�ݭ�;����ȱV)�E?^�+�����󒐶���6�{�9�E�u-B;�S���]���'�q�Pw���ǵ��쒡�㸯;"q�Q��_)	���r�\�dK�5yN�E�3n�_K�4�q���y�8T���%�Ѭ�~�<�����~�7�L�2`9��e4{��Q��<���{��ߛ���c�i�O,k��lDR��#an��gKj*��nC.[�����X {���2����@�HK��_!��w J�mgvX�#��i;C`�R��l�H<�輚�����pb�F`b�"�Y����d>w$Z$�r�����?���L��/��=���XLߪ>6&a��WG�,�ZL�Z3Fl�	M��y�ix�
�@ŔT g`�w���3�� � z(`��l�"���,�����QT88�gg�Z��t������K�a'��G��	��>F�Be���v�A&�A���v͖48X���i���ȧZK�E�75``(�������i�"��-Ő�-����x��0*�����V�i�}�)�X^�?I�8cB`a�p ����W��ȢzP�v��Lc����U�>�o�wM�gQjQJ�o�AUb����\o~�����_�hiP)'�#0ũ���H� �m�7>UD}��_��A��/�|~;��CLW��s�u��֏u=��}�]-(l�Hce�3��ւ�����]�,�#����&�v��Ї��RE���N�9;�E��3.\��,pk�M���F�!wD�L*������<��Ş�1�:p畏Tt��[t��@:"��l�*��~��V���V�ϝ$�P���,��O0�I'>���vR�V:��^|>�'<�s6���8y��4�5
+�CI��4w���\g��$�YS���P�9�ؗmSE�å��G�4�:ey~��D$͇�񃎁�P�.�x�4�v�Й�?i���	dM�� ��Sհ#	��F*YP�2(�-{�-!uβqeE�.���a96c� �>|w��b��d`�~ ���Z�ub#�j��$�r�ˇnh���n?�s %�z�( ppN.:oO��{7���l/(>J��N�8���rbb)"T?�\����Xw�Uz�T���˨�m��wCee�m:�;��1=8N�����A��y��[����ܩ���!��"�����M���y?fz��W|@��Q��H�RE�5�R�d( ��'����,a��,��9{H���-�_"W3�!tG�s���߲�=+� ��+}		���ܨ�S�5�Ϫ�@ȧ��!������9r!�k �~`ޱ$'y���m�=v��G�d��㛄S����]���GH��%��Á�Y ^����G5��ɜL�f)���Z\�in�x����v�� 8�����n�=(�I�!'E�-�fr�ͮ���2�`�#��8jB6�j�H2���U�~J)C؊����}��Y-u�8���d9im���s%0��0z�:y�� u���93a������J���+�N��s���'I�1�R��Q�AL����,�v.7HPWp�Oar"�5��A���"�~�jbа}hm��Ɇ�x����;���@Ww�Ed�Z :٢�n1M�u�4e�˸���eh�@ٴ�4�6�����<D&�'	�iƴ��~��?>ᎆ���qqw���.��Z��hK2I�v�;��T���� ���è��އ]�E��~^��T5v���[���� _Яc�)�)��Oߨ�\K�*�(/�p����kW-���5w�G��3�D��ҧ�������pN�Ϝ���2|�Ӑ���DN�Y��������}�@Sh��5�D�?�t�����+N�wթ�p������K{D��l�PQ��f�N�#XZ ��B�)�
�C���W��Q�����E�8�}�$���J��`�?ԩ߇�fV I����h]�d�l�ۯP�­rˁ��!�͋�1�#$Hz�F��	?l�Tf9��Ӊ�U.�����H�k]�[��gvF���������5x�����դ�yh!�FℳM�aƅS�3��S��w�B��q�)P��� �:��?6eB�>�6���܅��6��4�U`��<xPբ;����ðl)�����1��}mw�y2,vO��й�	�զ�*H�AF�_$��[�*�&�q�:��t�!����_�UD�P���ul{�E�7ԣ�/Z����XQ�����V�U��ٸ�9�H����C��ց��K8�
EU�p�7��L~#�kjDS�̄	��ӏ���z���"�P�Wov*Q�0Q���-vL��8��C:��Bf�"tҦ۝
1��:*[U\�����9��B�����v����h�0�!˝Oi�U�{��.�'�6��}o<���T-ahZ��O���v���M�կ���@w߇���Kձh'yĉi�,�v��2�"[��Y����`R���y�%]O�]�����Д�lwP>KS��`w#��ݗ��2K�J�U,�ڮak�6A�%����9�}=Ŵ�o��	��w���Q�V��y]�����T��F.�	���2ʰ���2QL��	��V�vC�Ls�1pB�ExS��w��Iϳ��A���]E�E�o����\<���t/�f�%��n���Z8F�!N���7mOZ��7��u�G��o�-� 9���&�X����=��N9&�誟b �4�D��L4ؐ���3���[-��nR�L%�-a�ud�6L�!Y���Q)F��G`��'\t(п�&`���9]��AB;���L���=>G
�t$]��#b#s��h�̴����4Sy� ���<�K���dC����)��`�7o�::R�<.��n�^>��W6��;�Y3Q��҅���d�T�A/��O��uV�Ny��M��|F�yfn!b���a�Ρ�i�H35�@2rn`��:���]��F���5#M��=/Jή�`�oC)pxr`d�ϖ=�[�S����ِ8���/�w4m�+8��.��?�0J�*�s1lBy��X(��@�M�����K���y ��u��R��!�'�\�1kı�eu�1
�3�P�Sʴ6�Q^�q(#��Ε���N���}���*#$睶4�ƯH��Q�+�)��1P�>#ƵPb4��Hѡ��`���0�X�b�?�bA���ۭl�,l}���2tu˼[�9��XަU�K�v嬝�%��]�;5{��lҐ�s�B/8U�H�Yw��V_=���@$w2'8�F{�U\��Y�d�F�j��.%B)�@5����yAT؁^�Oi���#b�L���D�I{v,��2k���+#iGa��b�#q�^pQO!|kH[���H6I&J�8e<�E��"_��&M>�O<�����hUj|71�,%\�r��p=�LY��=�%�N���(�#=� �<�rP8���-�趯c�S���#h����YD��<�1��o,8�%ܜ���	� 2o��Q+ھ��c�AJ�Qe�r֐�����Ŵ�o�I\�7�&!���1��`������H�d����Mj,�͵k1���Jvh��Ə���.��>+���y��0� \���H$�k�$�]o����Ƿ�.l�6�1=�p�iع�!��A�\]-�E�a⤈aH,�eX�J��D(��q�:�͗+$���ε�$hk��԰AͿ�n��L�������m����Ӽ ��-��~�8zk���4o��z��gxm��wY�t����x���t|���%X�>�a�5*��b' W$�1���}(��5�J����
�c�/2����CP�?&1jjp !`����TA����3�M���pD@��~n�>���pBo����d���R���I��۠z(���R3R�?�&��{�
R�h͊l����0D�?��bi����
�c\�|o}����<'�����1�y�����9[%��n!�el\(��֡L�;�ߔ�*�ſ+,�	�-�
��Oܷڵ�)\�-G�fX�,��.��o�֮��4Ӆ�q[v2C��d^���ڽ�/K<%o�����fP���/���^v0׿�;K��*��GJ_���&w��&a�g�ʱ���*�"��q.�|��1��t:�ؾ�.��e�>�z1�;�=h<�=.��9,��Q�h����ƹ��Z/W�ϚF�������,vlA�֏��I�d=%�h�7=y���P��0�A� 8�^���� �R�`�7kL��c���r5�����+S��A|�X�z ��H觸'lTH};W�S�9���g�HE��®_���i�����D�׊nW#���*�z]q��~E�}�@}�J+5�K+���ߩC�~���wŕDnH�&Ӄ�g�	��>IJ���\)cƁ��^�Y��y�}��� 9�B���/�:��/�x�՗�R�<��ʀ��}_�D�b*3��ej�H��*�Ql/�2i@_�f x:�&)��ٕ��ͽ�fTƘ�X����Q͔g訰�����`������v�#����SC��ĠX>�R��G�b֤43�,rر����)̩y��		�^��ګP �(B�?��ל�P��:�8�{ÔM��Xf�Z�L˛S-��UV7(�:�.�֭X-��$#n����.��9p��C�DdL��d��&��^C�����L�`d��������Qn6�r
��h�PnQ�f��7RP�|���fG���u8/��HelB:�|ٴB!)ή�H��F�z��3B��LQ^�"��U�����d!u��_m���/�\.렲����->��e�Ke��s�d�nҵH���WF�8�`���"h�\2MZ^���p�r�#$lu8"G`��DSO2���N^J͢o�:f������l�p��^��@x����O7*��o˼&1�IۨkV�}��2���6�c$���(�����߲�R�4ѹ��I���`�u�r(�	! �$Yu�	�W��z�<[%�2 ��bw_��|3`�[����Wk�I�����Vv戓�h#{T�f�$Q�����^_����~7�&�$�>��6yB#�B����S86�d�_Cg�{:�v���W�V�4�5��#jj*��$R�����I/��<!q�v���a�V�Dm�<�Nξ�D\�]�R�R�9���@Nc��G��O�QGY�
�� vt��r�1�X�?~�4#�{�Imᓽ�F�"_$�L�M�J�&'
i�Acp�%A�x�n��"|wi�Ǽ�^��Z���KH�UH��"'L2LnL%����r�Z=��~'=k�?�
T��D+IP�zXh��6Ew�)oß�5ls�^~��j&qL�Va���>���������ɕ.'�z�F������*�%C~h�ͺ�-7��5����T��\��~F�d�W^������Z��W�:�X9�'��[T���f򌢡d�\��H3��L�qN;��O��z��(Gn�F�J��y�o�c��}p=� �,��C��yJ��?b��Ӄ�j}O &�q�%�s�x,��N�!����0i���: �RG�T��������HED�'���d�?18�Fn��NJ_�\�"HĖS_A��^r:E@`6���u���X�r��rj� }Y����x�@؞h��!H�~�E�B�rP�'����2GI"�d��^�%�@[>d� ��J������{hdP$MgW�]��\:4@��T[��~�b!6��aGtN'J��	�۴���%��I�%6h�5A4��$�+X�9�QpPm�����U#r�މ�F�,��R�����7
ֲ,�tɨ�!���D���oL礧9���bH��
�	�ɧ�4T�U%���5�Sj���R�u �W(t:�@�C�JZں@WS�,�4�#�?���͚�#L'v.���knJi��
!�oM��_��{>6�R��!<��2��X�Eƿ2��'�>>���yN������ԉ�]I�t�����KoVӣ�^vLhMWz-��UH�I,9��̤�����!Ń���	&{�0�9��!_D��}��PF����_5u�a���d���x�+�p6]
��}}�Is9��d{1]g��V�J�/���Ǥ`���w閒�e�Ek��Wz���z��gb{�H�*OŴ���1��vJZz����
� S���!ڍ-��ǉ�р]y�����Dm��C�,#��+ۙ���i�2�1X�VJX�����{�����P��糹���?DoϾ���1/ra�bg���C�g���2�/[2��,�;(��&������J�H?���rkM�(o�[47+켞ڵ3�)��V�2�U���J5J��N��^8Q��%�:J���O��Մ�IY�@Z�: %-B�/�u&�i���\�ީ�»��;���Y�\�/�9�?��D�c�Z��/~�?��u��D��cW&�+�Zƕ_;x����'�iؔ�:�4W�E�O�R�q��\7�wyw��Ξ�Le�X�8��j_8�Ua�{c���J)b�4?z���3d4������|�p+${Ea���EUj�'O83����:�ۮ����ړ����hb�J��S�ŀ���*��ӽ��J������K�9�Wt���z�X��OZ��G��=�
��:�{K�P���䌪j؈�Y�K�z����?C��N}�����g92���qX)�KG�x�]}��K�\����f۝�y�vɟl�{��OS��H/�r:�r�Ujmq�Ue�B�4p7G5�r9�Mh�|�Iw���n���,�6gn�V�/E��i��Ѣ�E�4�r�*c����t(�V����{�=�;�'�"��!�u��Ţ�Ұ.Q�b��
������.����ϋ�K�����1�^z(5#�~町�N��.�	�NY:`V1�@Ph[�wZ���#��s�H{t:�/�2qk�$�_(;4J���n�.瀢���N��n�	��leX/sz"��+�X�ص']���~�8����.{�����y��h���v���7�����C�v"�S��>�Y�	K\��W��=��{�EfI�4�ߚ[�$S����7���*N[\�)t��T�+O�HTFF����/ �7+�%�?��e�C�<Y{M䙜*�$���'I@�V-�d@�L�5k�W�>��x�{��.�e��c3о=H�ܧI��r��j�
��/3{���!����w�P_ԋ���2uu�$���i�&�����n��[e�R�Ō�?FA�>����E��I}�_iaG���|�����x�>�����ll�d�A>�W���_^C�a�T�F`�B̷�eL�6R3�\feE��M!`��[Xh�A�k�%�]�P7E�l��s��КS�V�vr�U��0���F'��V,�v����^]b�=o�
�ܺ�H�>j�j�ֿT8ͩgzm9�ӄP��@1hBr��9�����+7x���k��f�?��() �i}g������d�=B��d�1T-LHi:kF����?�ȍ&>�$����Z)�f�WĢ�a�`�c#�R,��������p�U苗SKU��2Gge���D�r�Uڬ+��OƘ}�K|���͡�\ڑ���S|���I�ہd@x+�ޣ��l�vo̵VQ�eߚ��"*@�dӌ�ҕ�8�#d��Aۿf�ʳ����{�����<���:�5�9��X���l!���p�R�lC �0��QB]#��8]�P?v��7$�[t|T-��@�{�;~�B��ur$얒�Uo ���&&���I^ȅ ���!�A�K�>pK~nf��X��UN������ ����o�(�u�*�wH�$���V���OA�6D�EeR�D��L��ER9�o�wOu�F�%0��\kf����^a��/g�3��T�g�`29-Þ�.��p������^��5�k��j�.�03���Dz��/K���4`9��Ӟg���#��s�k6��aT �ɞ�A��|ð2lz�k�]in"U���c��M�<|���Dd�U��5��.�>�n�e��@N�wf�w|�D������LÃ�=jz�ɚ�
�Gs�8ZY��4>b���h;�}iH��?�>�/�Y<|���q��e�Bhe�Lf��8z��|莞�@ x-A6d�G�kPwypm�*r7��t���f���x��9�����>�@��IRj1�6@>��=� ���8�W|@W��vo<�Gt�)��#W�e���崖#���zy'�[l��*V�a����ٖ��-EtkKJ�p�xR�Q/�����u=�S��Bp���V���(p���V�&�*�_*  ӷ>?Vrt�Ӛ?dN��L�и4�������hR����6��	��j@�$��Y�_�ˡ-��p��z�yO��m� � i��`#�m�P��@���y6���Kk3\Ġ5~�	H�<��ؗk@X���Yvn�c>qcJ�����c�y���{)'}��з�txx�A��O���4W�h�:ڹ, �E���~&�DLE9�rYS�8h��&m��5N��d+�����V�=�|��E�̮��1T��͈��!ە�9�8.CLR�Ł% �˅�%������,/=!���8/�o�X��X�I��5�yO�g+*����d��뿮�	����_�ى_���ۋ�3����2��j��n�[iX�F����8�O��J�������`���	�P���fZZ�)l��3i���^�(g���c"0s��Y��<3M�#&1�z�
T�0 �%$�9�s�r��]�QȶN|\k��?42]� �*�@˜�4]��m�g�ɕR�Y��X.-h0���	7�5��|�ܷm@��(�=��è!P~��1��―Үl�!��V��pA0�Q��%�E��S�K`'�f�N��0[nÒ���"q�8ݯ[�������X����@��M�\2����lq���e�Q7(�i|�`�'�m2�eM��X`��o��-�dl��G���X�'���S4��oEN��B�+NW�!IV��F`Zق��K��:�6��������i�Ң�q�n�(������6L�j�|ف#�]�x�dl6b�u���<p�y��^%< @�(���-�	���Γp�F���/M�#��M���W�.s�v��/�DX����0X樯ԃ�S��L��W2:�+��c2G�zE#�����c�l��a�/J���dD��-� d�B�8��ޠ��`1��@�w��N�>�_�@JE���ע��Ĉr,�MS�	zM-����i���%����ߜ�J4��;錸�C����v	ZC�j�-������ؓ\���6G���v�R�a�;CV_u�2��uU_�Ey�1;�8�2��QH�̚����g���1Z����TGb���ck��˰$/��X�B�U�0Ád%���-XX</}F����k�>F-�dHP����ޥ�<���XQO�B�uegңy�A�uf̾ר��G(T#��LJ��#�~!���-�Ug��c��6��U��b�����BE=�#e PdR^���DxE	j���B�v��0�}�r�!$��ƍ� �G��ˈ���i�&��g�c�ң6]Zw�X-cC�1*)$�]HL��
�r��bG�.���r1�S�H.V0�5g�:��x�G+���X�HlB &Y𳞚��.BB���O3�轖�f��ᩋ��L09B֙=�9!��~pȢ� 9���jk1hNV0x�d�=Y�����W�0Ճ�G闁�.�>�I�M�@�$뜘�,l�Y�)ϭ��:�U���w�=8|�Ɂ�i~��쩪����8���\��pc��-�/�9�����?#N�&F<�l�ִdXt�g�0ė��S�JI=%�]\h�U�����s��T��̦�Z�`�ff)^X���.�*�[8��A$tjJQ�>�g٩* ������Y�&<�}�@2�%�t�Ep 9����##���\K��O��2OG�S����r��&Mc#R|QvU�:�J9�%��@0G��ȃcB���0W&��n�s�v^6���_���-A{�E���^��W����g�g�LWg�4�#�! �t2+���>mZ�ۓ����ū����E�^H\ֈ���u4��)B����J�*���ѝF�Q��� ҩ0.7~@� b�����<��8ؒ��j��"�㦪�/�)��o�����m�����{���0�Q��"4��oT��أ��h��jd�Q<�Vjtx�'��0�U�y#'&jX���;͝n?i�� �J��f6jE1=���Q&�ęhqс&%�}�ۍG�}zc;ty��n�� ���1):��*m���Vr^��+L{���m~�Y�b��Q]�uRzOe-jx{Y�5���䞖�G�z������>�z�%�Ư4: ���9��i��� ^&~�Q�ىv���]�k��[��<'c�zj�I��Q�&|���.������P���D�x�9��c�z�{���7!Ӆ��+B�|,<��G�-l��HfX���]��h�2�f�l��9C	_DJ�2�I��[�.���,���y6������v�X�C�Y!��ѐa���g,�ߩ,�&,41�ܕc�%�*P{;��!�U���H�����<�^vd��(%���$!]U[X�d�e����W�mf�yS�0#�ת�B߀ӑb�U�v,���@���.�&w��e������wn�a���7Xř���w\��q$�ٗ^.�ږ-+e�������m��ʵ)x$�q��HHP�~U�u|ɲ��ܿ���'���o4���B\��?�����\�"�a�&3|�"kc�e����\w�巚 �#�;
i!��(5@U�}G�{��j�Ϙ���$X�@�ߎ`������{��yb;��3���G�4��v�z�!���zv-��gDC�s�A�Aك��n���x�e/-�t��g��KHVK)_��k8�?G��N��	�6���Ppl��QN�`�n+���;AkC�ͺ�tCd��3�v�7 6Y�pD�5J������*���K�N���~_0���Ƥ!,�����"7b�5�m���/��&)6��]�)K�s9�^4�Qt�m�(,�R�@��s���yxq������������6��`�ǹ�F͵���k�qU�	M�/�#B��\!�4�c��(V�5��:�&�~��: �>�P�S�!ȖHQ`��ǵ���^]\��EE�/l�o�N�z�ՆרA�宰��r��Z��%�ȀG1�v�1���8�,ӄ�2���0���*��2	[�$� 9.s�%Hww�V�N4	�oG�����.@w�m�؀֗��#JB�ov<�Z@�m��j4�c�5f��g�b[�˃m&���*Ux��2������I�����A
��WH����z�!R/@�&N�EA��������F9U^�8A뜕������t�C���}ۏ�!YR������iG��x��Ils9�<j�\���C�#��Q��R�B�X�\{U�y��
[��cQ�?��iKs_Bɲ�����D��d8�{C��&���z���霣�8�p���З}}�W	Ro7���w!'�I{�in����+������v�Ple�i�u,��&GY��9�(��g�Z�B�_]ҳ�Bst�o�6���W.�g��˦
�ɓvc�T+S�hӼ�`> F�ټ�mv���8qO��"�;nL{+U�l�6WT��bY���`"�BG䙄+�ė�f袱�U(J�0��Ȫ�L���g4�w#����=3�bx�z�0J�q˦z`R�#$����׺T��$�A9�����dP�dʟa�wt��^��UvK���{cH�k>�Y\W�v��_���,��;�u�a>lǍ�e�o"�����G@��xSX�����b��RX�T�w��̬)�S�����O�Lk*3NaQ��8q&�Ι�b�K���Π�-iF�`"���}��>C����.��Ҕ�:����u��b.L&�m�@�Q�j��e��*_�C�D�]M1A��ٺgs��ˋ�d�xR�hi�'Mc::��+���J{H'�ɽ�����I��}1���*N����yǬ���y4b֎��:/p�}��\O��J�z�mJ2��ʸn��ʨ����D=�F�<m�1h?{����s����=��,)	�%t9�:h��gBM$0X"�u���K(�#o�I��3H��7�K��l7�D�xD����!q�?^H�N9H�)EG��Όt�>�b� ��ZF'��U��1�y�"�l;��	�)������H�H��4��xS���؍��Vl6�^/ȭN���<_��չ/��_^V#}���h֖�~�,&к��C��
�����PFo���+|r�ɗ� ��T8���X�����,kn>i�	5O�YIWk倘`x�\S=�&c�y�� B��_�h솹���K�H�~�}���j��~Z�"^ӠO����Y�����nt�v�L6|bU��2���Դ����致��p�-�9��zz2)�/��3vQ�[]��7y��N{S�uZ?��+�+���{����!�Л����=�%��H��"��r�Mj�ʀi����fӿ�g�Jp�����A�\�H����8�&����$aU��s�QH�4Ń7�i���QcZKR�J�v7�3�w�4N2�G���;� ޏ��{-����HmGW���2i,�w�	��+a�a{�2����GR�]�]���K<vvt�;�_�l�IU���.t���i��r̈�i���H�˅��F�����	N	ftH1D�h]`Fe���ć`�+�	������`��Б��T�h`��H��G��+��#,)� }6��ƕtۼ��H `=_���w'i��-Yq��]����b"5��W�k�b�o������ohq���8�:!b���Fj-&3��3��X~��#J0+[��uí�17)rA:�����M��h�=}:FR�1��&����{S�/��H3*(�Vx��O��c��Tn�P������\���X����ze�4lŶ�|����y�1K�n*z�2�?����MEy��H5�C�NC��g"�k�O�"Qʇ?�&�rƉu�n�Ϣ}ȶ�0z{j~>��K���Tf`_a�(+��⊞M�s��P����xr��k/������B��[�놞
9~��:�3}�>rFUg6y�K�Y�a/!�u�{�Z�7k�k����}���g���*�t��H���|%���q�XL���.3$������R��u�!��~x�jk�Za;�!B��>�
�R�5Xt�m|Bt-��8e���m�l[�nQb�E�#r�+��-�����	�V�ܵ�O-���"������1C�>p-�܎4�m�ӹ�4?eL��Q��������a��a=]�"D��sX� ����p۩;�T�,����MI/m,�����߷ھQ|�+|�C*AB؛�	{��7�uj��}֞�E���K���9�|��{�ҟh��&z,���׹M�"嚚G%「wU%�j�j����<�*{��2�e�g�7���b�
��Q���Ry��˻=�'rIP�����N\΃�N
*�?���$L�.�EN���y$��IZ�Y\������p:�]=��r
R�U�ϛ�w��}���A��R�C�~8��u��(���o�D�$�;〕B#�؎�W�/�h��o�����]{g��8H�(	��gS���=��Ϲ@�G.�+��S7��^z�\)��e�
.��"9�X/J��v(�_���C�(���Zp����N����6������yc�Ĺ�hJ������EF{}b�3`ֈ��P�A���W/|[���f^�&��r����
obZ��Q�0�����zh�BP�Y܂��J�2k<Ayf6�ʀ�,��~3TD�w��
�6xV�e�W��d�x!?��g����ǆ8��^���~w�t��YB?�ݧ6�c�M�$��F��n���ao�զ:I,��sM��MJf6p�A�~��k���
E�S���1�l�=�W]6�~fh'�v�X@�UF~�5C?SV�+����Q�����6���ݨ3��'v�Ru���U��G6]~���=q�,%-��o��>����R�ܸ����g+��}w�P��j��),��wr���9�/��&��a����ȡZH��:�F����%V��8�<�v#Q�a���N���5��&8'���S��5�}f�)([[�ù0��X�Y�«xj<N���k��:<(��H�o�GF��ɮ���JaVÝos���J�����뺘FA�(J�/r
���f��~۪�o��;{�p}�a��� �r��.2[�ٍ���	<T/f�j[�B�ap�rr����V��Ȑ�ʛ���MGT�Y+�L���7Ǵ�e�b�3��I/+�G�?Dv�Uj�ڤa[�kxsJ��s��΢?n�l�w�w�Z3�rv��f��T�䛱�|݉OȼaU@��Rg�~��}]3�F.*���c�F�p9D}��b���%�"����Lz~�X�6��>�/B^hc�oF�E@H5	D4�0I�q�볺����q��[אeOr��(�.�I�2�88�A�)�8��������{z�
]��`7�9Wk�B��	ׂ�Fk��e')�e��7�ü"�T��EG��3��9=�3�q�  R.��@�wm�JDqB�&巆�����p����\-�|������wR6�" ��da�����zt�MZ��ϳ)�O��ӝT~.��;%����〪��B�əR�@�/�0��ބ��H8{�)������ғh=zW���l,Y,��S΀�	��gk ��`u��Nu
.���<ɵ	ڰ�׬6��d�"t�o�&1�N�^��1�)VD�i<z4��Ҋ՝�C(�� t:;���_ɱ-�6�m5LoZR���VD.[E���XX�`6��g���(l�'"b4��]�~z:L	$<��~��;�s��D<�H^p{��tY���VE�D���!���Q,��8bd�_�}@�e��k+̲/q�$|N�y��C����4�D����K �]P��y�Y6�}�[�x�a�˭?���e������f�A��?���*qQ���Ǭ�R����#�k�9��2:�~���t�η\��Y˛#ǤL�(M����5;D+����Nㆷ�	���储�XQ�A�q�y�E��Ƽ��](X����c�M!�l���.Q�B����/�2����2���ӣZ�'φc�-p�w��\�R F� .��j��֖}Vݼ���t�s�X&-�](��ԫ���X��0e�XK��H�=�z�mHHL�2��5�MGz �L�5ĥ S(#� Y������u���'� �^��Z��0S�w�1��
ds�l��5���/��rw��X�-���oE�h���7���jh��Po#�@愄��� ��D����ṭ�	^��k����������8/���Y�9z{jU(}7����K��v�q�M�4�K3t��A�}�_��ӭ�)�	u�Ў��N_�*�CR���&��:H�R��%Z#*�/�ނ������C�"3���6�<�I.��w�%h��j���l,�s1t࿶
�!E�X%Y�T9��V7�)�5��J_1��.	>���=����h�|��+gi��.5�m�$����&�!W�MVW4��������&�tq��]�,��A��R�1���1���9�
r^�X�*��
f��x�?�`ݴ_���#��Иp�����n~G2Z�L�������M��R���+�Z✔ǾbC�8�[�}���I	��$P8d��*��	�xT��ڡx}�?}�E��{���`I50��w����s|��X��>໰�:Dm7�ׅ1Y���,��ߏ.�?(TZgM;:v$�c�)�0pg�ڪ��'��[�l��A)wu+���XOe���7%��9s��<����S?�3�|�9�ΰ�����p�C!\qI�L�(Zӽ���K��.ב¾�x9��lDu����:��R�+�\������QŦ����鍄A������6;�!X�>lf)�$囅���xR�y汰�9�="`Q,)۷.��s��W�vRh5T2�"�
n�?�����>^% �ifw�xڝ�ݝChʳvu)���K5�-�q�$���	UƓ8� ����S<�g��ɪ��A`xJIF_����`��l�S*ք쑴M���`S��VĐ'�ǎ�4�5�'�6Y����b�د�z٪���s?�騕R��QL�6����EO	q��R�8�ԯ����w ˄[����7P�G�=�����V:�:o�����m��bzL�Z�6TT^�#��M��S(�(���������nk?fY:��a_a�eA�r���g9�@~[j�g���M[|����-K��R�ח��蘛���jUr�S����O����ʚM�}O��&��	=�R+'���V�lyw�	f{M��l*7�c3o,O��}R��2HJ�@��C��Z�`�����5����R4i�<�7I, vLc^�<�g_ g�l�$�D4�Z���Vo��ģ�hD��.V�ߗ�l�Y�Î��3������.C-�|��m/���fY���^S��2ᷛ�o�p�˂�A]�I���B%A�G!&zAx�bWd�ҽ�=������E=B-K���UY1������<��3�vOW8�7nmZ�׆� �5X"�U��gB���X�5Է\��9�R�w�V�z!�����-)�R�}l<wn-�*.��!�ϗh
^����4������s����AL�>�OƮ��Js���1a4���>�ۄ��O*�;5E���+����\��	���L	k���%-�Y
"xW�ط"+>�R0.��9:	H&޾;sV{��ƽ���Q^�O���3V�����~�{_1ݹ'<�!��JI��N���6�&��-"�L��#}[��Ҭ�/N��YgX�eDS���+������r�����MRT^�u��ޑ���
����c�p`{�x5�c7�!AKp�(��}��61Q�/͙<����o���K��G%5�<-()܏\l�,�� �Y�U���Q��;y��p���8���j��P�IebcϹ=���^��fu'��B&[*˞��8�c&��ǕpHi�ȸ�D����-l�Qc�x�7r���n7������>os�<е�?/�0�����Q���tP��M�葑ƣP~�Ge�fOm�Q�,&�h˭��q��,�D�HtKfp뿆��C�?V�$�&Zrw�F�ð�*�/*�Ϛc��E��#�9V�~~g\��+7�iQw(������#*(z:>Z|_��p���L<��
(9��']o�Hǡ\�2Ց���d8�ݙ���Lda&���cw�uL�M�,�4m7�ȵ��������:퓺��'� ��ء6Sne�6��P�A�V���>U
�j����r��YN�ZFT���c;��[uz�v�r��.������#�� ��sh��Z��T!~�lK�cތ�!��!�  ����w+2Rf�����o\T�U���xFy�ڑ��nu?^� i�~Ц6����n�좓7Xn`?ԡ�<x
��!]���3����O�Pk���Չ��WmN(a�p Vѵ���~|�ݱ��Z�Wp�Dl����I`�%JU�9 'j�4A
�� ��uO0�r�59�w��n��Bx�@����t)�v�BF��<����n^�W�8ǭz�^Ú��h"`�f�D��.\d���9j�a<'�6آ��Q{r�G�{S�)ix�:ȫ��źD'���J����m��6�QYy
�:���@�)�2XB���d��`���gB���`��7�ó�Ud���@DH:��G}d�$UY�#:֒H��F���'�5HM�n�����%%�RC)b�ıo��u�9}~e`&�	�uf[l�O�$W}{��@iSe"%hO��5�IG��W���txv���^=ʄ�O���1*=A�/&�{��e�n��v���5 ��N�v2e&��W�a��^ ���
'L*�3|92�Gǹp���J͋.��F�0�_� �
��.p�ƅ�G	k]X��h|�r�_�y�@����L��poq����T�//?���i|���`~e�����17q�5��#���9P|?��t���I���,�G���E��ذM��*�@�ĜOM��=g���Q;����H�l������ �z�+qG2���+d!��'Ψ�av%o�6~Ƞ�75u�m����ہ����zH�H[r��@~Z
n��ƥmjr��a6eu��
����g�Bi�2l����=��c_ [�}�U����y�SG���WlT�g�� ���ƞ�r�~;�*���J�+���,�y�[
�ЧN�K�lyY��sO_ ��}����J��s��k�T*�6δ�z2�4�Cb��5É��N^L1G���͟���#���ġ��X/d�UM��`餣9�^�l���k
D�
�;M%����~΀9��)<�-*�~�RtS�x��F�Q�g���JMf���0�,�Ԗ�(��y�L*�Ih��^Z�>~�7춈�8*O\�30�D����p�01�r-��
���2���@�b��X�eW'����w�Y�=�2M��T��|xS'�m V[j@+��2`��4��g�IT�Z#�(�SM��B������0$�7�6i�|��ޜ5%��J9�*�<N��9d<-pK��\��"�c�\������ )ʈo���u#m�h$�&��#�Q$#��^0N�Ӂn9s�Gdp����Z����-��fwC��ų�,ӷ��mejv'�ƣV�o�ݜDq�4��g��?�P.���|B���� dk�t����ml�����n3a~���of"c����]�դ�_z�m
�F;�y%0�5S�22Ѭ����	��^���hn�n�� |����K����p�.@�\l`��M)�X}:w-�PɛÁ 3Y�	|cì�����A� Ӑi�ƨn.�!U���$6TZ4�z⏶o(N_����)������ك���F�j��A]o�Š��G�i��!Ԫ��|��|f>h�`����ny��Ab}�D�~�fd5� ���Q���Z��-.��F��,�Rђ��\�e�ce�����9Sޞy�t/��&�d��:�����㡼�E�����u�E_�g�O�v�y�t�:BI��>�2ʍe+Ǯ������5���0|#�Z��Yj31O}R+iJ�3K�=,آ0O�;�9`��9T7�׮ [9��'�,Sǡ��ܞ��C�N����c�^�%��dȞ�Rt26,�E������q� ��~�J�?�MSN>\��ކ\h��z;'SOӞ;91��t��D�Q�����HQN�;�Q�f`RW��p�4�����1���������8U��� `�o�R]Lo�����2"� 1��`���Q�.U�`+��'̕j#7Ҝ� ��|����s͕�"wG��_�5�j}ķӔ�����ܣ��wp��גOǟZ��,��p�Zpz��	"�\%F�$�Ö��K:��v]"=ڞ�s� �m��z�����{�Y���6W�
�Z L�*t���V�4b#R�l���ƙY�6a�@�$�G#,��P�@�U��D��R��~���a�+�\�+�+v�?����#��ap
�Q$�?�ͽ�(چ��[�	
�%O �W��k�k��ĮSl�r�8�N)+���B��ֿD�[� �G�����O�ê`��.R�:j�!'�,�j�ضq�~4~{�ސ撼�mH���}�bў7n���TN;r3����X�nT�vx��k��h�@�������I�}(/d`���0"e���'�h�Ci��/��j��9�A�Y_}��3{�z��X�.^��l���6����j��mS=��@�q\��lk�bk�s[N��p������Zs�g�@n5�܁sKD���M�$����}N�܋��&X��aL��,l�_��?���a�{*yoN�s���CZL������n��@��v��Vc��۱'S���P����@���C�����a#�5�l������qy׏{V)�������5N'�~�ș�³sz�d�p-����a�_2,gD�xA��(���'��'vrP�-e&��G��l��t�P��j~-Ic���r�G�1�W�%w�@�%u�^K�	��w�@U*@�o�	���M`���[�2�vn"�;@��$^��A�^��5K���~��N8�0h=��*��;�r���K��-�bT@�<[��u�#��'ߧ���o4�i*6��yH����ط�NS����WQ)����1A�P�i��W�-%�u ӷ*���(��g��}9�d�'��Q<:�$�XSp���������6d=�%P��(��|�
M�)�N	�X��c����W�Ɗ�`���[��4Zi	�5��ǔ��l�#���B�?��wu�\���/E+AB�E��y���y�T�o 0��_����ӭ'
Q}+;L�;4Dל���WL�qwڨ6�I�U�5�&�Ԗ��m��3�M��Y���+�Qi�,__�G�[5��X{̱m��{���ͷB6>v8mA_&>�Yh�&d�7�[�"J������O�������y�${��	�g�Kd2\���1AXq�+�	M���^�zѬ<�zHZQ��8=�1��I��tX�v���Z�A�2�������+amB"�ƱE/����ߒ�`���͈��1�*%$���ؖ͌��l�����;v>e���]C0���dl��[�w�c$*/ܡ\b]�L*��B��I��K���A�K��%�1���j�	%�Ѽ}� �D�;:_��Nf\%���h��,�W� Z�?�J�xp�h��Z�1;u��B���rp�������!`}�a����O�Q��k�ۃe�H�ʣ��
��~�����E�"I-P���X'gB�Wlfeu;���<�Z׍��b�[�M>*�Zp ^�3{�6���C��_�����J�5���`,�;3�WC����3l��5O���H��"�ù�a
D��$݌�<Q�uf+
�p]�k܋�`P�Ht���Y���	M1�bv�,f�{�L{�`1ׄC���������Q�):�S:��2����=�D:��}O(�U�da�j�|�D5�zm�q-~o�jLG�w���j��c��0��F�t�Y�-�n���}��Ƕe�K@�����-l�&7����6=��|���
�w�?�PIt�-b��"hчH&j�؛� <ra�^�Ý]K��2C�%��iJ|��Z��ף��+Y���@s�/��jy��t�C�X�s�/� ���~����!� ?�B��Vڿ�`5�>����>a��cx񄓑�Ϝ��3�3�PsH|�2;�ww����)'�����{�^��t�g�ݻd멷��$�#�ml��`�ա;����s�bt{RdG�jp-��� ��b��;�~OG��D<��xv�k�l��Dgt&���UM=R�V %���J�zcE��h�Ba����s�2���z�OBi\��xF� >e8_�����bF��N����g�y2ZCB�iN	��c���n�C$Њ%�Ǐ�\�u�������U�����l�����^6h�̷A�|���e��$��y�@U��󮵠[�+ɹT�E%�Q�G}��e��u`�n.(��v� ~-��+��Ŕ��LC�|����-[U���NE(�վ��ݧ-�M�{�M�t�؈���4�}�m�+7 #
���bX���1doʝ `Z���Z��ͱJjqLd{��e/ �}�F|�o��.����Pě�ωo��T��3�Wfm���<���^%{'X�Jҍ�]%kiYi�H�4���`GU��:xA�N�ܥ;+�fg��㓰5�B�D�����1�4jM�¨"���B�wK,RG���	�0��y��@+U8q��7K�^� ��X̏�єl?�<h�����n��=*[�:�O貚,��&�7i"�x2><�}�#����������Zθ�(œ�hf�rjL���t��o�g�4�)3�����\�ط"(�̶���ƚ��*�m�w��$���`np�6޺T�Ḱ�~������wO"�8_��˟1�gb;�md�^2l�ȅ��e�����h�j��`���Q[g�	��[z����*P�.8˲1�{�[`��,u��ޓl{�7��3���;?�C�7Y��R]��z�C���j�ٌ8��p}\���q�4�i�y����㡊x��2��&K�bc����н	]�ˌ6%�d8�G���ʬ=]��{Fof:zR��>U4y���sS`V w��݁��?W������-C�J���xW�v�����tP��ҠGdT���&{a/��O^�㜕��ޒ��n�9!]Ɖ]�8S	%����9b�����������Mzm�{����|xU�)-5�Q�&&�*����H^���fkJ~��:O��(-qO��_�+�}�Q������sq፟9�5������g;��t�ԝq�u��b섚�ر��Ϋ�C��h/q ���&�-3L�������|�UKz��d�)���c���k���m�Q�<;���-��f}
��3N";���]�͞�}����~�Ȟ�u���h��s��aD	�kL:0x[L^Ż�¤~,ɜ��L�B���Ub�k��la��E8pf�W����`����i�?A�ǝ�N�H�3b�n�1�A�ϸ��!�+�wL�C��`2�qxr5=����§�d���$�`�R�h�.7[ކ`�&ƌ�yx;+�<(=�7����,	F4n�(�Tq�k3|/)�F��8��nA1u>��5`%��y�j��l� ^�fI���6���Ō�����@ЎJ84(�)Y��L .Z�T�G�4ik�b�E��
2����p"@��\/P ���z��[&���<�q��9_�0=c�܈)��xjB�.
&�TVT#��Nx��S��^�c"U�KX(�e�T��O�{vy�խ��d����R��v�#+���3*Ѐ�.	>�\T���acV��gK�څ�g�J�q̧�I�<�s��ߒ�-j?��-�2��[x,5N:��x��|�/ pP�����H\8��^)��?�լ(r��fJ��)N�>Mr�f^�($�����8��٬��u�fִ��O�az�T�l+Ǣl,';+i�D��1�f��.�����~ĳ�*��}L!$ıP.���T�0�̬of�V?�%,J���Ɇ@_:P��f�Y�w3N&�(���A�Z�z#�C=
��[��E|��y�@�*��f藄��J����6��n��S��X�]~�岄2�<��&&_?#�m�?���sn�{��ޟ�1p,*H�R�0X�&��}
�_����߻���!���Q�[��X�g�#
?�Z��u�f�����:p���w��/H����ѴӏŁ��%Z#j�1a�:���}栽&p���w����:u~rc�s8��u{N�O�NX�PKndiBY�	�p��Ε~�̅�3��C�������5?�W�}����d#��lϪE��
:���0xԳn�Q��)����*8��*���ñ��A5��-�?��F� ������Mu�a�١Cy��_����Z����N'J�4;���sy�-ad��un�=zA�v��E̯������1������AK�DU���⚝F�j?dμ �R2��'�Eb����\-�Z��Er'��v{�������n�=��T�O�{>5	�v�
�����X.{>��78�u���%��:Vin�݇��̘�,��b6��'t�v�?�s���:���W�E��#�*t@�� B�EݰO+'�4�?�m�R5H��^\C���<[SV����c"+�$َaB����hye9��� ;�c�^���Ԥ���0�Ղ{�Ug���-�1mo"9��"tz���=ի�f��=Mo�V���|��t�f���y;:Y%�ơet��n��V����L6�'I_���8��_��c#������=�L���`�q_��rO)�<�n�̦�����t�+YNhʦ�I��D݀��-n 7�"b�M�_ahz����O� f!qP�����qͺӶ��/MdYBe�y����e�!�q�p꧛����!e5��!�iن����x~��9�4�
�hq�UE��se8���(��g��©�o��c�����!sP���(t;�3X^?�{��s���E]M�`M`��ЪL�w�=��T��O��q��?�g�~LNm��Y�zl��E���qt�LP{-z����T�RۻOO��,-��i.���G��񍠧��M�\jz�[�Ȟr�^?dom��؟Yf�m�� l2�O!Rn 2d�*��XMڤ��A��+������ICr��ꔷ��'h���l_�|�ԏ��im`��T���H�W��č7
�������O���&9�I=�G�(����)��H�[�V�&��P#	���7�4����I5�\�}��L�Ԝ~��H%��LA��Ċ=j�榹V�ڜ;�B�)hi��*9��s�]�ߨD1��A(zA�ݑ�n* �7�"=��o�3��`��%�����	�!��_zt#zi�"9#��NL��#~��B�#��q	p�U�o����'<Gd��
��.QI���}�"�c��Z/��P�Twq�#����B��W����6`��e(Cl��ǅVzL][�4�Z׊jq1E�al<��yjY۰���2�z��yH�Q�[X�u���d��0�I���ڭI܈�W�S��d3^NTc$o�� �%�yz�ʠy�s{��fBLI,��SS��橉ءX��9� vS���Z�G��|w��d �T�����d�f�C�(��3��/D��'�/��9E�ir�_�5FˉC��Mq�6��z��r�i)?��#�����2�z�i��H��Հd�b9U<��;_��Wc��/�oA�o��e���n����e�0J9>�r�L�NA��f�T�k���}�fz�vڃv�Q]���Kb&����9�|������y��0�7��3q9N3�(�<{�l�ҝIVi�iF� @���, f2�,^�Q����f�lt�)GfZ|��o4������T�iҖ�:��9U�_��N�f�gU�uе��a
E㵁��D	e���b���\��Qj������r����U����F���ۧb�����U�kv��)�$�#칬y0�Hܠ9E}}!�T�J���3��JkF�H����k'n$�|�!>Y���i�n���"����f9��w��L��P�.X�v4�SSf�7�"dQ�
wԽ�"��@L�k����9Wc7�X�|�c*?��4���=;�;��]�%�g��]U�a΢���pp������oJ���.ߌ�lU�'�ئ������O��Gz��ѭ9&�
�]2�s����d�_ߵ8!�_�p�c�[_�)Z�a2�繀�M7-��g�s�@JE��U�����s����M�c,�#�Y�j�`'�R!宂 *�;��%�=���I5�y�����=q�GM�M�$�9t��$�Xr&򍃃ذ��GKh�R;�ԪIp�`�$	ih�x�8"t�":��]r4k Zj��o�N<�" 5L���2��:��	���u��@.,�S��42��h�x��z��{h�%4��uիW4¡Y�1�,����Y.E�Q�!rI�'+��c�m�9wTy�L����X���,Hr��C�H�aM�C'@�}�1��t�w-$��ɦ$��Ň�����f"l�cM�5Dk����ɥ�?}/�wfV�}$���B�V�)�UU�xߖ��[���C���jřyw��2$T�:�L%�6Bo$Kes30�N?;]���\@~$'�����"���j
t5������YĊɘ����j�:o�fk�t_뎼9v��Iy���d�<=!����bNQU�}� 1�*��'���j�I���@�]'K�/������|7#I*O܁,��I�������-��ZΗ>wH�x���u/c���!�m�0�v��}�~�¹ѿ, �v�T	d.j�Zr�0�����1Nƃg�
]���	m@�8&��[�W:p�hy'o���r���H��=С��\:G
m� �Huؠ���'����K���	�k#	=W��+rkxO�$S���!�_��R�T)/:R�-ӯg�6�3�O�Ԇ����@���V	�]ë���_j�c��]X� �����j����77O��� �|~Q�p��
s�E!���v���A�"D�'�W����WA�ዺr�^x��сƲ� ǝ��^��k&�ހ���L/K*�ny	,	鷟��.=��</U;�?�q0��z�L@�]��O# c�\��?�q��	�[����ǵD���듇Z� ����6(8���&���|+�|��RO���H6�KÙ�W� �_�&U��Q6��C֜�h,_r%˗��y��� �S�$q`2
7��+��K/�ä��iM�DF�Dw9c�A�D������
-���u��o��ǰ%�(�h���5�~��L��EH��`�ܰ`��u|�f<��{�?�e])��P9E��/�p��T% f4�EUN��B�rݞ|� ��]�����l��5��d[a��:�4t�6����n!�J��yd9�:`��q)}7,�R앮��D���`���O�m�����0�S�ǹ��}2AӞy��������%�j|�S�V����H��]b��GS]?�!(��Y���:�����)��a5~�W����Ƞ$' �qA�<���#*��UE󎇚g�K���@m${�G��� $������Y�7�C�RYT�j�A^��Ǐ��c[�@�g��%sCI�#N �MG�Tx	��W&�?B�nKf?a6�x��^��!~G�wr�5a�槜�doi���=$��3?\�	l��Od���:}�#���J�Oq���P�9^��_�~�8���Z��2Km�D�遨s��j�~��m8Y2�a��ᰐ�:�`\U�A�n}oى��uatO�;��5��!�Z7��2�%���sz�_He��	�G_"\���(О�ǡ�U��^�Y����_���!hQ��^��jU<������b�����-Zo�LF��߈0�<_�dx�Y�앨f�2o f���v`�ğ�2�-�S)�
Rb�~�eT��r@bF����^x����`;%+����=����n������H�U��T��slK�l	����mdG	]����]��;��x�T4A��
��$�{7�9R�>7uņ����-�����tQT-zf��T9��$���/9|��Sny�v���~�+�Ru*�"��e0?cu��@u��A�:�Cn�,ʒs{TJT$8�eU����W�;ZY@=5	}S���o֙��&�7<
�r��7�+i�?�&��c�Y�0QC�l,�c�ȍB���3���u��^-�U&�Vl��N����`�����U1���o �3�(:�`�U�#:�t���ǻ���?�_r#�v��ҡ��|
u��D �a��`��B2�V/ְg&�<���L+�����PSy=z}�3W�r�P}�0S\&�ud��W�����FD�vhX���C�n�-�V�Z�������\~#��ݽ7o��\�4�(?�$\�9�����i+ZN��`���Xi,���X���Vҝ4�J�!x'OTB����t��I/,oak5>���q��8�����=޳��e�2<����wi�
'��,�����/�£DA�3�;�����> �>�3M�"a�\n�Gb87Qd�[��͖X��=���c>�c�i�1^�9��T�P���H0��2�RՒ:I�Ig�k&���jX��}�0k}�����Ŏ9B�T��ᐷ���.%֟�ԩ�Z��9=�G!4��c7@aK��}nU�?:$|�\�������D���^��쁁�I@���c.gn��j`-�Z��k�:F-�{��>�Wd����U��n�+x/PӤ�\;m�[���D[��
�o���r�Ml�  ��Cp���8g�L7"W�����9D>�GL���n�u��-W#. #oKg0͏u��8����k��J�u�/8�0�e��h=�'�Y��\ރ4N:�Z\� �tJTaG��ю�|r�ix/�-o#-��r�������0�d�$ �Y�m�Ev�X˛�u���I����� �ӋuH��t\��_Q���-L|�L��WFJzB<�B]Iڲ@�6��w�;�`��)��������bB�L�5�&�B�|(�Ԡ4<�$�<�	��#4�+�W���m8����Ϣ������lb~l�,E��V�������{�r�颀S�����i1�$��A}��ls�e;{Qrӈ�#9�i�x���Z�}�*���Hl�`�{q�	�<;�sdT��S�~�u�}���5fO�x�H�eAӌK��t�%�	�.��T�����$SS��SRF7i:�I�.\G�~	� v_Qc������i;���r+���|��pL��Ǿ����']	�ޥu��#Z���\/N�>�����#ۋ����Z�t���0z��x���<�E`����A���,r����Z䦛�M��9����ߖ�y�c�!��V��k�۱+R��j�԰+��� 9��f
����TbZ5`���^6����Kl��&�,�E�+!�amqf��<�M=���W�S����E�e롓� ��7*�철�/a�RtMv��*P�T9��)�A�<T����=̏��ML<�"����\�'hz��5!����/\�.�Rs��q�S�.����n��rʎ-y�(>�|��9�(��� ��h.ϣh��J��A�m3-�?��h�37��[�ja�J��~�A�F��cۃ�#)E�u�-�Q�p\*���=,n
��^*Ĥe?�+)��`��~�YF�e:}�/F����n����CnL����O�)lxlx@�S`,`�T� �̾�F��I�6���Pˈ�w�~����ʾ�-Y+}�i�ꮊ��1���b�kt#%�P^��4"�,�`�X|�0���Ư����p�G���+�;x�?,h��Lr�9c!cP_s�\>�P���z.T«������Y�ͺ�y��&M�!�w[�w����ň}���nEk�� �c��j��(T��ty*F �ɒ�6뵁�*s=��u~:\�(���ֻ�����`7f�$���fV���� I�rԿ���.Ξ�&��\��P(~�8��(�>�,2�,�`{�c�;U����C\�����6i�W�b��N��KE��#��k�	�l�T�FH��T[��D��U�3� �v�z\�8�])�G��Q�8���V"m�����%��&|�m{��I�y�՗{ iM����U[���5U�����v�2bt��g��CL���$FQ�p�-^;<i�O�8лy�Ͻϧ�ok�����=@`��\^���U��C+y\�o<�8'<m�Ee=����K3��)�p��%.)���EAj�}��b'�s�U�gܣ�Wi{[N��N1?���=��6(; O�WK��G�������ni�Þ <_���Y^/�HB(�T�?����b��p����!Y�\ұw�{����W@��5M�S�����?����%��e�B8��3���LZ/�6����O{*H�2g0��'CM8|-��b����#��i؁b�@<+��0go�y6��f�Ԃlo�-sG�6$����Y��w�����JpOE=�ص����F�# F���G�DO��~��Ǥ�-8`Lae���/Yu�8Ȃ�Z/��!0uɆ�r�alV�(k�N��d�,@6�J�����f��^@����G��d[��FɺU�"�>�6	G Jq���.z=$�r���O���e�l�����