��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+�Ŭ<� �{�>U�%Yä��+��̇=��[�C�5a��R�����ҏ>�$��7{Bv0פ`E�
tơ��;�{�F�V5#1~�A�ե�2M�ڣ�o���GU�&��q*�t$�\�bsu���"�b���gۦ�QR��R�]|��־e�̢�?��@�Y{�S���O���Cnp�S�/��U?���yX�=E���R�$YU�H#4 ά�x�3"ZR-?�����=�!���\����q"��ípB��%K�\h9.A�QY�ŏ�	��u�w72��'��a��(?�i��aM��:�q��ؚ[}d�-OnI�`~��v�EhOt�UB��ʌ�5���V1}�0��wךy'�X0��7����oC�D�n��\7��Oْ�wA4�g��`�ג��Tzx�:/T����9��i�Ar� 1�5�s��U�W%�eb�ׁf�m�������#Pj��]��R=����{��L�=B	�s�r-���J���e ��+�6r2�܆��x�
�6�?5��O�J� )�W1�P%��>_��ͤ����@�*(mw( bF��=�
���ܧ��v�.���-%O57�UTK��;�Y��U�($cv�gF����A�};${N�u��o���j}"�S����J��v}��9��d{�K�UB6��]\��3ZSN2��&�#q���)�G s�p7��@UE�k�|h��ܛ�K�u�S�?C����0�x��y���rF�;)Yp>jk�s�P4h����8���3��(X]������9�%��sd؅>F�еl����3�a�gD������Rla-��e�ڜ�ٮ3�H��/Exx@�;%�*λ�Xw�4u<���T��w'�vbP�DŐ��:G�
�q�|D��h�`f82'h��0z��jS,�	��_Hָ8̋h��|߹?���|�ā�Ʌ�-8�Ҵ�;��m�P=��M��TM*o8�8����l�D��5��f����tW��˗Yh�2-�*J�wDoZ��_D��j�^�b�F�+��gOج���SMaY����H����H��oE��3?r`����cfkЙ�=���BU9	%u���"��;$N��wM�	����ݷ�'Kk*�q�"�_��A:����|eD���$�+�<[�-q��t��^��;fXd��T��>�'V���DU��zl���>�Y�F�j��I�T��n	�ligi|�z)�o�����J�����~>�3x7�{B��3���K4qH;��vs$]�ψ:�=r⫘�`�6�CT׋�鴊D'kP��^Y�F�������y�㑆:�@�F*�be��� ��ߍ�/��ڟ^�����V9qk�����Z�	%mlw��Ͳq{��I^�@���#z��<BX>F�B����-)�x,~J�5N�&ܧ����<����N��'�.CE
�����ZpN,�}��#�X%��S���	�Mo|�5�@���T轇5�{&
�]�\]�q��:Ք6��$��c(�A����X�~�B��,�%f��3;0��|s `EAn;��ih�f/U���p�R�S2�2��s�
Nu[�ɘ���*žz����v�+�T�u8�l�,��ұG��^w�WdY�	� �m��{JO
svsط����\x����'�6�<�[sHQ�iu/�?�x�?���5�;\ȯ���M`Jye����^t��ȿ��٠�h!���#�-�E�t85CrkǛ�� �N??���֝T*E�y�Z�/9��x:������.x��6�<����ǻ�F�\\�D��pk��|�7��MvζQ�� L��;ʠ�:̸�]aq�5EԱ�>,�rйZ�z��r�e�����h���!�{-[�H 1Q����0f�w"I�)7v�n��'��y ]�	t9ՠ��?Lj���Nx��쮷1��� e�Y+���|��[@4�譚����`9_�"ڗ&'Exy!v4�)�� O�p��&�+�nH�ܾ��}��Jh,]�~�O����urQ$�������%�'VZ6 �����M�W:Eri��i+S�C"�n��S��jL	��C�ˣP{�l߄�4�5����)�c]`6����S�*�R��JN���`�f66�W��+���n�[������R��ʤ���!�*g���߷�&��DZzm�o��@��Uq(ɘ��ǯ,sw$��k�m=��gܑ:삙�0g;�K��?�$�8u���,}����g��,�1zNlW��9%��=�g��턲����U!s��'��c齄R��9Nr#X��ړ��!����ē6_�� 'Jyң�Lڹ��9����k���#����Mڸ�%.������YX=A�x��y�JP�`Ќwn�0)�3���rY@g�����O2���>cz �V����x~z��8R]f�����jw D��AЙ<����k�[(rB+�c�����9=�ԭi�#���"@��.�A�6���S~yL�� WhL"=�X�D��W=SŘT��W��&2�}����[*�ڣ�#�3��eO�R}�+
T���C�b�]Y�T_�W/��0B��4oHd�	�0.-C�i��ɷ��h�#{�H �y'���y�rĆY���@WH�E��S	��ݯ;�R=%7̍Rv,�i�E�Y7�+��ô�X��䑶=�w��<�Pd֡��zg+- X6�q�4
�S�x������B�ސ��eeҞ`ꌇX���>JC���ƾ�c�%�Y���u���"/�B��l�E�G�"�;�>��d�Bوk�A]S;C'�VK?�Ǒ�g��δᵼ����j:�(r4K�3�7��������P/�C���,eA)]�K0rgk��j����"�X�#��M�Q���[(N��,���vB:39��:�V�Y��>����ق��Ufn!�>[L|�BO��?���Tzq�d{�M�+�����
� �"�WՏ��Q`�N�!ń��SP���9��%�GI�"�!_a���e�O���^�4ə���lʡӚ����΍GxW��������)�2�f�k���$�!2�G�P���r���R=/`/��ˤ��NS).v�3�f������,6=}h�gV�GS�g[u����䰺�V��,Bz�Cv����t��ju��uŧ�Fgu��A������u
�nK����i������f��0����,�����F��66�Ѷ�3���/�Ї@�1�חZ���-��C�ݍN�m?f�<