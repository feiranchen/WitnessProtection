��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\���=��sl�^��V����Y�D�?oqbN�H��/�u��;�oqS�\9����)j�Y��RZ�x�h����*Z�Ű4�_�E^�&�<fN���:j���p�"n3����V�P�T[A��'��*i��~LYWϚ1��ͅ��j�B1����/�0�Ή�b�0fς8�4|�A��UO��b��s11M �����-y���(�!R�j<S��*2'؞FSE�Կ�z�b���W�޸=.:x�B�k��=dL"p�e�C�
on���eD�'����:�*���y)�ؖ��(���(����n��O��Y`5k}NY$H�x�E_n�K�q �����<�F2q�aV�=�"�By�ƱbU�n	pI���E�a蜁u�>�)���=���G|�.Sa�R���,��U��DoJw=ZV�@�񹗔�K/ �)� ������i��pO��EG�öD,c�S�nB��r|�dl!�@�6�uw2�xLLW^8s��tf��[ڰ��hL��	���/����y2u��laC� hA���㓐9�=ٽ�t� pf	I� ���W�CY�M��/E�F�V���/?;�?�'�L�(��T���`����e.e�"���,�'�I���oԤo��k��@[r�����6L]X�Y|MA�6f���-Rm�&�qE���G��u��_� צ8�юtot��(�ItŇRD&B�����i�w���ID>?��kU�V�p��nޖ���m�N0��L8Ed����K�����_Q���H4�W�a�y#ܷ����U���i��!�k#����c_���W�����YS����?i��95�QWS=�lv&�˸J�`�� �A���R��}~���T���~HN���uOj5�o��)�?��x�����s^�`n�M�9����x?�z�Ж^��uO�k�G�7��B9�9t	�I$;�>�	�0��
L;銻��*�2x�/�`?���X	]�Y�H����
06�؜@�o>�=�~���+hk$`�3�.~X�Eg<����Y�Tq���/�����P@յ�P���,:����W� ��X;����JԖ����'����`n�k˝�"�O[��nt^
V@eNA��CpxQy�.��4R�|��j��'���'v>
䚧g�$cD���X�!o��@hp��YNt(Š1�6�'=�%��A(�����s� �Y��2ve�
�l	&�X�Խ���!���)�l��V���������(���g �= )~�p���J0襽�v�s��d��|��z�Xj�������M��:h춶<�8�2�4YM�������j�BHԖ�_Y*a��-�v��v�Nh\�H�y�v����&p�5�p�=>��a�L��h� ������x�^�5[��������=a���g~T}{@I����w7m׸@;"Ti�c�F�fN��w2eT�G7!	���M'�ih��tQ�F!z�����M�
�iZ��ޞ�l�[^Sk#R��
G1tw��%��� t|���ܲ����Q���`�С'է�����1��M4�>��f@U#��߭m IP�������o!�b]��og����h��"\Z�.`5������Yc���F�ZEy����c�~f�+F��x�r^td"���}�)U���l���<������ubL��I��@����]�"�o�fu�BJyc���-^Men$�w����d�u�D<��u��j�hrn*�%��	o�w8U{��g�}����%�hO�$;��7i.�Q�]�t~~�b��U�y���oܕ$>]E:��&`�}e�	z��Z(�NG.8,�a�Dr������V����:t�$`J+��x��IuRe���W.7;𵏛VW'��F�X� yX��*�b��>��R�ll1� �U[ᓺ3?���6*�s[�9�܆&V�-�`�?�[l���i��R���^f(J��[	��C�79�,��x��t�@o�����1	���=F�nc���G�0t�72]��/+J�:�t�z��dz
%|珞0(�]���3)�4(a�����EE�F�[W :����-24_`_���]��f+����緎@�BH]���?��E����݊���G�4mzb��%?�c::?p˞���ݕL�#�������àY$u��z�W'�I���%�p��=@l�9���[�h��	C1v�Y���@��+�/�\�G@��º�dgZ�c�Qh�n�dY�T`��=#Lϼ&��>�C���Ŋ�9}�S�5\��]c�[����<뀛��=]�v���Fdp�ۓ��U8j�`	�9����D�zZ�Z��b6oJXЮA��Ԧ<ҧ��E�q�mk�<����,�CM� �.���m�grJ�iN�N)��{Q� {]1�%<��OQl&��l�<Ä��l���=��o�+'�#"d�L�'�뫜�Ng8���C�:j�)S�nH~���;:n躶h��q3TX
�?tC��tK��>����ѐ�4�,���G�v/E�0I��m���Х"&3�VE�\���$��Y�?%�d�5ȶi��o�����^3��j-�e8���$�M��a:H(w�k��%"(���Ӄ��wJL2�&P}���9�P�L�	UR&����S���n(ASe>�D3��D��0�k.y:��%���I�����][_/�v���=�4.4o�o�0��.�G{]�gp�Z�]jS'iGO�N��K�"F�0r(���F�7^$��G+S���y�����$��+�����Zm��洠��,6���c6����n��k��k�c��ײ�T?�!�X"i�
�����bi���w��i�~v�]"EP��q��o�o�]n "I���xb1@���f^�]Sg�a~,Ū?��bln�.��'�D��= (w���� ��qZ���-�k1�슂�O���1ċ	S=&�B�2�w���3k7WY9�=ѰQ�g�_��/�#��rXJ�e�_���-�9���Օܢ,�`�ڧY����2Tre�f�ab��ꇢ�$�0|{d���}��K�j���XR���2#�$��*��5l���H�&P�;�B��T���%9oMU���'�Sf�G>�/?
�m\�G�\s���#0Ȑ0�]
J�K�.i$'�#,<
�' 5��r���п����F�����^��J��b�=�,�W5,+h��c���]���Kى����S�U���'I����U_bhF*@_�Ah�ر� ?�5]702���&��w�C{rx��>FG��rq8�q����������U)wR��j~,�cZ�hZqH�����E/�i�;`�""���Eԯ�$H5B�⦦R�����2䔭�b��*T��Sӏ�5�=eR�#Q♺�����)BB�)�(�c`'n�6;7���<0��ϴ�$y�L�@eOy��J%���L}�� '�ߢ���]�"W��$EI�b� ����-`<Z���چ��))`έ��F��89[��f&	��:��>{������>k^�;1�=���z��ͩ�3���^��F����e񕖥�!�f�"�Z�B1![I�;�I������M���JgeE�wj�2��ș��#Tv[X��Ll����|/z!t�ׯz"K�b����ȶ(tK�K�ڕ���z��:1$���w%��V|��E��F� BrpE,�@׺?��Y�*9��Rq�Z���uq�D��(�We��ꈈQ ��ho������*<�bc��dq�e#҆���E1=p�pS�m,)rq &�_8�:ߩ�
<�w��!�it��������ҟ$y�=v����ݹ*��үSD�������q�}XP��.M�0�k?����+T��Sr�♍r5]Z9����60̦�)0��O<��	��utꊯ'�3�}��x�2'�r\m�g���a��L��[�M���bͦ�.ݾ;��vN�qk?f�4Nt�	�
:^+�+����M}��<��~�$�U�=Ƿ�&f3�ց���$=���i�{���}i��w����Շ���p�ǡ�2(�5R��C᫢�ɛ�)/W*�Z��#[)��szUӛ@ܕ�-��C�<�����cIR�>�9��ACkTcdJ�]��z�i�gxo�^zKz��䲽�g�z�gQ�0=h� wL�˰�Ӈ�j4v-�ng�8V�қ�&��h鷇"��@�9�=�\W�U�z�6�*�!�cieڭ�ziDY6���)�f#_y��B���[�pV_>�5���8��j���V�{֢vP�\Z�.�2��zƵ��4��G�7g\����]��2�h'�!��Y�w��۲��=�v�Q�7�����X�z���Y��N�&@i�pN 22x�?K�G�N%�ÄІ���UvT:I���)ϑ	��A�RH/06 ����$�w���G&�F�+W�v����M�dy�C X*�aK̋�� թk�{J�U�,���O��e�U��_�]QD�a��G���|�k�Z'h�m��.+��Q���%|>��]E�	��gWW	V�j�\1Ռt��W�WX����l��F�r�}�j���8W]ƪ�,Ya*�"�ȬT�r��O��f�,���=B_S~���L�qK��o֖W�N��C��a���{z����������3�>�"Y�昽���*���Ǽ�%���h\�|����i�-H�)��d�,;�ߕ ק� ����w!�C�a���)7�7Y��-�(��E@���t���ǵ���p2Cs�CzI�]E��@�~']D���B!M!�nX���-^�o�&i��F�Q�&��	I��)���_&m�L�i 3��CN�'WW�-b����2[\1�s�	D'Wm�uX�?�.a^DI@�-[�`��:9�f�M^nE�N͇�U{Of�X��Xq�yz�Dj
-P6b3)ψ��:��0� �Uy{���f2�M�ߕ��	 q; ���S�{9��Z?�g��"��e���1�K�磁4��0��-���#U\K�޿_`������B�!�Ysf<d�a_ �4�q��̘���M���TH��)Pt��[}>��b�&b�L�����<�i5+�u�]�b����B����_=��ܙN�w6�+}Xn�@���m|�od�m���-�8�a(���5s+ѣ֩jW���}�4[MŴ��c� �X4`D��oaa$�?��i�F��&��t~�.Lnx���uwm��9��u�xr�E�o�(`��,�E��9��l��a{�]�˭����*��'K��=�E!��m�����՜S���΂�����Ʀ��c�ݠJW�&^�P��)y�4���SL�Z?V���Q:y����K]�D �Z^\��;@q�>^��������Ķ!�)�I����JD֑h�qF)6�&T��_VE!�@�r���Vk�,����`���<��P�Q]��k�n���1n�ێ��ڳk���3p�;<��}��µ[O��m�7��xZD�Գ�m�k;�����y�����#{�g�
K�`��Ns�jI_:ŗ�Ǥ8�zs늈�eh7�I���Ծ���3
�@�����UD��O�h���ֳ���X(�5��~h-�2[d�ͯ�I�����#�}�4���//dÜ�`ѩ�s�k"'��i,�"����~��M�d�/{h�o��0Oj��d[W�m�#S����?П?��br���(#���""��($4�8�3J'���$y�
 �N���0��Ih�JU���[�c/wݺ��M�Y����ù��Q	��C�S�|��	��r�)?U~`mV���(�a���H�	��R���X0�eu)�ɇ['@o^�T���7=�n��c���y��VHz�D�����
�0�����A�5��8��(-���Xb�]*�3��%�NZ8BV8A��7�.����ܫۻަ��7�4א6��+����*�fM������@��� h<�Vm=�b���Y��!�e����A?
tv��$#��b���_��솢��{h�)�ʉV��<N?���4@?�'(�o8��b���i����t�J�M�Yh�)N��)�fC�(C�e�?�oͽ�>&zDN��|;��/�D���{�Er�iFJ)��,����z��{~��i��>�}�a5S�����ޠ��|
�3s���aU?�FߑA�[��x#�$12��4���� |�L�|s���po:��%� + &g�ehd6��x�&�.�@�fZ�{Ad���E��l7��a�6�(��K�� �H�	�t��A.���	6���)���0m��pf$N������i#6vߢe��X����c��5Ġ��zj:����n��IY�\=j����� ��k�3���@2���r��_���÷�夭�_+AY��·�G�WXKE	(�n�dI�Q3�%�$�����a�D�A.:���2�޻�K���Njz@J]�'�W��/ ���N���k�� ��S����$C`,�{�F���n�&2��	7�%@Y�FR�3Ut�re����5#�)��y٧
���3TyU�^(���pߥh�LzT��2V�Au[rr��;H/q���A�C1!߹m}q�]�4׫r���d����E�:4���Y2nm�8HhI�Ӣ~b]�����ӟ���^�XM<q�F��f���֖;o�����X[q=F����J]�Ju��F�Ve�/����u�>�R3�xgzH���!�L��h�6khy����J�����y�JQ�b٧cOx�?`�QYh�,�Q�uH�MW:g�ŭ�/�3�J��Cy-�i���TqV���q ��R;�+%{b�@�Ia�$�sڴ�NS�1�5bk��0�S^���ףӎ�4�$r�T�UE���ɇ��
��\+;��M�E������e`�$)N��Uj��,ȡǂU;M�B�W:�|G� }Zl��ϒH��W���p�4�Ó}��}�q�$u��v��ۻ�ڗ y�֢��Z �j���C֚#��{SZ��p�\��H����m0R�F�V��:\�����k2��H�ԭRȖ ����H~��RU��!�P��!��k` j�Z{%���`NK�<V(��X7DiY��b�_ҟxY$,��H����pNN&G��8�/�Nѩ2mM��"�����`��S�ŘDr���[�vJtڇ@�8�*=Y�P��IıBمst#�J.;x� ��<n�s��ٵo@�ܛ2�i�Ӿ��.��.�>�ܝӚ�U��J���+c�`���aLV��{U�͕5��x|�&DwIb[c��	���a�v��>�>�-�WP�Ԍ�����1(x�(55�H�a;�TI���s���z���O���C�?��е��2$�'�U�1} *�[Lk��O�Du>�;������L;?L[�t�v��X���U)��`��.c�s�W��K�Y�'��s]�j�~�kQ���lm��L����!���������_��Zd2؞���/<2�{9՟>v�/��9`������M+���I�(�V���7�OXL 52�Q�.̺���~��
�����;�.~��p��w�� H.���4��<�/ez̘{�f
c �XL �+a����sĉt�b� �῍���2����+�ō�qĜ�O�~��j*�]�fR�&{{;�,�.3���4��U�U��\�xf�����9
tla��i�]̯'�5T-�������N��5���֌�^6��=j��&2��-Q�=���7�\l��Ť��~O��`�!f$
�#�g����,,�20�5�����f/�BT�P�M��,˰9��q��� !L��#��?�h+�_��1Ŷtn�����$ю����V�9�wm�X�T�e�O)1ٕN�6��
�;}�@؛�"�&�y��a7�4�aN�)!L�T����V��ϑ�q���_����f�Y�ڮU�	p%����}���N"����\��{���hjF��|d�e�_s|{�� ��h�ٸ.dZ���ј���Em�]����?�	��W��ܥ5��=W�5����0
u8*�G���߯xޱv^�yǳ�?��Aꄪ�k8���̣;0W�.����K��� �ߩ�i���]�雞ۦ��B��7�ǫ#�^K�� ٍ6��y����d��(��Զ�%.z���3�h5�?�Yq�����)�W����2����,�m�+H�s�8��Ch ��� 5��zv84�iV��ɑ3$�Ʀ�X�����3�ݸ?�51�
/�z���T�ub�k�p��x`����zG��^ހ�q+��BI�����|W�o�0����ƈ(OG���s</�'��x���K��Q� vٸӦ��!�����Y(K����3/=@.3��ʹL���t>�U��}zT�?A�}��R��
[�]��5H���JEC�ʏ�*�R�Uw̠:Մ�m�0X�K�?P*O3^Q��'Q�oJ,�AQ�Ԓ`�o��l݌�/מ�Ӂÿ���P�z��>�!o��@$��ja|A��ݐ��|}`��Qc�(�1��|��)F��}L�� �����qg��2Y�7n�U)����kݼ�
te_RXeA�nM�`��κ%��NN}G��΄"�Sc����C��v4J�{]2����Sev�� hDmL���,]�a�ѭ�'���S��?��|`h*e�� �3#�Ls�P:V.�
�ݝ�"�z�M#������ڔ�
��Ŕ.Ǎ0�B=f�Slt�7�!Q�$���I�?�*�R�(��>�^t�6c��51h�<��*q�9q�0Q�1UE;�<i2l�-��pML�oWx�}O�(,���g��xk'�xU�+����e�	�"x7��:���*�"�N@㐲J�o��Oq*UW�@�W�gɷ��M�%�c��yY��V/��]$�tɆ���ZoE��Wro���֨>�0��(�&y �Գ�d����[�2����@y�"�vE	Pْz�n@ٯ7�H]�Ym��X�C�?QzT�h�9!U't��؁�7{��~�~O�%��i����;����MI�0�W�����=�!o۞����=Hs�،t�9좖�]�嗅��z���q���MO���?���Y��(ZZ�&���9ҁ�CEx��f�>�#	
�!lE@���J�`x�e_��^Ox�	�`���� N�S��������Ts�P�=�V�
�<���w<iP�o��uHWSb��_��F1X�/R
R��<�^���	zC
��$2f���sO��j��\,zϱ�WU���V��!Hy7%V�	C�E��#�*F�����&w�%ͣ;q���%���¼�?S�k�J�!�B�&�U����������ƫ�&�tN9�^�B ;�oɗ'�5όv]zT��<F��^]���5�".��-c�R �������ynxz�f8%�B�}�½eAq��׳�b�T�K���)���vkJ����F�H��h}d��Aw��O# ���<h�z��\bEyo[Y��x��-��塉^α���*1�٠[�=��n�W�ZdB�|���x(X{\!�V6�	���l~�B��Z�����i��}�x����nSV����o4�50X�6"��绩��F64ƭx(�=�~����\l2&oJ��!�s��c�X����F�A3goļJYj�ں�C��&�Ԏ���y���W,� ��
&�<��:=H̫�F�=-#?�*����ؽ)NN:z7��=2d����>�!D��߶x�Ŵ5S�r4�O-}�a�6�U�,T��Y�i[؉=�AC[F�>
��v����N9�'D��I'>.�&��O���Q�3��F�0��7����Ogɇ�`�Ni�Y������$h����t�rt��	)9��$(�֤��+�+w��_��\�w�.��d�)MƊ�n��v�,��*��P����uM������2w�P lۊs�8����"O��XU7N���[%�����'_���l�i��,��.��b���[�u��@�9r��6/���FA�"ý��!e���/�Ng���[�r}l��|.E��t���m�vMK�g֣K�߫ ������H^S.	��=SI���.Z���x�3М�~޾wF�M@��ۺ��Xj� ,�8�0�Y�^Xdz���װ��\��6������e��iU�Ex[��&%�y������	�pc��@'Ü�;�/�6)�I��x�:m�F!����M�צ�(��;X:����Bu�,���k?���f�\\�-˥gk�|�(�y���*�
�&�h����UѶ�<������TKC$���Oޝ%��Z�.u3�C� ��\y��X6E��T�QF��L�?��U��!�vE}-CC�o;��M��&�@rKbJ�����@5�?���E!����D�$�&���NrU2eU�:O��=��q})��a����*!'}�L�R�ë�{Hn{ʨ���$��k��sG��Hl�ȜҜ�y_R��ظ(��	p�Ư<�}�Km����Rn_~��Q�0�,��1ȕ2�7��E�|��x��E���1(V酼�?�d�;�AA�H�(�����ƗD��E��L��V����m�������Sÿ{�J������6���N�[���g'x4v�������i�����Y~?��e�D������`��, ��c/�����`��!�?�47o����8A%�U��͈,K?Ɋ<JϮn��b�r� ?��v č� �v� ��N�}(# �>���Ӵ������H��P�]P�jS��4��^�)"���'�4���v���o��� �Kio�M*�Q
���H��^��Ƴh�*c�J��LKRWR �{g��BAS:���Q�%�T�[E�eӰt��|c��p;�⧝��N�N�����:�G�z�p	3� �� �)ހ����A�t�*�Ӽ�ȠUu#���y*<i�EG\����q��Ra�I�أ1gs\XTv󌍧�N)�����#`�J�z^X�N���c��lxUm��T����R�6��WN������ٯ�>?Wy��p��=��&���.�C޵��"y�5�4]�D�MZ��\�
�����p��k����f��#���oB�Aݣ`��m�����w�W��bg��ۙ?�h�� i29���
֙�?i�Ef���L�Z-�喿�N��hSr\x�x��P&)%B&�E�,��"r�ox����-b}
_z�
�ԃ�����.9�ɑ[&L����.�8v�=�-vmZq�_@j����Q8�b��Y���hNe�����U��� :���;Ue�lr.xL��^@��f��7��,@ѡ����<��g�˯%�^�vEI���3$��~t������C'�N{�r��K��X�k5��(ݸA��r�j�8jnf���6/�,}Nl]�"��R9�'^�T83p~g��RSlo��@_u���� ؾ}C3�C�dY���%�0
k� A�#�.ʟ�q/�R���*�sYqى
*/�[�5!�1�gnBf�f� �I7��ƥ���(�2ɽ\��Zj*oiMg��0��>�k�+d`%e���6kA���'l��B`�86J�o-����2â?e"8[ˬ2g�R��v4+p`� W��r99q��~��qX�T�B�����)L?s��	W-��#�zS�ߓ8����~P��2��!
S�ā� J~��w�a~��g���6V�<⺇j�u��/tt_�I'AC@qa�ٺ���[�ԯ���LL�w*%������[P�M�tÅ�A����U/+/f�E%W��!D��q�d% 5j�B�0aE��r�8�,�(�d~^"�pK�ucI;n/B�����	��8
=���}�JU>���9jXBr}"�w��r#9��ϑA�Y��Q��_ųK�~O�
 �j<�`��iA�F=8�yRgc�ٛ�k2=�~�xQ{&� ���8�~�D�-i���Ԅΰ,������b^�<h��2^`�o�_b]uG������~��H��=|fA`�-���8j�9+/&�����F*^U(i��
,#�Z���jF�	��F	���hSS~7s"V�"Μ�� F���X��nRL�L����!$N�h�z�,�̻�}T_��C���}�V��1Z�0Ë|t�#kk�7g(�c�q�"B�d�8������E]���RL���QiY6ڽ&���=g�(	Ԃ$�F� �o�ku���/
��6?�%OCFJ����f?ǙK5�k����kz���+3��rM\D�[�H��~L���� ��4�������}�����0��Ťm@�)����j��C]�3.�n�~��6jD�`���Z����)3��	^E���dn^�Z:��`7P�$�4�$����(�L{��]-]Ӱ�[�}dC�����x���lq|��^�QYq��{�u����)�S�表Ͼa�|x�%���%/�3���?*$0���qgR�,+��}�0Haf$����i���'H�S��&'r��#9�J3Ԑ�=
PB�������� �PZ?�ފ��ݗs����]�..�M�i�u�{��|T?#����j�����UW���Q/I	��L�Ջ��c�9[����+!g�ʖj���BI�V�aȡ1��S���w&�Ɇ�A�_U+j���^���_���b�A�ш��LI���=?В�}�(���ꢷ�:��̷L���<5��n8������q�:��#��F}���+�J�%�OOV��<�X���$�C1�4����0e������沎MI�r�E�P����1�i���^�`�N�Sp�r�t��t�F�x;�������c ������ŝ���GKt�:E]h��ә�"i6d9�+��"�j}*sv~$�L�I���W�]c�Cr�,�S�^����&ođh��?�d%1��	�|�K6�G����/����c�����!n�/����;l$̲h�L8wV�5{��e�I,H��y8]�a�͑}�Z��� ����z�*u��_76'��@�+­�C�����b5)�sA�Mɼ�-�6��n�?�}t~S�``zB�Tb������+߸�v-�ӯ\� �e�J�W��ɍ�������K��6_���9�#��5��NhHy�y6m@��|�ʃ���9W�%qĄ_J���JOc�5���8�9�u�ρ�?� ��Gf���1�������e~�n��h�o��5Q���1p�1�"	��մ	8^muoA�S��}����e ���S�|�=��*��:i�)n������v��=�/�<"S�kRTc����3,r?�MS����l"��Bۜ�� GEI�6VTBT�,^�;[w���D�=G�ĺѺ��[yC!�\��{���=��	�ǚ�i���`R�.� P�X�vi�L
=A�E�3x����͋� deW��s�8f)x2I�"d��!�c�i����K'�n{�(F#y撰�����йI2m�ˍ���2 =��g�_�5���@��<�Z̫���.+W��B(��̈́q>��M��IM @�Ke˕�\s��S=�hK�ʃ��G�Rb�w�U�*?��	_��1��qLp�0�N��
���H�i}f��!��Ђ9�u�L�H��2����(Wwv���z&̼:�7O��,�0������&���������vg6�K	&8����ʀ����z18�8=5|�y�g���U(oԓ)0�۬���z̜&6bG񔸐��4A0oK��_+o�8�	S�H<�����2{s��F�t;z�ɼ���G�]6�Y�3�k�\$)P�P��;����L`��������f�2uז)�6��J�yL��P����*���{�A���V�PȻ�����
�������A9Ҳ�)u{)�5�Q�B���v���^RC`�/$IJ=w�2m]�-��8h54�����AN�r�Jb�d��"j7a����jw�nM��.1[�Q|`w����n�	��t�wy ����*��az���B��RuH�$�{���D:���=�n�|����H�מ�F4j�ZB��?No�?o�a�#�ɬ	�7d],�.�s�F8uq�|��� �r?1p�2��9)nO�0˨��v�Edp��ۦXsw��R9񓤤��^;C|���_�#�/,���k�.�E�$k�K�Yx�ؙq��]��8��"������S8�aue��m^�d�T4��@H݅M��9�B�������p��ٰymS�X��u��
}���m��=_�:&l��éx_l�˙*�m3��~�;�X�_7�۪&��L�^.��ʐ���=tZ�.S� �qk��X�Zpm5Xa�Uܼɋ�
m;jo�?�q����a��2�[�q�E#ճ��+�Ȁ�՘ �^�L�Q0{�W��pD�6>yPK������ >����$�
/R�c\�_h�/!Y���ͷ�$h�S���W瑜��UMK N&0���0��%��.�ZJB��sQ?o�s���b�:�	ʾ�q~�J	Y�l�����]?�����FARmU�K/��Irc����F����4�pǿ<��A���(��d&	[�D���)���xFK��æ�;����Q�*�{�"��*1(!X��2@�=�LD�2�HD�W������\�����[7�m$&?�+]�ah��I����D�	�3R=`Nt�b1l�L�6A��=���_�o��w?noi��w�I� ג���lن(��@O.���6�N(_�|�����g~�̬�]Q<h��b;>&@�`��l�Z-�p+�e�� �(����mK� l/��:��1"��1��τŧٶݭ�o�����b9Ն�&�4����c;a��mH��ې�a�!I%D�և��VM��o���:��;	P�:V2�Dס���IB�d�����7��L���enG>�AЯ\:�@bdt�W�4��뾽}N����Sq�LuP��,� G���ʿ���*# |�KXer�@�F�/i��t��#2�P��xҼ�\W0�?��k�0ce�m@��4H�����<�
EB�˜5����d�0~7׆?�?i�I���eei����_GrL�,b�p�v.٣6���"Ӌ�cb`I�A��:�U�`8E�uw�f;����"�Qz�`�c�'��m�L���(��q��G�@���gI ۹�x����h�[v�����u��}�8���s��]j�6
������< ��c��W�:P�	6�%�s*h��&q�(��~]���Ԓ�����dzS�&�-��=m�=���<Z����%���֧U�V̙��Վ�F���N�ю��G���:�����Ng�$��0_5y����9��]�FݏLOM]������Dbn2�0CX־�� �[�;�ͧ��lx)�iTW	رtG�J��r�k�����8poƂ[$SC=�����"6��4�n�G_O��@+ً_��z����=W#��k#��@�J!l�� �(Z�[�Ԛ3��N�h�Q�3�,d�m�[�fO���N���݂�˲?ͣ�8�P�/���%��i��'K���i鎊�� �Lvg�d�d�#,�/jb��V'��\�{��9.0��q&��(��07H��L	Ӝ����8L�R���zz=����V�I}7v!���o���e|�T�<"hW��Bt�
������D�Z����o���ֻ[�?���t�g��?��7�.�؅K�a�N3,ǐw�у���^:ޠ�.�����<�r���c;v��G�n�M���kuU+�ݶbb�~QO��|[U� 6k`����E��㠉����.!�<���˶#�(���K��_Њe����aRL����uKW4Y�e?.
:ӱ	=�r���;����z�}��N�B#���	����L톷5�hs���;�Y祧ʧ���&s�M*�����K�)!0�wq�o�%�;BC���˚����se�C	K�Yb����[�e.ka/W�q��Q��l�n7��<&3�c/=���� �)H`U �0�w�-�]�]�I~=�?�����P�Z�JJ��<�wʋ���JdW�O�KO�l�^r��X�j�����I��ĩk,�59MV�kb9��ٕ�)��wg�����b7g��x���D"љ�ór�zDw����0���W�N�f��6�{1r�d�1�R	�c�{��f��0g�s�;]~꜊��T26�̈́M[�u�\nj�~,�QU�"�_���
����B|4EY��웕e�:�Z��gA��:��w �(;fm�[�RC0�;w>P3�C\� ���"j��Gf�ӗ�AQ����"�iЊ�#ǔ12�\��+�q�0C�Mʓ�����h�V������
)�t����E��:җ�ob���
�~}|�r0���btm~]UͿ{��3)t��1��n�c3�J��b�h�����'`�P���^Ng�/�%�l�R����m����Z�*�Rɇ_��E�����oǔ�ޠ-x�^7!�_���ۂ�rwآ�
��a�T�5�~Y��,��N޺b]��LCv-��W�?v�I�rÏ�d���q�JN�Z6�W?s�a5�@�qp{\+/-^�|��f�@e-����!��ZK�>w��ԡ	6I�k�^���Z� K��������G�yw�����w��:�?|��#6���*U��_M��$M��Ʈyb��v&�d�u ��i�#�Р�K�"����� ����x��Y�,��AaG�5%W��fިR�Q���������	����Ώ�����vT5�4���5���X�]!��xBRN���9�zU��&���Su
�_���+D���	%Q*$�GaXܹ���F� �VM������md���.�Wj��8/�:��Y��<	}����qQLM�E�A�	sc��m��{f��ݤI3Oy.�0��	ݺd:���pi˷�O"ޞMy}�!���M�;;D��(F�myET�!i�X�{<��6�n!U*q�j�\h��a��'E��|�����31wo��>������g<��Ol��@#	����