��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+y��mG�^Z�7Y
c��z�&��p��&���B���
���ס�9��j] �&�#&0Wh��p������[������Q��S�{"j�n�n��O�K���J1k�я��)��X G�4.�"Q^�̨��
���ת������:��i�}���J1��yժն�D��d%���������6�,V��݊�#�3'�o#?俉��&�&>�J��G�L�E2U�̏�l]��_������兘7�?���mJA�f�T��]��z�$f�̛���a�����^>�eD�-5�����kᔎ g�Dc��&�0�^��{������p�G��`bω_
8�<�M�	��PQC@f�娬q=cEx����\#�3���]��Jn��_D�ځ�I��%���r�a�����Y9g��L�:ᚄ!6�$���XaA�����r�|q.z�9�R���*���|��L�ˮ{
�D�y���bnE@6��
@W3�@��(�NJ!
���5���XaC�!�\M�a6R>{�5D�F�~����(����I.��$�����Q"��z���P�P�`6��fh�	��%Sݴ��t����⨖)�k�ӂ����DP�PX����=��x�0?�J@����{��|}���Z�PH�P��8�֋�߃����5t�װ"Q�>��E�>[�*��$%aE�&<�SҦt���Y�υ"�
����D9G��RN�B�%����bR�Vk��gZ��N�|=�jg���#,�ۘ�� $an�1B��(
�c^9.�+��,�H�M��O>B��%��Y�Q�&��@���_��c>C�6����B��:�M~��d�\$��$
ਟ��������xb��E�{��@�R��]I,�@o��+��$�f�s�̹Ǽ㞟;_��6�y�W���J�/���?����q����SrY����v�WbP��͂M����ʌX�D���m ��ȿ��g���`�sr�]���-ԌR*�d��KpT�#y	Q�a�f�}�7mƫv*+�ZÞ���]Y-��Ü�S�J�m/'Ϗ��N8�t�0c��P�P��4Z��ӏ5Z�y���r��B�?�v)�vq���-l���7�Zfj����׵� ��T��"[ܖF����i/��Y4Hh���k#v��>�B�m�����6�a���i���@�?\2��}���q%;XЁ�W/��f�oC4��#��3��E�P���ɻ��@�Y� �$�E�i�`E�sL�	~���g���⺣��_��ie=A@�A���>�k�"aG�( Ėm��S��,��s'BE@�<wrr�֤\������D�7M�(IF���Fs���'%����0�_�����((7+TV�7�,�n5��?W��A[so}У=%|�[��eX��u�uC�D���/��O�Ps^�+u��^�~�\?� "&��� J�-�9������$�ux���|��9�jM.N�ho%�T2mE���k[)��[/�c>����S	=4,*���Qφ߆M�ydW����I|�2p��QJ*��9GO�� ���6����S.�,�H��&��y�Trc%FDw�֎��l^���i�z����J�!6<������v�wE�I��o|�U��l)-��+��}��{��o��pn �����v _�Fޅ�H�;q�}�����j��*H2��QTY�9{/|@V^=(빩�G����i��Zz�M.��~cxp�r>FZ�b9	WDҐ�2�/���ά��Y�#�q=��Ӄ�sɨ;�ϛ���M�vc!N'C��5r�����L@a5���_�[0,p�k�\1*�^u@�����/��İ2�u�^�2����r��w#x�Ú�.�^i[��|�'u���8��|߰��@�G���m��u����Y�.�iI*S�L�LRU�>��/��ڋ�!]��!^o�+Cd�]�ч�kE*��`��Aak���z�<�dZy�y��%�����Io�JM��9�i�Y�� AT���p"��s��%���'�n��R��)�ŭ�����W~��]��g�~����b�S8�b�.�l�=�=v��Ods�R�k{�����8T=#u`��;��������v; !�J����>]�g9��^�Y�ʬ���{	��nd�L�ĉ��A��S]<>��-�x�1-��z|O��A��mk�;���+�f�����y�m�C�Ym2�����ӟ�����rR����iGrX�jXo�	i:�:�G�v)˅h��̰}�%�D(��xeF�����RI����Yi���&�qS���+��fII�4��l����-tx&*�/cg,�\�YӲ �:;�^e ��q<c���	���0כ��^�Q����q��>����'|Tݍ�=��w�je<���� �2�4�����-��,y��'$�¦Y�Ր3���k�u�Ji��jC��i�/W�k#Hv>x��M]�`��{[ΌRg(at:�Xܢ�.�i����C\�a/���t1����ꔬ��Ɣ�R����x ��.9H>��^e���O`�?{:ļ��%��N*��	o�υ�**���\��������I���GM{���)c&��9��}V��R��Тe}���a���_�Q���*7i�L��w#�S�ԑmU{�̬_�������࿻�&I��sM�X�����$����q���ȱ]��"�U��u��en��EBZ�N� 5