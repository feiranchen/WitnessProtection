��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�$7�&"�K�;���e�oG|!.O��b���nڹ�:9@F;�`Z��^������jy�ݧ�>��P4�}�����T�
vs`����o��	�u�����ɹ�3o��>g�|����̓ @�'K��<$�N�h��?Cr�*-�E��O���0;���6C�sd�5Յ�Ц��ߺXV�>����F0�6M�=BCB$	Q���oV��Iz��T��fsW��{�ПZ��<衶hwh���M�2�D�0�a�c+�U�tH�W�R�e��j)�o�ȜV���"�r��"!B
7�r�o�!li@((�RׂE�p�r�����t�lG�7)@8^+h������E�=�,n�]U��gމ�����07	"�ʡNP�`|_klŹϯ�:���A�$@��Ι"_OS'�52/1�(�i�RpN�r�a���ܗ�]�S�	[�9�Z^�@o��>��^��-A�
x�fD�ȝx}ӿ�,��/",0G��K���!�lᆲ��M��|��I1,��ǩ�H�`\t���A x�AZo�]�r���N;�%ά����C,H���JAf��;�`3K)x���bE���@c- e�m�qܪ�^nV�dAlV�ST�j�,݉���i�Y$@~��<��ٶ�.x����1v+� �N��5���r�~���ƭ�a�WӠ�69���7c�����YEb�I˄(����`>RMF�__����B[N����^�d�߲�2�������X��@�����*G�!�Q��?�s�]��/gW�{Y������Ҹ1y��_HI��
�`�6������1����`���*�|�>V�3G�(���|��E�L�pȍn�`:�͟�����A5�~p돔�52�VF K2���=�#� ��&���Tv�X�&u)l�����=d�X5 T3�`sW�kj �|���HQ�-���z���hm]v�VL^T[l$ס:	=�-�J�s�Y('�O�lx6Y�����Kp�D�^�ۚ#��|-c�2/#������:"���m����r�S��5>��W ��KE<�
U#�3�>y���&{�P�����	�1�(�~��w���31uT|�)�z���n�������b�BNJ��/kc�i����;]#���V��� ^�"����oK*_w�9R5g�e+hr8���艧b� ��4v�?��o����g⊸��u�f�1��vkfS��7�����a�->G�~T�@f�J5�u�t�e0�0h�n���J���u�+��_D�52�����q�l��^m�6�;'txڅ�eH$I~ L�m�q�", ���a2�s�>�dJ�mLƦ-����U
�s�|F��=��i��2��qE���`��	�\�����U�E��4?�!L&u�e�'�������?�i֧%�_̟�)�*�?��tS 	��9��!�ʥ?9������� ��*я��P��D9\/t��HfT��别dT��*��v�ID��OgN�y����*�G��>R�G�e����/	�h}P_$�me� 1V%��m�R��˸����3�a��=#Mʇ6Z�ʤ�*xְq�	��!t���%�;v�6����@�����M���w���v��a�⋍C0�%��#���Nf�M��LR*g}E`̦��/�`yn�w�!<#�1"�����t)�z��A����8�l:�w��v">�X�84��2��2����1���ؓT^�L���WA�Dp���ὓ�d�QT��ShV� CJ����|��!c�
��Ic�t�u��(��x!s�P��v�W~�O�|r;=�K���C��,5N����ZD�|8X;�p���C^,�+�H�����H�W�$O��R$�>�� �c�E�6�`k�1��y�-�� �er��G ���.�J�$?x@_ �诱�U�֯;��A�8q���U�4�V�~~���4!���²���n)��/��Q�.$�F���[�C��o���c�*����(��5<����m��J���7?18)	ݢR� ^� �W'
k�ǸZwg��Կ��={Woq~�%dWfO�� �ޗ�W����;����4�>�x���1��uJ�llߔ%����s�:�����M��BH�_�)j�0:�w��lK3����
:%Q5��w�F-~۬
l@H�k�*���ӫQ>���|d��c3��SE��n���Ǡ(\n6�Q��0XC߀��S��}����Q˗#�?�=V������6r{��*�4a��WP>ض����{!P��Z.��>�����&\��������0���N�H�Kt/ht�]]"v���ށ�L)�[�������%� b8�i_�Z��;�K�)b���W���������CYw1���J����7� �c㎡����a:3�O�Uy{ںp� ��S��М%�W�n��2�p72BN0�s����������r��M��^�wؤ�&��K|r�3�
�����)�����>f�+9�����,��[�	��m����4 6�C�$,�eyW6qD��p����qX�:����]oeT@݋fC0��E�p$�+ܨ��v,f��>
e#��� n��z �_W-JG���bv����Yx����"���֞�|ś�`�+<�FA,<�ؚ[pP	u����f��p�:N4�])'n鎉�:��3B��g ׳��eZ���;>9���p�W#�h��A4iE�sv�ndď��t�G;2R�����B���"�h��z�^MM�T�Zҫ/~5m���X
e��L��̭؞l��a�0A���d��Qɇ�%����Pi6jeF]���3qߨM��$>4�UA��n:���GXHs@d=f��S��� ���Ȟ웊��3��^���,� ��ˎ@�A��S��o�ڼjg>����*j۾��^����ˈ�z�*�GH e@�r���G��o�2&��.M�#�6����=��΂�#O��H�n�4��ɖ�B|[MHFP8~�4ԅ�\ 6�s������2�Ans�6V�pS�ha>����`�Zs=C�6ޑ�σ)sת�<`�d��%mgUstZ�p����2���K�@���5FTn��:��*=��Z��v����/�Znkuf<ƣ�pO�����~�3I~����H3�aE�R����=�BDA�q�[ͷ��BV�<�w�4��!Y<:��~�����c���gGz���Сo�ҁu���]?Z�y��f5"r�j+�1�0��o4g��2^P-s���I|W4�Tu*�B֎U��c!�=�rw?��M�b
0�.T/&�2H2H4iI��S��n����^�K��h|!Q{\6���-2��\�|(�DI$�"��޷�����N���6�O�㙐Q�N㦎�şH��yu�!�^qN~��0spF�0���1T�v�#�)O�R�ꄑ�t�A�����"�G��'��؍"�*gW��qؐ���!�Яc�P].��9�L�u��K&�Z�]-����
.L����w?Ė?O�M�}�y�GG�L�B�/���C�o�Pqӧa����p�4���[��Q��#�9L��*��Z�����΢�'d���a����{zw_�K3	Gwn�z��ǒ謥��e��T����U�f1B�]S)������&K����]�/�V��[.�,���K�H,�z'��l�̒���U�_J�Kn���LHb.������:��"5�E3]=��`�mҕ?'��n5&}%����`dw#��%��ThE&'`�}?�4�bib���&��h޵g�b�Z\��yb��a���W��*<hR<�-�ݭ�*��PL|���E)��l��h�mn.��}D�qt�`�31D�8���>�T����

O�P+4=TL<<��˰2�h�o���e(PB�ؗ��ge�N��E(�/j��7����l��4 �k;����M͏Mu9����b/2�.����*��L��4K��s�j�@]޷-	-ws�g	�o��w���e#~��ױ��)�8�>d�Z {�L7�#"�;��HP�B�2j�$����otn^����r]<�A>�x����'.sV��U���sJ<��m��.r���fq��uC�ٰ��T�Aի��?��F�V��;�M��)��?��M����+�6]8���z��v�*?j�.�bV/vv�c_�?֌�GޔN�+�T�~Y���7Ŗ�R���R�%�w�d���H��7�8�G�8��{�%�\,�:)��q� Tk	w�T"V\�
�E �jh�Q�kZ�� �P+�9�_J� ��թ�)�_G�c�B���[q����ˆSٟ�Q^^�Nz�,��zf�6���~����d�m�gbT����ˢ@�y͗��R�����R��ih�a��$.'� �M��fXQ��OY�0ԛ��4��*����C��顦�A�'z-�����[D��s���D�QVF�e[W�,�z�1v�([p����L�z�Ҝ��T]��&�G�Q,{���QI0&@� ���s' /��i�&/���h�@il����� ��{M�J�lr�-��^������!۶.��X�I,G7��A���}�f"�u	�Qq�7��!�|4㠧�甂���q9��F����kT(/7�~@(zp����FIh�|9�]���ރQ+�P&z��)�B
=�|3(�e^�����{wG�P��ܦN��$�[��4�C����5�r������g���=[�O<�!�G��S���շ꧿s�6�l/Y�7;�Dc w��=�g�uqP"� �n��f�P1��f�~���ǂ��8����2��7Ic���X�\�^X���^���}��p�Ph�'Z��٥���⳸A`�q)��D���z��$�=2�O=[�J�*t:c�*��T��B;��rGJ�<+��ѐ����V�éu_�k�3J��q@�+�j�nѬ����߇�v�fi�7<�6/D�M�T�;Z���N������a��H���W�ͫD�f�xC��(N���2��r���~���u���B�ΫN�Qr�ݮ�} �V7�����Y�����Ny���W��%��QCE���u/�.����k�����}��d��[M��|J;n��h���T�Vt<k�`a�	�MM!�qML�k���\��^����K�е1.�����'�h�;��,�	S��
%����Gtqr�o����p����0
`T��X�Y�R�ԇ�$�KA(8垲V1�.���A�����$��ڢ�#��G�I��8���D�}��(ƣ�<\q-���MB����K�\Z�;-cN����[�%����w��Nn��\$K���X�ô��"�
/�Gs��A,�sp�B?������h��%ӝ���?'7T��G�"�m9~d5���(��|�Sr�f0�s�{���<�k@[$�q�v�޾�i��s��fw��9-V7����ڱE*[Hg�^�eE�G�nK������Ul��Z.J��}��9�Ea?�S�d�N{�I����^"�mu�2���±�O��êx�"�����D:�W��$G�?�h�|Q)�K��T�J��6rd(�A4��?ӜX�2���B������z^�7�R����#�w�րy:���Z|��]Le�2�U.��p��Q�	�K ���!:< ��ݰ�M��
5�0h?�.VЭ��L6~N����Ƣ�Cx��_T�<����Ҏ�������c�&K:����@!���Tw0�B<_);D7���%������r�g�^����5�C�$B���N�Y��/<vv~����bW>UC=�Ϯ�O���]�,x�����%�ElＡ�Z�V���(+p4g6�a
��a��U`J�Cb́I�oO
��L6*<����R�ۋ�3��0Y��=��BJ�,1Xeoq�u^�]F���gn���mJ4�N���p�jָ��С�|ù���67j]J�~E�/�	o40��Æ�`%�y;��E���
�����1|z>RƑ������;C)��V�:k��kc
����7������M9�s;q�����FӰ���}0��Ť�6��'K;��N�!��ih��n��,�1����6�j5j�2���y�