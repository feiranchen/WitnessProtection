��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ{� q:4�ZH�]A�u[�����[v����hM��F1���&��؀���C��@�F�zuT��';N���c͹��3&�� W�S��oE�d�ƺ��y�ݣ.&}sn�Q�		{�4�ZuR���QsD�/�b�P!3�j3�3@,OW�ZGc#Y�aF\���y��;?�t�3SJ;dy:����RR��\�t�0�����'H�D�Ll�w+]��l�@����8J9�.��d�b+B�Y{�bح�v����e3����8@A�I=�7FTA*�7̦�vf�5T�u�	����+_�D2��/�a�>mx��Ad��8m[!L��{�o���Z�4�*%'Ͱ{0�щ:���(�M��5�d���������=N/��h��7t�S���*`;	G�#,�t?Վ�nv��PTv�"o�$�lG��I�S9�[�K�燯�_W=�X�[����gΊ���PY��?�K�!X^dK�M+����d�%�?�rR'�&E8��h�c�#-9d� �V*�-ǐ��+�?40����ꕔuy�K-L�_����}� �#�J:�C��{�C�H�m��W�S��N�����5�V-|��>!:ؓ�I&zg�m!����[c6��<R'B�t�C��+�QX]h����`|[g{~z?�/�����QY����P�-����?𺝖n^ȹ��}d�*d�����ȹݲ|�K��i�sj2=��SQsh��]��X�" �{`��_��$�i!Շ����ߢQv�p�TP*��B�,���T?����9��_�:ǪS�S�^��<��_��/ў��B,�\�ь�)�}#M٪a�pQ��l8��-�7��ú��Y1�:\���e:a0o� �h��r_���<"h�Xw|��H\9Ƴ
Y�M/v��&���5_�nxP������Z}�`Q�d�ü R��|^�@�9��E7�Yx�T�����)Ф�Wۦ
�y�f��?DâS	C�(7��w}�A��B�V$3�R��#k���A=ң�cT�Z�O��򂹳Y{|�b�Dw�b�����86WC���L����K�N��_�ny6�%a�u$��G:�0JS�:�Zl�B��S��-
������k1#X�2�!���>��3L�]��n� �qW�@q�C�ȏ�.S��Z��]�v�o��o4��0O�����2A%����P�m��.M���@�gv��� Kq�Yn+���'���nk��x�?����4��� iG����6?s^ od����R�ip���=ͮr��В-�,���H~Я�v��-$�+f� H�IS;CC���q3s���0��;w.����+��4�M"G��q(�J�u�8@{�ĸlيj�I'P8X>�x�����߬���z�qSO;iD�m9���~Hw����S+�hN0X�P@9�t,�c� ���к,���f�讽Vd�Ts��2�9�7��G'�عզ�����Az����Η���9d0�;��#�A� O�&미�fɮ��R��k�cZo��%�I�� 2C�y	�����x�D�y�Ц�����<Yo�K�_����C��_c2"���X�3L] =C�D?��0��B��>a烌%�R��T���\�QW����S#.������^U-��DV��e\m+�$3�1��wr	?;����mM�;db�7K�����1��M������6�%HYa����=o׏��`2ċ:�R_��FL����k��aE+m���4�K��d#�O�ܒZ�G)8GFF��B�Gd�0�u�L��3z,I�,�^�?��7 �3C�U�!u2���;Ddf7=W?��4�%5�  ǰ48���X���۪=�N�u�\�Lh�g�p���7�)��4�)]]�ڧ쟳$)��o�B���@0UDW��w*%�� �iSx��6��ͪ	�Dy|K��zZ$?4o��S򪃾?��`�z6(��=!+k�O܍��:t�����: IC�u���Ԭ.��d*E��agUĤ�t�,����]����KɆo�� ܹbV7ߕ��w�� ��V��{�,�p�x���Z��������|���'�!�3�U�%ƫ�$xD�nkL�Di=�M�(w/@��K �����a�yST�R���'-.�[�ln#Y�`���9�jI��^^��$Q^�d�ϊtmj6|���˒���!&x� `E�]f�����\�[qP��͓��x�`y���ZUGH���X{�^���s����S��r~��(脵�TP7������Ϯ��d2#�Ȃ����<�ha�>w�S����j��/���V|i'1+y����?aP��_��=���)����묉��}����a0�j/�������ח�9���X��G~��Ekn��|�����{\�c���!��7��ǢZk�BGb�:����#Yx�'����cu��E9�\��o{jIg���ٵF.��h���ՁC *L�ke�4��4Щ�_�È���PN��W@x���!I"zd�@�����N��(�����wZ z=�!�"[���qn-Ԕ+�?�v����_O�u�4�'n������S��D��4{Ћp��4�b8������p��mb����&C��+�-6�(ǌ}gn�ds�_����	}S��^�O��G�-Ų�QŰ��}�5C��l3��9��+�X������=x���4�*w6��.A��pnL�%�՟�D:_��nr1Hw��V�HEFa�k��D�54`�����7���!�j`��k��� w&�+V�J���\n}�R�H������"N(�h	�v���hN�$Ƀ*��9�e���M!o*Ix�c�Uv���o+��Cr�	gc7^�y�g��ϩ�[�BG!v�/��O��Or�h����:Ǖ��N�m�#zf�kOq�(.v`��M� �� /%��d[	KaoC��/��И��'���*��~ln�xn�6�m��©�i��C���y��З0�o�GX����ڟtISX=_��U����zk,����XX
�<��B�|�:K|��bG�>/]�/�+�sg,�K#*~�r<P�YӃ���Nqs���E�TӢ��b�K�Z���#w���oې�Ժ��j��^���!E��j� �%��֗R�?����V�$i�ֆ�:�w��~�_rI��Pl�(,UZ���U�휷�4*u�Dg��-���'US.1�6��4� 7ۂ�vL	u��!e���!Teb�yK�}d�D�Ϧ���9���v{���o�̅Mvo�H ��~S�ǿ�W�ļ$ /�Abm���o�`���}-��e$o��ax�xX��gǥ�d#���7͍�Hϵ%�y��[&#种����{x_�mS3��՘|
�ފ�[%M�B����a�}G���(sΤB�/")кtxu��G������T?]�YQ����S�BHX��<���K[$��6E�ݧB�4�G��2�^-� �b4xx*Eg�k��h���D>�D����V��$ ��Ԍ�*U�iP���N�݅8��xT"�bH`)⠿�K��GY��B�i�M0�p�=���j��W��UOݷ�c��d���5OS^G!M�k.Fʽ԰�ՋbVzE]�!��)v�{[FGL~9�w{�ʜo�-n��dQB<�Pt%���S{�~����*��^�Ə�	��ɾ��V-z�!�'B����S�v���|Y��I��gl!���b%8��I�&���*�z�+d/��I�q�����Q5���\ͅ �<�V���=jhw�P�	����!�����T<��}�ؖ�`FV8�b*)2bKT dP���