��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h���]��ZBq'aN#y�L��,�&8RG/���.Rh-��/� "	m)p��N��ï�li�δZ��U$�/���зk�BR�:���M��BCz��I���>D��ߍ6d�m���:�!���s���{}��ca`�f!L� =q�^�� �fggK�4��[�$��1�)�f�p���لt���&r��<p���Q�H���H�����%-Z[����*��]�Y ����I��F��4�[3�t�#U>�̫�����"a�9�Ls�k�C�Y�l��d�eH�����AD�"{��'YQ,�v����j�|��0���j�<���cZO�c��}v�Y;r���\_ZZ}�� �����d$4`�{lE��;Nu
9�U�) ,�i�n�7�a��^iG<5�C��Ր�𯲴v�(�vQ�AW�G���LhI%���B詯Xk����,2y�.M����I�9� ���i3p�h*Uv%��ᇜ,��t��H�\�����
�X��e|S�DN�|/u��6T�TH�W
9��}���^{e}쓁��5���h�v}�4..�Q#C��y3�t�Al�� �.��G�n̻e�Y����:	u�o8�h�K�-̉!�D!�����m�,����~���D�+�������3U�(����/�~U���[�����쀏s^Ӧ���GOm'+�m�}oR��&�B��e�IK���D�<�]����R�#����߮��ϟ����(�9ͳT��ޟ�2�,��3 ӎ�pl������txC����V����]�Pw=�ݠ�G�lY�Nx/�����]{_f�چ��ߋ�N��3��7e%���L�����؄G��?�Ԭ/~�*��M�k����([���x�/z31��k
��V%#W�o�?(���g�P�����=V0
��t{|�Ү�u����r����~�Ė��'���n������xb>[�/�X�4��V����j��.�������j������կ�dD�Yy1�!aR��˫'�����	�(���;���g�F�J��{��Kp��駶L��{�)� �wu9��3l߿�h�����,]C����G��=:xC��l�����"ijb` ���a���Ĭ��^���M.�4���\�}($5���n�o�*�<��2,1x"؝d��얅����]f+q��������#��-9�[��F.?�<�h��	ka"fN��o�H�[؈��̕�c�Dq�4(,$��<���r����=�y��D}�fw��嚫f�5�mmA�ƿu�_�(�:j��)�h���E17�B��d���(�hu�$�}�!(yT8j[����Ga'��:q��@�J��R���g<� PӞ�Z7%��`�� ��C4���{=�n��ƍS6Z��� ���SKB�-��.wC��i4bY[���T�28�8��ӻ��A�y�i�N?X]d5c�(>�)uc5��Jʠ�"�) fj
���Qd��J�~�7�B��bsQnLFx|��=&Y燖����i��ߥ������ţ�٢��M/�&�*�fAP){�:$�7yb��Mզ7ػ�����ى0Y�
O^����R���ޜi�Rt��f�?����kfF�65X�CC��1��;����-4��E�\��	�\UOU|�>�7� )=Ֆ�8�I�<i�xlL*�ȀLw�yi��̌�T�C۹��;��>3�e��O�'��W.��<�5��x��i�X"�bf��@{P��kev�@�N�=e1S�B2��oc��K�՞��m���0<&[��fA`��Y󕩗U��4�e,G�P���w?�&ؚ��-�������,M��/���"(�m���&z���>0�����DP�q^��U��_�WW1�=��D�Ti��H��ԡ�*�ܜt����C�}�v��M9<S�WWj�~��Z�e7{���1;8�b���^^h�D��r(���ݝq@@D�@�C_7kh/��a�x�-��o��$�&�8���nŇ\Y
��$H�Sp�mwO$)�ȷ9%"#�{��
/��QoYB�%�;c����Ŷb�e��s�m��2���M��J*=��N��!��rf�v"�s=�m�`���_�作ڔKu�˒���+��	/����Y0/;�ˇ�S����x�ȁJ|��N�;kwmB3�>/�B��o��?J�4�������y�Y��ͱ�7�2\:�$���V�*XIWF����Q��y����$�b��(?j��=�UTzP\~p��P2�*(	a?��Y�+"�m����2`k��kh&�i)�B�o��.�]�ʽ+~��B�j���[�Q��Q��#[�K*��v�"�I��Y�x����ʗ�MX~c ����Vē�������)�y&�i<��,�i}��H�QbObh���䤿���
�;�\;�p�sFy�V���+��{�� ��^�%��'���#�[�h-�����F�Xn�tt��孹�������
C	��g_�c�����{&g1*iժ�?�W��l��;md�������A��b2���8h*��0|�����q}��^���Mt�Nxw�?��<�7�=b�g��.'0Fw�k׵9�ڷ&�/3����Q�ST���_�L���*���Y$��W�[BNY�)B���iPyQTviݦ�7�v��Sv���J�����gxm�El,&@�I�v�l��Q�>}��7��赎�F���4s��ռ������u$w���U�wT#?�+�qU�%�<��|��@��L\
�
	 B�b��C�I��C�ܨ�`3���:z���S�J�OJݫ����bo�w*ވ�	���?[O++
-�H������6�)��+�!@'SVtd"���x^-ů���FpN�u𛉼(~�tZw_� H���I}�|7���܅k܃0?V���m����������ڊ#Q���K2;��9�A��N�i���H��^BG��iZ<��f���vN�a0�3�Ms�B�\���g��l�g��.zwJ_���\"�7x�PT�*:�c��H0����1Џ��}�Y�`�SN�`��i}4��(��21O<�1���4�M�%�0ox������9����q/�Fj�W,������w�|д�p៭�Mb(�:>f�Â���Ԭ0&�$�e��_�����
���<}ܗ
vjx�������^��3���b��lj�����	2��h|����]a��:=�J�uy�ق)�e��W�˰(hFXE�6?��FE��?�`.��[�\�w�_*=A�g�6�ƴ�d��R!gMP����/����d��@O�C�ϝ�^�BG���(�������_��ˬl��[��9�Cƀ�*hn�XJ��.�#Sd���o��� ��T���z���o�a���X�1��@�(2:�d��x�7<� �� �vt�}3y<A�n��|�� к�D��4�Ĳ��C�/��]�e�(�c[L#���<f��"��%���&���)��VD��r�n*=hL}nt X1w]��/��@ř�����c�Ԗ���BA8*�g���H���2Q��,[��3��N����󈮗�����s&�$�+��<G��-G�$T)�L���N�J�DU�i<��"���mз�ӘV��eT�wb��+����d��S!ʧ��za�϶:u͖`��!_���y(���l⤮����SV����傂W�q�;��u�h��GP�x��Zf�������_����Z�5�zu��S⥊�T��=��u��g���Ƹ�ca�ul{m�v��>xY�`�e��7���_�ʠ9��Mo���g*�q�gWt� Qm��o�o���/����\y�s�J̜�zb[��Q�B��~�q	�0�f�KZy˲��=����;���r3�7蔟μ��>����[���o-*�F!�Gu0x:�;p�y2�g|$l���%ev���v��R�(�o�{ω:q~N�V��Q��.��$>�k�G�U��bP�*�<=��V_!tf�{)۱l�>�{dR��7(5�������Y9�wrC�FgW��U(�a�����7Ξ0E���(S��r7�4잽W�Ub�h�����r�1�}�T".H�C���s7?�-j<��Ⱥ�lm0��J=8q�a'I��72��s�<^�4��4l��.?����3�KP�JzF��_.|T��H��v��)o��=.�� ���HԬ�׾.C��E����˛v���;;_�N Vaȶ?��m��fSwѽ07�9F�yop	��K�vx�Bq|�԰�񮓋�>��s���C��;E��0@���K�fxR�f`�Fej�ő�Ӧ�o�2��36M��C�^:�fQ�^C���Q���G.�DE�����§�B0��1E����>�-�Ɉ���M��7�U )@���P���G6�d{�����d�^�&ħM,'�D��sE�WVO�9�!Ƴ�Ԅw��K�`	p0ށ���.���� R��4ʅ���*�е'�6�ZjV�2��i��e��C��7�����h~2��ZK��|�����3s��ϝ���(Dh7 �Y+���f��#y��"ʢ�5Ŀf�n��-��)t��3aE^�5��s�g�uF�B��Ȏ:.�xwﲓ4;`��Lb�R���:BF�RU�&��p+����eG<4SK���e�J��q��]�cʆ���i ���Z���Z�q����h3�X�ꐖ��r$�����6�sc}[ǢrP�6|.��!��J$�Pvц����8��b(��8]#��e#ֽM}sF�E�����-ҩ��-B�&�^J>s'�"��E]��FAK��Յ�I���7D:H�#�Ȝ�9s$/���ԟ�F���[�6I�
��3/���\0��惨����-��kgʡo�nO�%��Z�IN�oYͳ�X��G����iPRX"/`���8�W�J��1��^��;�Xtw?��鵲#��]\_�Vk�H��WJV\�x{s�Y��7�l%q�,�;NbR�ZX��[�z�S	D?={
��<�3ؘ��D�e���n��C�}�{�5��W���
kkR�����?� (Ih^�Ԣ��r�$���eeo`7�wջ�_��9�OzjSR�rR���t�1�c��T8�	:�^����(����ӛK88J�����a:��ƀ>~�����l$ϵp�Q8#V;.���ìU������K@o欶1<�lA�;A�̩���`1��0�������l�X�c��N&�\�eOD���1��ϙ]E�(�Oډc�hN�]/e�O^��6f�Ι1��?a�֞�mo��}���#t��]���m�rx��(e��u�^��T���D5���g�r��G�ߚp
[,���/>�iiz����TV1��)
)�`b:�q����}%���/iHK!�)�k��e����׵�S��5�1�f.��p;;GX_ � %�.˦��Ĭ26��������"��{C�~�Ț~���1R��lx�)-e�HO���|˨ҿ1ʥ6 ͹N�Mj�D���E��:�ǃRH vNr�wo0�-�o�j _k����/������8���'4 (��@0%}X(�X��m��.}a�xA:ۡ�{�u����7���t����/��l��4����n*�r�Է��D��xj�__�j�*�c����5�1D��H]<���3H=}Y��ю���j��ˡ�P0�a��I�X��T=���x���%��7����={����h�28T�}�X���c�F����Ў4����eĒ��^yyI�iwO��Վ��b�*eB�J���"t�*��)/���W�����O���=t�9{1)� �^���� DŲ������R�V�;�L"�F_E��RK�������e�Y�a����^A�����/�OV�p��1���8vo��6�J� 2< ��bC��zܽ�^
����]P��9b��1c|}k6�����q��4!~�=�|~����������%��a�jP��Fz� ��m4���W+o<��F5& �sE��k���;�b�b���7��ܜ+.�)�璧��%���k@;�GyP{z4���'F3�t	�.��gh0Ih���8��^�?[�����5G�`�PqhH�nvZnGU��m	x,{l4a����^���'[���3{���O����0�����Oq���u�V�����$����ё�U�g�ϋ+�$�(η�T�xG7y�:�բB����d"���+߉�~�y����	���G7�k� Ǖ�b�̏r9P(�H[J����+��=8@t�����������:qƑS�����W�VŖ�d���^���v0���W�=��˫Y��妵��_�yYg��Dx�N~BPTm�L�%��Nq��L��:ہ�LJp!�,�Am�ų�U{	4c �߇��vƬ�n�p������G��	� ��(�G�g?�rL�lC��0+�)�{�,��&�f٤��\�ʩ8�}�E�lT�_����Q��җT�D�L/v���싘�l����)���1�M��}�,-���ŖA8���]�n����T	�N�^�s�p�±�͝��w��vEꏶ9�R�����C��1U9|t��*��)G�LM(v� ǺvI �8��[io)��t���tHJ����oY���]��u]��B���D�;�Xۂ�&ص��0�Q�g�q�P}��١�B�;�sP�wud��K���K>_M^�χ��b��dȃ R��"q7j�|�v��uЊ����]o㟰�@��L�)S�{�Ʀ>_s����90�pt�At��[{�_.2_5W����E�u4�"�bd+��y�&5P�!���L�#�y]�%g+&E�U� �4�I[�qr�7�g��6�2Ҷ1�f:�Ѵ�t�ut4z�?���B�?���h��#3%v��y'%��'1��#~�Me@n2����B-�:���pu�׎f�������ot��_�gΪ�(%T�	�㓕��[�ejM��������?kݿ{?*�#P�NA�2�����������"(��w�.t�B�v�g�Zk��1�,��~�4@��i�TU�,��`��ny���H;G�D�ú���U�)��$�v����L�cA=�e�$_�K�n�A�S��w6笆�o�����%?%<c���ad*g�d�u�=l2N�a_�(�����$���|��n�t�������z� {��9xЊKM��b������ʍ.zL�Z7.�����n��ؽ�P��$Q2�Z�)�	cy����p�N52�;^��!p
,��sof��3�6��&�U����y?B:B�Mm��b�GFx��/%�tl\�������;NNe�ů�_�3����iH�t³Ӥ���1��	��W.��(��J��ǣ��K\�16/H��)8�1c^+�t�,�5|�����h��_�f��A6>ã���ǥ駨� |��F�޽�������<�O�pyI�$�DZd3�z�F~�k��<�Xd���ȵ�����^��RO�q�ǠSlU DqP�Qh��RL��U��-�T� ��W-��k��6�P�:v��˜�e�'��:�d%^��d6&yyG����������H?���J!�9G�R�jѷ������v�j�j��8�0d�s������PQ�Z[��,�*Gfᯥp���w�_�S�e����@k��#	.m�u���u4ɽ�,d
�xz>5���f[Q:f~���9��HV�X��f㥵W��B�A��QANە��|i�����]9����Zd;��s���oӳWK4����ue�8��|�IĐ��)܌O�	�*�-�I��qcO�G��I�[x����b����A/�uy3��H��o�bp,!XUk��s�G�G���քӑ�iC��m�	���R�jMA?��9 ����2^�@���Q�S0�.?�_������\�=�u�[�wtݕ�"��v�irI(��#����'��z5�W�e��;�p�LZS����]ޮ;����M?u�����BS�!�.�x��q���՟��|z�)9���
�G����d�x�f'\��~��V�r���<
;�#�l�؋���e�9��T"K:�RQ�x�L}v��z�=_�B+�H����;~YX�����kØ�y⭫���t�k��z:�������_^�P���3����6G\t��$����jɡֈ^��Y�ԡV��ﻷ�G�f��/�[�	`�N}����m�r[j�Ԓ�mD��#U����x\k�b"H��c!A�ķ����U=�nH��xl�}���[�$h:+��DIz`��8��\��ɀ/?��h\.�c����'����ΗJ�od_��%Ծ�V�.D�@��YP�kv|���pIS��nх ��9xB����� (�_��!��;K�Fr�\�`��x%]{�P�����2���O��K	i8w� g@�c�Ʃ <� ��fUN2W�� ��o�ȝ����7m�9Ѫ����HwY�V�2�vH���2�y�(�id���~�%�7И@	��M��%8�8�M�"xI� ����Q�0�z�p�[��M�����&U004�b�_7��jQg�M�������(K��o�uo=d@����Z��(l���i������V��U���(��ڑN'�٢п�����qd�<���0�s�?څ���.�J�6�;�C6犨�m�v��-t����`r:#���=q�*�2�,�� *Q'mq	�U��ji����؛"~�j�qN���h7�蓑dz��-�r ���gLza�y�C	S�4�-1>h���5�(|�YL�N [��_��)ef̠37��.�%O�n��[�a|0�����}��7��5�F����	�~('sk����� "�1I$U��X���`������W<^� ��T1Zsy[Q�� �W;`��sKu�?*��1����ͣ��5J.l�,���O��t1� Ԟ�!c7Y����h�NtXXM���n�pA/W��t��y8Afĝ�<�j`pXuq������T�`�o?Ɯ�R|-�nJBw�;��΢�
Bj�^�7H3^����������^�����pCФ����7�dp�kYBA�5�P����/3�n�>F�(P��7$�&
�/�a�c���6�c�w�7�8�l#�?�PC��6l��g Q��$
��QB,i�O�Y�Zω�n�h�+s	x�ǻ�^�C��@"��0k�H�/�|���m�z�̤�2��m��Q�8k�j�վlVB�gÎ�����?�V�@��Fes-�pY��+$}SC���OO:��+���������82���Vb��Nݦe�B�|B-q���a�����n�p2ϓ�7<K�����v���[���՚E9B��ڨ�EG����jS����2�ѧ��Q�Z�c�W���e�'A�ٗ�o�al��Yay��#�'Y���I�8vgϸ��T/h)��I|���h�b7P�b��$a<�#�8��X���z�>9��l�3�����S�̰Q�����Pm�xL��0)��YL/R����m5�v0���0;�綃e�ţ�^��\��.�ČVa�q#h�v��}x\��|Gm?BO�0�B4̛Ef����H	��� �����T��	��&�'͖�k��éD79����}Y�Kn�)�����.4���/o�ߦ�D��`4�7-�M�Z�� 
�����QV���@f��v�D�>;��dWS��`vj�.��8�ci����i8
�kv���]T��*4�B R���Mσ1��smF�,(��0&N A:��I=؝��B�@x='?��^B9�W��`72J��b4SRu>O�,�k5m�ر����Xt �-'6�t/&7ѳ�����t��?��u����
�`?՘S��5s����!�^Cg�C"i�P���ڗ�	wU��h���G� ������>k<��Ώ��qh��"d�7������������
My3��NE�Z��p!�Q`$�[NxD��\��pW�)ۏ�8elW����}�Nα&�ʂ6�;�����G�4�r������S�E�x���ģ^x҂&	�Mɇp(�0�fV��101�M�u&�c�Y)��a� ��v	�Ol�B�`&*ɷ윑�
��_�b�P��/�!Sa�:|��uq����Jc���Q���}{�)4
7�J`�PV���{8_����dq�"�F�>0t�4dr2\PB��b�塾[�Gh=���n��7b��U���C��b_s*�:�4���O۵����O5ꍧJq�	��^�-��P�-1P�-}�C�2�@>��{E���w�����~A[O"n��;��oc~�K3����P2�#����E6�f���lև,K�E�j���p<x��u�Q�H�G
�Y����)4W��4�G[����U�Ya���O�l�n�[+_|!����������{�c�T���1�]ܞQa�"�N��Lӫ�/Z.��l�OT�"��d{XW ��E�u~anK*���	UmU��K:�NZ}��nDt[��@��J	�
,�$������>���d#���YM�Y�.  ��b����8U@�Sy�߸��?�{M��п[���0/�<o�=�)q!�t�F�#��2!�J�.�bcH[(/�����iv���+[Ȟ���ן����D���o���H�Q�*r�?�)�S*���pY �Gԍ���yPN����L�S�|��7&5�zK>02�
YoP��>J(�=��Л���^?�.��c0l|�eg��W�Kτ�W�H	}�?��M��r���/f�w��"�tK|5������"�C(����S[}�~k=�������T�i�k%騧�`bѯ���,�[�+\2	?�iN�o\Z!�"�R��G�B����>���a';Sje���S���5�<���C$P>+��hF5V��m��n�4FE�3�Wt�L{h`9m%�r���_�S�hfU@$,�q�ۈ���(�Hfy���۳�|�'�β���@`!�������du�#���ѯ�i��{V
��0�抢�}6�jQ6 �r�����6��� ��.�v][��g˃q�pu����+zUn�E�&�u�����4�{LY�"�.�I�W�ӋF�	f-��iZe�����JK+��s0�ׂ��ό+/��/��)���[2��	A�eأ��H���!�=K�� �iL�^�ۑM@��/���1.uت�c�=jjMah]3���q>{򇼜-�<O�r��f��n��7�1͢�7�'���H��#�hz�E�Ǩ�|V����2��\Um���	��la���Ka0c
�<�FM@�4bP�Ɛ�o���5,��Qq���/����LI_ùO]�i�d�;�%h4�|m����,�|c�:=m��/ƣ?�Ȕ5C������ ���������{��+E�E��%3���;648�\�zKY	U��3�Q� "3@��g5�� ͐՞c��[V�N�u�%�N��}���/M��?(g��Z!8�仳v��G"�=x�X1{cs�k\C��c�Z���.]r�b�-���ǒ<�4���&Ӄ���Ob%�Rėi�?��/ŝ��C�<j��đ`Es@��ǃv�v���Ih2��6u{���[��H}<�-�2��Hکۡ��f��$[�3�P���ew5O�)u�K�l�rN0���Fӽ��C|[Y�Һ�SW��[�Ǧ��+??�dN-�rc���Ė�{�,#G{����;~�BR��j�F��6<���"�f�rC�)!�G�X�R���,�\G�&E�0n�vu'@�3��r������̪B�:�ޔ�`Hn��rÑ�)�HSt�Ӡ���k��Ϥc�\���Iȴ�9�ĥ�ƾ�5���"�3-_CQ�z0a6����k�M�R��K��?^���(�&��J:wT���:��><e�Q��M�i:��L��T����]�$w�>F�3Ԟ��ھR�⠺]�z�g+��t�*@1B /�C��c?���.Wk�Hi���i�ޠ:�j	�H2���N�hA��c�*z7�F�uX�1��/�Qx�Xʆ�4鬿7_��\�蹜0�]��؏�=�2�X1�O����J�H����	��������A��)i6�V.r�̚��Z� �����o�~�(,���>bW�۲�V�s�^��fy%|����
�1���4�_��wb�b���ͯ�8�d�~ﾷ��e��31n������q����!�&ΔɓC]��Jvf)�+˙��"h,�S�DTWp{)�=T1]�u1>?C���g���8a��_^�)0I�a���2m +L�&�����^
0$M����=P-��\"]n_�ɹwP��:bw*�A,Ȃ��dg�=���{���g!��������L��.sW���+c��/���T�I�c؁?��9'⋢.�"u�f���&��T�ׇ�Q��e��q'h���B������g�������r�X'-��Sü5f+�1�ʭ�B�����+��@����Q-1�cP�^6��Y��7�6hdr��%b|�`�O����ӏ~;�\�.�9�ظ����!��ǝJ�E���N3�+iQ9g&=�4��]�uH!�[�@�ƙ�q�%w6� �A�Y{m�ZHtI�1���:Z�K��khU���(f��Ƴ�i����\��ډlN��1e  �WXHM�n�x����&R�,h܉A��n���q �a�ß�c��qYց��OT��ױ��2��5���\#[�1Br>'�fA�B�%��z�8 �����ѹ!C.
����ئ�b�-����:����~bs��������z����C�9��#ͿІ?])�h�'KC٤~��r/@n}�+����������Z�ѕr*���kr�>�ǁ̍D��27b�'�祹�a��4����6��sz��$i�����r�8�y�C7<D� ���Lܠ��A�bAv���{XC�d�\iQ�*�B�ȇm�V'�V�q���S�.��U=�����S���럙g�D�Ԩ�ވF����_B���1'+1���B�?O�@���aמ�jc(�]�~��w�@o��H"b+e h���/��� p'�K���fZ{m�Bg���n�P������}Tn��y�Cض{ Zx�
�s�u�C�TW(���}ϖ�X;K�&t?ͥ6Är�1��w�!���2E其���N��������@J=�$%f$������"�/�M��Rrf���i#2�����Z;�N{�#�;;ߧ]�������MK,}LS�Co��+Gؖ��@gH���~�Y)#{�9�)B�r=͛��ǽ�@0dЄQ ��^H�,�	?xdw+S�ȗ-��k6_2�m]yƍ����T�]�Ҭ0��C����+vw��(V���}';86K�� �c�g��@�.Ч.��_��6=�>^GbǪ`z�Q�����7���8w�k]S�����; ��.��{G��Nkuot�.-2���j4Q��.�����M�#:F�@=x����%��S�3K��N��w�J)��W�R��_�I��B؛��端q��Ea��=gZ�2�	G�a�%��p��p��Q��Y7;|��2��@������8iR�/Ȼh��Ϊ�D<�A���F��m'=�N�ط��n#��2�H�tG��B��Gk�u\FQ�'�|�Q"�%���&W��d��d�ET�m3�sG�ؼ~]k�;B�%s�m�o��1���,�_zI�gڕy�3-�G=���%߄��	i^,�ܶ�F��'���t O��e���ގwʖ��ʵOP@ce�f�y�He��F�ʅ掇���k5�H�I�M�r��j�¨v9A{�v�w�$��x����_��Y�i 	g�h����f�p���X��B�*�����?������0��gm崴�����G��E~a�3X܌S���hӥ��{B�Ujm��yL�C���F����]�Jrӄ����M~s�iK�y��}���堳a�W�y��(����%�iQ	�6]9��EÒ�q��5W�PÙgb&�L�h�q�B���Ql�0�n%�R.� ��JBܕ|iD�X������B�)�h�r._V���ro~+�2}�1�cpBy�#���1������o�������쳸޲Go6L'*��BP��:Ay��C�}��ũD#�?v�$.Βl�y>v���AQd��f�&�l����'9��Dt��
�3_�	I�Gh~��7��D��� 
{3$V����b"�6�������:�I�e#�')X}r� �����%>�a�%��
pi��I�����
�u�������G��.~�bUHw�'ʮ�>{��4���k�$e�0�V�i	0v�o!4�������On����_��;����/Ϣ
hQ�..�c��镎��q�[Լ��y#of^+����G񃒷T?�-������m=��d�J�p�꯳�'�3�A��R�eP��Y�r�����Y��V��zp�!֮��S���
{o^�����a3�oa���:(<�l$e]�c�Q�S��$�D�Z�O�l���H=��dw�cV�\���E*�?N��]�q�b��I֎�y�5�5���*Ќ�å(�� y-f2��(�f	v��_L��b��P��NCfu��D�3q�vkV�*�ӕ�5�
�X� l&B�fh�k�L��$0� D�b�z+�M^w�u�����PG1	���j�+`�SK���􉽞��썗�̫�n+w����tn�d\	�y�������aŨc/G5�	�����Q[/�z:p4&?p��/P"�]0'&7��w#M{�}������h�A([�G˶����Ț�� S�8b��������Z��l�� �J�<��D��F'!K���>��1%H���E��~����c��W�7�\������^`s]���Ƶ
��y=Z�R'�2���	�Ȍ��mh4.t@�*,�S+>����̗[�e�K��/���� �&W��L9�g�a�PuL{��M<?�ڦ���U5������]R���[�����̂b�� _A��_.����Q3��l�Xm�ي؆I��Q�Q�f!>�5��[J�:Cn:K1Š:��ʧ�6�7��o��Zĩi��W��BZ��*1�6N�Mo7�-rx׏NLD�Ն����#)���)���E�H�֑�GLV<FY�io���O0�C�ܮ���x`O�8��1|��#n�HF)�ͻ������-�������T�Db��I	�3׹�_¼�!B,/���A�����uوF��zvk܀�B��:�W�I(����T���>׸�.�!��_� ��n��t�����q�Nzf�z������Į���a=�<p�5NF�磸����̾E���V�j�\S3�{zDl�d�~z��=z?�&o �m��iR]<�b�V�_JR2��FI�ΛmQ�~�6~J�3���,{�,�2����ͺ~-Jƶ����W��+� {+�Kأg�QM����w����y}�9���ِ�%o���˳<OG r&p�l����Vn��)�C|�R^<�i��V����mA��t��� �3�ĺHS�g {�uO�;��Q?3,`Q�[~�� 'V��s��V�"�K�{l�XuA'5���Cun	�MW�|#W���s�o����p�U�1����P��C�zscM��Xr;����s���UD�7�E�=؈ \܁�`�5�)�`iԞ�F��C�l��"-J���)��V�?���p#9�ݜD 8���3����貧��%��v��#���ף4 �V�� r�;W}9�6z�m Wx�MR���q�|�1\h�����aA%�]�9^J���]�ǀ��"Z!Ī��y& ��]���XGW�˒\W���^"����ɢ�<�1 ��{�M��8ب��(c�ν����!b]���z��#쯘�G�U$j�x8-2�;1���}���Ƃ|yPX:-��c#���GoC�������.��h]���NM�}�Zz*��t�?���W��T<Ɩ+rat��]H|d�[8��*�X<��vs�yO�퍃m�[���q+�}��0�[�'��(���W�Z�L�c,� �>Q��(-^�u�䁏ӹ�c�h�qy��0bN=NJ�\6N%���1�pw9qPs�\���|-ɋK���,wP�
%5B�3�Vm�+�N��l��KF0	"��e��}P�#���j���فT�4s#�Nȼ�[�'wR`^�~��G﹑w*Dρ��gfI/��D�-��(�X��9�~���#����l�������c6�(�R�����N�����0؝ i[�E���Fv�%�S�̉����<�停��=�O��8���x<~6��v�V���H��VQ��\�׋Y/�T;E��͢�$��h/�_��0��+��Q���oį�����$k�5U��*k�+ ���Gip�{��!���Ű`��l��jx��x�OfX�����^�9BK��ʠ�b��C��9�4b��aOUǆ���<�?�>gk���khO�A!Sw��
?m�=(e.�uuMqդQ����~ڥ6�����-r�J%)���pX��9��d��7��қ(z	Ѵw�Zլu�~j>�g!;;�g����P�-@���|����-J^T��Osj8g��v�|CdZe8�ǋ��,�(܈�h��H<�o�����T���T1;"C�
}�Z��s۟h��cîc�MY�Z�bm�J���,D��e�b4>�+��]�+�=l�Xu&�b�eO8F*�m�������;B�;yPJ�4܏u7�͆�.EC���Es��Z�0��r;��t�z��R�hh�诨� 9�h�����*�u�����%����0q#�ykk�Ux=�a�s��;��_����Sp78��8О4i�&����h��+n��ó�t	G��y�P�t/���7t:�u$F�j��#�y�V�f�.���-�s��ɉK�
�]��%�
�[bZ/,�z����Dv.^�S�z|!{w������UAE�P�VU�i��7��QU�[��i�z6
�m�j��g�}G���Ɲ~��3��yf4� �c_ա5�fU�W>S۠h6�R��C>}a��ޗc����KGwH^����J���[�M&��j��W�C�R�+L�}�͙�����jj���
��l�K��������~�1?9��
.)4 �T��:f��Ŋ��u�^����ӖQ0=4�o*�Z��0kHuP��1��(�n��>�� D�x(�L��&�z������z�xo���AV��'R�ä5���A�=5�L���(P^�?ܑf���w���� �4BC��'�B|�R����K�g�.U�w9�p͚�����g.�����@�u�]�jڭ��x�fjy��F�C^;{�_�k>��*�����q����;W�ڏ�+��a�n4��)k�I�&T:�F�oˀ�{�����C�Z:}ŶxB��o�X��V=���}�܅_c�.H���RG*	T[h֓(��)B�\vh�a
U��0��SO͎N��3a����+m��˱ ��,�jH�n���m V��c��5��H3��bD���In���|W���6W��&Vz!�"�⪓�d[f�oV�.�?�7�6�8h��R&eU�
B<$9a��A0s<���6�5����}7B�������\�8}e�Pm(�eB�ĥĀ�����(U&zಐ���e �65�r[%�!'�Q<X�#tn�����"��Z�s�W�ړAԀ%�>JZka��:���T��~;rpt5�M\9�i4y���]F��r������;�|���V��g��T��8ԡ4�f;X��hׄ�bY�w�R��9<a�����J���0���g730NX=�OM�٘ �g�:f"�ٓ��Efo+t��Jg`C��4=>���*}�*c:�#z�n�rt����]Y�dQB�%&X��t��CjQ[�[H].���B��V���Hk��0��;��J(�q ��f&�Y���H�#�i�IR�	�<���N^ �j0�!W�r�Y2P�y�b��6�T�3��mޜn'Ji��f�B�p��m�i�q��J�Q��!V�Cr�����L֐/t��ʫ�aw
�vK}��N�+t]���9z��+Js%�U%т�j���phܓ��}c�����D�^$=%�N�q��/5,�sM�v�k2��{��λz�n��czs����,�P�l���� ��49vU��Q���	J��,�9�v�E���vo�{����,`�`���Q��^� \�/K?�+Ǥ(���<�.��8�V��a�S:W����Y�\2������8���MW��6���O�pm<C��/�y����O�i��V/�	P\-�	^=cSC��g��v��x f�v���w~���5��R�I��G(5~�	1�=�b�3�#@��?A��N��{$�=�o�\N".o�Q]���]5QhSsB����Ɖ	�j���Q�*�sB����$��Z�{]y�b�'ژ���w�K0��,�V
|�.1�����W]�kp�v����S�pbܔ٦Ë�6�4F�8�!̀�ˉ0"
�@�s0Z����}�0Ȋn��#
�X��)��'M���Z���uk�6
��z�!�>w�f	$���*0s�u���i����4l��Gg�ݲ��c,��*LI-ϡ��m��!���хL��CTy�\�|>��:|�4ULy�w^6�6�DO�K��X˴������mT�� �����P�H_�-�3;��V��A6��ؽ�5�e(���b-z�N���(A''*��)	�)AFb�Y<�����~�;��B�-C��K$S�4�A��#P��C�h����Ϣ��h.#��d�)�ĭ���N�ѧ�7�!�:ܝ���ڭ��1���Ƈ	F�����D��@�x��k����Q�Y�a�Ǿ�\�	�}�֕�4EL�ɝ7���?Ƅ�����R�T�q ��u��,�����یr"T.�x�# ��6���b7�4F��� ��t8�����f���hh#�:Y�!ϝꅻ��7&�
#��+��, S�~n�<��fN�dhZ��>4/��] �ׇ����u��[����5�aj��d�ϝ� � �]zC�P>P����_w���� �I����_L֬�J�NO;�ْ��a�"\�NflYk,c�Q�q,J�ZX\B�������:κ����Q�LWƔ���@.�d�	�^}0�'r�X��v����`�܅xnH]�j�_�<�a�f<Ꭱ>�ѳ�?Zסc�]˲�;���|fg�9��4�ЪkK�|ѻ�W�#]V$�K�,�C�0o��sq�n6~?������ [_~���g�\>9�q�R�<X[��#��Y�2�y��uV#Ea���Ã_�l��Jp��0��lܜ�:/;�G#QK�u��r��I����7��9� ��Q���gw��*H��e��-��ʵ|O��"ދB�4��&�pZ 9/�[�)�N�]������k��,;�9�����u���(O�/a�}+we�Һ^����Q��L'�T�bg�
b$�S\��a�x�Xf@��|w"*FO�&����/%�-�n��3�ߋ�����f�xW���q󔮪�7�Ąk����e2��swf��Ѩ��#�6�:�͑�)���g�{*U�3bW���a=3f�� �[�HšU���Y5�9Lu�p�"E��X�l]�M�s&An�"~3{Bn8�dT��Q\�+����Ye�yIp�*>p�Jbܫ;y���i�g<���'xkr�߈��wPz]	UC'��/z[��g�ǟh���=:T����9�GtP/"�Cn31Z�9%�I�~�/9>�7p�����5��{1ȇ+���"�!g�\���J��T��H�p�����Y^�?���K�ly20��|_�)�S)�zr�@���r��U�����X��?�L+CX]�E�H����Ʒ�:9 0f� �
��L�b���F~��e�+Atl�ܿ�����v���]�EQ,�q0(�K�R����Nuٱ����-=����B����#J�,bp?�n=�����D�Л�`סîK��ҷQ�[�n�c!Q�P׭T�{6�� ��^i���2XC�к`�U�B��u�1�g�:�b��KUC��6�
q�[1Ԯ=Vf~��N-z 4P��-wc��!G>��@�qW�F#>�=	��v�0E�9/��]`��`S8�'�6P^���<�P��=�T����܀Zh��6�ER��j�w�k�>��"2�yc�/f�|A���{ӟ�`���0�,��d��J[>��ڏ�7���$�����L��Bl��Wmbz����畵#��ٌa�	�Jn֣� �lb�ui�r���ɰ}�~.���W��T riBn��\|�&�(P�/(aH��Tr�`�W��B�'>v��r圎��D�hw��p"����4�l�qaPk�;Krn_����k'��x�F,����.��Һ6�W:�~0��,�i��VAG�9���w�+{�Xp{�&���{:6�F{�7A�U�����Z�����WɆ��&B���RvBxc�d7ʲ�Th6�%��a��e*Vrlv�U?*�G� xx#��	�QN�n���F���:�^��j'�z���yy�bi�]%Brſ;T�k��5@��d���A�S�5����sJH!7�J"����g��ƿ����@��#��������0T�
��LK9�$DN k޺�����������b���U�d���AgJ*��z�Z.i�%v�����r�p�@*�ES��u�����e�]�eIw�A��1"�:��JUrg:�	|�y!�"c�U����<�VBR�5����%�A��J;a����Kпqjx�z7O#�O����*��_���l�P(�g�I���1�^�� Gj*�������w>�B�@P�(X�R��J�����}_C����M@���;�� �P����������$�>TI����Q�M��( ��]h��b(1 �ax���,�@��졥7�h���?s�u3�s�P��&���+��v"��C��p���p91r~Ʀ@b�u�ߖ���J��hlg�!��M����!M�A��}"h�t�ߌC��Bo�"&��'��1��(����vH�Lݑd��Km��|��נ[��u!5���K�&DY�}�	��#�(u��C�*��nL���Cj6���c�!�8�IR��|hOţ[��[��
R�V���-c�ߓ�.�Z`�;����
;=ZG�S�(q��`� ������K������#0L�pq��k�@���A�ς�B�fn�F�]�3gh�8>�[8��<z����Q�.�u��t�f/}g�$ҩ��Zh���d#ԐM��Iabp����.~]2�� �>�@X�����eKB��BH�N�N��� l���G-�*?
��l�	���~�0��z͵�+�f,���6�[����*��Rq�����cC�Do�f��R���i�N�٘��+`��Å{��k��]w��j �'��X����`)��h֨9ώ���$��m���g��~�Ξi�wJ���J[�<�"AIDc����?Y��Ie{��%�&B�mW���a�/?SԩL�,�����/q˩!�xV\�/j��P����:��P?�rIz�U����w):&�5��
��G�����@�n��$�wb�"'�4Yp��;M��Sdml��V؜�������T�C�/��3p�q�
w��Yp��X��Y����Gq�@�/=]xZ�����"m:w�57�t`?�D׮�D�$�4lT:�H]��S��[{�-?$*���p+���6,2}��'Qގ�gk�9	��M����s��No��L��*�8��8����~�I�I�C�>!`W�wՊ���*�}j����?�Z�ndSq��Hev�ulǼ?�}�`�{�P�	�zY+ۀ���ؽ����%Wk
����Z:(l���dá0�1i�&Ҡ卜�u�Vo��>������a�l��������yC�L�ߧ�����~�VV�X��زyGג�p�_;��7m�a�L�6�yS>�v�^����y_���ྂ]'޺^aUY�q��U۶bG.�
���b�C�-:#z\�n"2�z�<S���T��U�Z��;�w�l+��"xFk��(qh||I���C)�oƸC#?��!z�~>�9���\C���sR��[��<���9���pϖ���en+I-�o�9L���A(]�V���koh�Ґ�;M<S�����ȭ.8*�����=�}]6�4��Ge[R{��s9�t���t�c�M?�1g%����O'8�P9W)��~���P��a�:ujP�����l�����U��),�:z	
boz���雪g�J�
�
横�{�j�[MT?���TY��Dk%�Sc���c(0����)[f��/{��9,\��.,�jb*��#r�K���Ok�uD��J���{Ŕ��h/�N���#7�"��^� Ձ=	,��>H�	�]ݻJ)���o���"�����%�6�1g�t�.�������~������T�����7�����"��dh�~	6��fg���L�J��Ku
1kˋ��ZW��h�,;����<d	�����?$��γ�VUlf�V%_Oܞ�9��Ie�54U�.u��jh��j}c*k��bM��V�8��z�k^9�u�H_XX"=�h1���Hu��2n�f�.�F��$U��V��N�Y+�6�C��(U�؇�T ��x\����R�B�?"��R
e����:��q��~���y����[m9��}�(R��%P�ڕ:,�6�?�<�ƔPNnh��>�ѝt�Ƿ~��k�
��n0g�GVA�/��ZWP�*8�|`&�C/`�%7���ה#k�x���:M��Ծkd�ތ3!�5��L�h�Edx�*m0��g1���?ɶ¹�d�O,���ӧ���B�Z�@ӣ�L9��,����