��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v����aW����8�]�T�]�6:v�&�CMl�g�x�J����l���WP�C8Q�����
��1wcf�H�Ĺ��.���I���v������> B�G��3�2Çb�ZS<a�M�b���>�tE�f��ԏh�����b7 Ql��~�^��_�XO.�`S~��x4�V�So`d3�O2)4I�ܪM�SD����w��U��%+�:h��:�1��d�Ͷ,�0�i� ����/�	 ��0K-O����2�}�V�����Rkp�r���� e]s�"���lZ��9������55����.(�̸�)墀#�Ľ t1��;���8��1���$�F�"��>��|��wS&U0�:��	�Z$�n��~���|x����g��$Ҟmk4j��B+'�N[c#n�*����?d�
kWm"��q
�cH��8�r�>t8�-�Ui���nEʗ#P
�p<?Ӧ��,�C�	ٹ�]��|�����Px��Xd���F2̡H0$c�뮷�ō�Uc�Kc���)P2Bv�"��
!D7׀��C�v޼��ǔS��4W�E��XB!�1��E6�CP|W&���A��4B��,�7�P&|]+�ٗ��!��7[�Ǩ���-N��@���{�A���З���[�T�PLjo��W�|,���<��s2(-#En�� .h�V��ǊO�<�Ҵn֒h�G�s�*��5[h_z�\��@�Y�
�)�z�z�t�2�K���M��fTT(��|8���O �|�EA��u~�E;���J����n�Rs����y�ɻ��.�I��: b���<�,��*~h(�u��.���)QI_�Hg�7sj�UU�5s�q���5��B�����14���ԟ�6����|�0|W��bt]��=�w8�����/k~�=�{�t=��O��dh�SL ��7D�k$�T$pk��H��o��a�g�V��U����qp|�a�iP�d h�ޏ�s(�W"���o'=�ƸĚi�4^����d��?���I֗��a;N��|��_,`�����#��d4jau!�����uh�Z���±�^z_���W|?B�a�s/ �ȫR0�M9���S���R�<ʽ�ݡ#�W�I�nԜ=��Pn�>Z�",7��a�]� r��8��	�?��糟>���"���)(;����w���Zxɪרl�M]�\x�"w�%q�2V�HU�~�dAf�m�$>���z���X�4����S�{��U�ܗb�m:D��L͎���-��y�?D�dR��|��x~%Z��Е��D�=J�ߛ��b��6.�F3�J �T�V�_!�n.�b�Q�B}Y���Y.���e�\�C�@��+�� ��'�9�vŔ�������\�1�K��X�4^1	�d3l?�N���u�G ��/Pq�g���؎":��棶���p��~��-j�|ԫw}B0å�������K�e�T��<h��&ӗ���h�v�@]E�~�/��a��?������a"���]�ȍ�h��$�?S���ů�D���0�\�%�T6���ιޮ̢�Ǝ$��ԭ�c*\WX9�;��7hNvD������Uu�����`�H.e�&��}H�W��k��;����xSw������>]��-q ���s�ȰH��3�3'T���r��|�(2ϕO�~Ă	�2|�w��@�I�<_H�͙,��ʏ�� R���DFeDe��Lyr�i�u�k����8.��6snz0�#�cI�����^M:��iʐj}q%�����m�������<�4�c�a 
��-����(Tנ7�S��Cg��vR *�r�[R�i ]^�"���ێ�30�!ɨ���[����.��Lt]g!���,���*����ěxq���F�V���$y"?�����P-J�=臼#I��Z�y}�jY�����l�R��j���_}>T�$?�?����{�J�U84��Xw=���R_s��D��e6�g`��v��ch�F�U��ZR@x��>%��`���Fǁ�A��ꟲ�b3���2��R���+�w��u��v&�CF���R�Ҫ�c��H���h��ـ��xj����T�������+jy�#�����8!K.�&�U��9C
F��g�T9y�c��6�ǋyMF��܆��d�ha̼a��H_�m���z)�l�!����(����҄�R_D���Ե�4O�p�w6�Hq�αʾ���)A��h1<ƫ�Ay�U��tJ��f"�k�fa�M"�SkVL&ɇk"|.�o!]BV}e2j�T�2���AC@e���F	{&��A�uv�>�W!ֺJ�ߑ>�	����S�%1��l�xG�s ��a���3q����&�W9]R���\�}�n՗�V)���-�ؚ��h�T��W7���yKv����~Y�:vY[aV.��|f�2%��f�ڗ��߰��U������4����%3[.PH��n�
�=6��xZ� �Kp����Y�v��ʜo�;�pD�_��5E/ �^&��� &���]l���g]HA��^���}$]8�]�� �Y�)v�R���S�Ҽ��}���3����ɯ�߽�A�s��s��2K�П{�8���pS��pB���A=VɢX�U��H�}&�Y��Rb,�I�� ��`Nf`����R��"�IJҊr��{��}��T��/<m��(����[�x�W�0���r�Y[?���������1ѳ��H�#ǲ]�w@㯲Cá�-x�ِ�����M�7?���
p���;�9��O������/e�J�[���D���)�Ԕ7�"�}v�1阚'R�nvؔ�`��HEP�!MN9��S)�O�s�B��`����s��ث��hc�"]h@[_�������m઩�r�
�P13t��P3�h�bI��{ 3���uq�ǫ;&'��$u��٥^)��S��V݄�����{$W���
=eF��a����@�c:/z68[]�h'&!Y˝���}O�4~X&��#z7�6�E�ħ���iAV�Z�_�VZ�GFf�K�F�Y��a�o����[����;��v
�������ar2���[�]�/���'o{g�ח������C���)������GG+*g$��0�A2	'^�\�E3d?��'J����M�<$�pfҠ�VG�$T�GW�����x8��m&ط�q%ugL:<�ɇ?BixN��������^E'�����"z�^��@��Lΰ����jBW+"��Q���S�Z�)����x�8�|:�#~��D�:n��
�{/�
->* �F8JIe2�����ޭ�s�.��
t�J�Lڒ��!�x�?x��z��e>9���G�$ѹ� W�D2�sl�<���Gw� �Ľ\!=⃧Z��l9��#��,��4�U�,�SEV�eó��a����w�t�I��&�h���E��-���'L���U�8P[MU|���DFE�_f믤d"�#�)��9r>y �'�}gOB�=s�r�0'�)MwB3�C{M������(�Q+�o(mW9��p&x��Gu5O��Ϸ��^/	�,C���IH��"�gA��KȊ9�-T