��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�xX�GPW��si���骿5�շ��3��\o����u�.n�Cez!�������8�s���&Ĳ��<A3����֛W1�<m�7�p��ۛi��*7q+�/	�:q�F=�@�_ڟ�]%�.���]A��>�-�X��;�W)"��uƬ�l͕�e6��m��T�����1�Fٛ����&s�t�\!��2�9��͐~@އ�S��,D&yA��/��!�͟���ii�ߝ|��%T6�}���^��n��8n�\tΪ7�뙳�3�w̍�hэ����WO-�X)�ʻ��%�D�[�xlwu�C���O"�� ����:�|A9��5H�ߗ�~N�J��Cz"۞��
��1�(#�d��C����c��y����j��-e>m�~��Ϛz�1Zh�y/�D�%W�߶1���rG$�ogqh�#kv.�Ϧ��)���ĸ%+d�Q�lL�+��k��R�a�����7���J>�h�������������o���<�	�l+�x^��L���қ���ĝ�s�!���~*�Χf1@��Y�@�->�d��@H�������o�Bz:�-RNmT��JcH��u��(QA�.�V�P��a]������,
�#�p܉�.=�*`s�����}P'҂3����iu�d���LOI6�EKz�d���pC,vY`��A<��P�È^�w#U�%/�'c��\{��hu|n	�Z;�D���9��z�z�,Ch���V�q���h�{�w.݌~�����n��@:�=�tid��ޏys쇴K;H�[�<�e-�9��P�nn�/�E���_�`=�j�e��@�iw-
U1�q��gJ�UT�\+��(T�Tލv���*���5�,����$�^GP�Z@8R��W���n��K��F-��
%�^
v�<��u0���7W�suD���>x��G�t.N,�MZ��pw��@	dy;�0h2 �eC�:}�U���]\�ߩ���]���-�HԦ�T�̿�R�b�R�h���D=	dm�/��w����I><��*ef0�'Z�3-�w�'�J�U��z<���\���Ŀ3�!Ri��GZ�#��9$��\2��n�[���P�u'��1�B��ޠʲ�V���L�tN<�U<�ZA����D��8atq���$p-G�0���ϨHN�h (��F�mTM�yc�����P�HGK��������0�P���q��/�j��L�a���r�BK��:sw�Ɲ� }����#a��~K��	�1�$;,����ڙ�,5t��B?�T�������f���I���?�~�o�$K4���@�X4K�$�1�D�e�cM����q���G��T7�-�lZ>��J�s�&�����
EA�.S5�{�5]��yN��Lto}��ܫƄ�� %�uH����G�4�{�7�ہ��V�>^��Y�2��d757mbgOY��d��r�����Lf7��h�����?�hLe9�>���m�w�csjAI���or��Ь-Oа�z�l�W�a��}�yh}q��b&5���u��p��E�mpiFL�  X[�WJ����I|�o ��L Rݒx0aw��j[%I��:C�P��b9��뉱�R��x��2��q�M7���k�h��fN���J�se@'cn��G���
xͱn�!��t�"��ҡ�#/ئ?G�/):�I�Y��܇c�˰m��TT��`q\>ʒ�e�����ߓ��'	ݩmE��!e̻i����c���p��-_���:�)0��\LW�,X��ގ}-r�.����m4�*�hi/�eF'n��'�wr���ȏA�l
<�ǠoX+�
�k�)_V8j~n�o�ᙶu\�b��7~����� ZB�Y=a������v�r����/�@l&�ʓ�� K�ZZ�êo��z؎g6�����Ӽ�$�8,±q������
�+������/�����٘�W��Ƶz�DHkc?�`ΕHk:��bb��;��8\�[�J ���Dޔ/ �!Y�X���[^0`O�t���N�@>T��A���?��Y��lc	"9FP�N�e�f<Qo�8���!٣��D9�RM��'e	I��?Dp���122#(Leec�o��eJ$���(D:����?��H��i��(;�2��-����!*�n+�k��Lՠ}"ŷ�����ݖp��n�+%{�>�Y�ww��dL��6�\��D��5����`,���u2�yr~:!|�W!�,K843���	_�ӝK����l�ɮw�	�根��޴���k]�.S�����7���������c� ��A.Z��Ay��Fإm� �ᑷ��YԹ���$x���U�*3%�����0]`x3���8V�:�Ǝ�aAF(o�����d��7.C�/���r���b��.�]�NY�ҵ1ӻ/h��afZR�k�o��{פ�UyQj�T2L8y�*�0�QsU��^��Ԯ=�Xo)�|�X}�fS�Ƴ�\E$e��t�&�� {�]c��p*R*Z��� Wݪ�==�Oi��Tƚs��Ͻ8�1�9��N�(O+�GA@�8�����:�b ��$"�aA�b��U�����<<��$_s�=c2=`�r��C�S�-�H�O����rmZ'��pI5��u�(�C��2W��6�jqCi�n�W��e�P�N:ST�l�b|����oS�(⭵_5�H�e��U��u�.��_�kܬ.�{�}����`X��[��$\�B��d����1;U�����t��S#���~�<��É�L�w�6}�=aY�c�m��wS��N��\���m��s�����?dP��1�]����%~��,�����O1��oO����>R];y�=Lu�[�������T�"�4�#�+	ݕ�y��]�>���Z--�_,7�X��Ο���������l<n}��X&QlH��~����[Ab��[�GE�Oht��U��(2�8L��ĝ��f �4��i�`r)���_�a�ڌ >�����.�)�v�Y��'�`��{O�i���.܂���"'�b��HP�ӕ���%�}v�7i�L����9Y"�u�%���TcvȼM3��F&�Vc�ߡfN%0�(��Lv�kwk��R��͞�&qH��2o�4AL�
 X��m��s��|��E�H ��Ӧ��ȸ�1��d��3/�[b�[�e32���f}ڎ�2��/[>�q׽�snNq]�T��q�1����9y�z�Fh��E���fEJ�ؕ'�L$��Km8��P1_n�I�+�N?6^*�L]ow�9�k�^핎v!i_�.��V����)�\����]AQ�CX�~U;��$I����/�ܬd�R|��-���U����AF�K�lR���5D������k��2^�T%�2Ij.����m6ہq�w�C�F�3��ia_:8�Q7�'��&m��!�,�,���-�[6Q�"�dSef�7����<�?�@t ����g��;vU�"�����_�w����k<��ih5pfL7��O�Y�P�f������M����桽_	���@#�YHǔ�~<$���uV<�0�rQļ�Csc�9������IY�6`�ĩq��&��Q)ߞ��A�Y���jyy����f���شHv�=���ؘ7H85ը5��zs|���2��W����(��?�9�U�����~żP���_\YRv��P�#���s|�YHf���Nu��`�~��zjw��똦Ac��k�҉�����C�W&P�'P5�o}#�D���?�~����Ñӌ�X53x��AX`���َ�����A��=��J�>����Y��2�P�F�s�)]��`ec�_(�/�0eO7?;�i��#qJ�_E���>M�g�6�^6nzgaf>�9e�}04���`��J��ɄL�~,h�}n����q*#<O\p��E�^���r|�7�& ���Əd46�n���Z��|�*����$	� �dnn:V����]1�ŵ�fà�<�DH�NQ�m��(T����Ք�iG'QW���K���
�h��bh�g?�-�Sh@�����|���e�����o�3�%.�2�ꉑ+5;v�����_m���7-��$�sl��+i`�b
�L3���_��o�U��t�V�puFT�<�z��T&+�w ��ԗsH�,I�Q|[���!�e(<R�I�9��.Jd��?�H?C��J2E��m8"��{���,�!a�Џ��I����SӴ�ZXr��i[7��x٥��Mɇ�1�7����<v�g�rQ��a�k,VA�\�r���,2z;r��?��9�9�F>Av�I�R�^���XO���st��5������P�S1i����h����
��c��B���{�����Α:E�������8Y���:�u�����65��k�Ȅ��<�d��+��ۖ���&��v����9v��n�O%��9b�C�������6�������P�jL^5Mq�������4��c���KW�9�����W�ZdS�?zu��<�%�_�R�!�p�ĥ/�����6j������3ԛ_�,0���-������d�K�'\{uu^�T6�l��l�&H��Û6>P w��~.���x!�%�'҄��7����2RAS�'���p�����c`���GK耽����@����_$�
�,�9�0�$�3�zcs]��q�[�UR�#����ts�	��ԵJ�I��V~e�A�����f�A�;�C(e&v���5����Hó\8;��:g�+��7e�y_~����H����AT��y�.�i�����#��&v�
�j�^���b
,$��*�*,�r��rǺ��ӬAp`�-�hQ��Q��5������8V<���y�%�gZ��<���R��9ԑ7�n1�&l���4��;�"0ؘy� 9�
����̎(��C	Րnb�'��/װǣ� ҷ̆ب+�Z�-�@$x�I��(�D���|���I��BK��5v�F����:+��+��=�G�G�jK'3�9�\A���P��2���)bNVrHA0�%�s�s�ր4����� �{_8�9E�[�f�u!{L�/�6K�q�� �����W��=� b�,�M���,���7� �"<2�P���_���h�O�g����|�^~8$��挰�73*V��� >D@Up��gBѮT�����Q�X�x�Qю����3^��	L߇�=�]i5��˥�U���g=;f�����uT��A�;հw��R�_�:��lo�5�90�7�O��Ժڍ�kkq�~Q������ �B��$p���^�~�����tu�N���+�߉��Tʪ����y/�"����0�Mȋ~���I�o)�S�d��$� �d�䡡�>���c�����x�4ъo���~PR�2!H
�8�S����t�6��z�+w�4"��~�(�d����~b���8���u��?Ϻ���-��M��z��ZO��xN[cA5�,�ޑ>yc�{\��N���u��4G�@�.>���g]P:�|<�^�
"�AA@�X�u�Xڻ�5�/�7�S������|��[1qBP����Pa�ܣT�L�ѭXWxu(�]@��5
�A-�I�vG������֯��8�������ko�S.@gۗy�4�b�Y��� �`rg�d�5Y�Pa��R��L#̷�cw����NTNa�\#ioe�"9�uZ�<ۤpu���~��|�P�l����O9<٪HjôL�1ۡ,XR����?;�+`�n��S�a2"���Q1�6��g�1P���i��|xn���ɱKC�1��ʹ��h���<��o�I�/�3��[ ��^�0�4�"��8�d�Jj��<��ir(|h�%[��|C�(}�6�a��l��h��|�Y�¸�;�
��kL��1ΐ�d�M�zv�A�n/�B�mQ5i��vA[X���D&��?�(b�m1}KG��>��F[�Ē�X��>�������h�[j�,	�L�U�z;�K�wɪ>{��:&�V^��_��巊&�U-�
l�ش��`|d��*��V�Ԇ��˯(w�L���O[7~�87�}���aǆ���K냩�[��������P��5+��g�f��g���f����pn�q�'55�疃b.�E�0�os��c���~�pFB���c^�r����;bIA�᮲q{�����Î����ut�X|a�==`�i2G��E<������p�o�i�+�3���[��z�����0�δI9��'�s����-4�_%9Os?#q٠}?�2`�����\�oq���.���6�",z��x�ض�r�W���(n�����6'�n�W�\�'�^��)�d@��5mG���@S�5۾���O���{�+Ζ'lب� ��;�E`���u'9�3�`��-}�ie� +Ye��M�&�Em�h�T^ۗ�b�WW�8-�1l��6��zN���n���f�BI+��엔����Ycz�i�%��o1�yp��B97w-��^okkVY�<b!��������� ��'8�S0���|��ϐ��y^������#�v��/ZE��q�P��2D4�1X���mM!�4�/w�R'��8s���"��,u3EK��Vn`���j��T�9E�z���|ծ� ����a�RV�>;�8�fa7Xj���N����`6$���C�0^���<��⻼[W�!ϑ�>mn�^)z��/�Ӓj$��j
�D�z���q��>�Vx�D���n�U�'�1���Ǣ��3ď��7v�֧�q����n��2�'�)�6yp� +_�VS�>K1��g�9�9�'W[Σ�?o��.䶽bF�7M�k�i=QaD����r�6��) #��P�T�w:�W�`V��'>�tG�.�>�N6m	7F����D(��e5m��1��76���dR�W����	���У�d+��w1�>Y����&��6II��K=F���$�m��I:�M�J�M�ͷ ��T�����*��suVB��B�M8�@�1XY@�:�R��A�@��a`%�/��#�6���Aw�}� $���q�}�ދ�R�5�~4��a��9�q=�o���\�C�b��dC���9<ՒO��j�\��p�Y�,Ю�a��K���p����Q�B�5mo �_^��h3-dc3g�_O���R���5�QyN�����)U����m�C��鴕����3��ȶ�a]�[�M"��$������y�K��V_��T��+�{�{���0��q���3�ϪF��u^p�8ݫ��o����� 2������������7��~�=���<�r��1���mmA`��B#�?��a$��}�p
X@�I~���*UG$�6��Wjo7]��嗈����jM\��F7s�Jƅ�ѸcIh��*�:��&ξ��e/`��z���&j��&]�"�-�ve����_���X��Nl��@E��3�t���p��>�7��ځ�����ԂB�Q�3#?%:,�V���k���ۍ�-Cֺ��[34�<4�!@��v�kH� �=u�)F'�J�}�G9ԫ�_��=�3k��Ş�#��E��R�'&�ڽ1��̙����5�'�ӭ�'Yi&5�SG�dc|&vYƋn����x�N�N\Ç�c���