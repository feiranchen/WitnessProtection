��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX� ��V��P�����q�G}�~��a���[ۻ�'��0B�
��d���d�a���Uc7eN��������#夯b�������W�D\V�L�̅�/wO:�jdmY؃ơ�Խ��Ӥ�L��Eğ���'����yY��7s�F����~��(����.%�Q��u8��wW�[00/�[!�6َ��t+|��X�#2{9�ǿ���k�-����i���dx�#�Ҵ*�'���ҫ���/�#J7����ru|"V"����}yj�J�{�㧒>�v���D�D^�h7��]M�GW��ug������imӑh�O�Z�TGi�a�|k��z]�Ry�>�״��(�mD�Hʺ5�[���>>�.���u�4xu9�<��i�/��k�\��w�{��ٟ�[x�N~���R)G��6�0��қ��!(&Y�ҥ<Qi]3�I���c�ٷ��Uޏӏ��i w`��%�&��������r�t��Pٹ�$C�*|�������ƿ��Y�*�?!�ؼgԜ��=t7���˅���

�pfs��[�`�_=����\���c��Z����"2[o���E�\�XБ+]囟7��7�	��o��$R�|?m���!��5�QQ�pT�("�VfR�����B��3�EQ[�����Cg�DJ�9���Up��D*K�)o�����tlS���4ځ��d1�hLd�(���h��^}���~_�'�E�f�bi�[mm�
�����������P�LIN�ߋ������i������M!$�v��i~u����(��;�Ҡ7��P�y	��}�"}��9/�gRh	�9m\P�[�����9���>ư��M�W�a��\x��Ȏ)E}�<z ���_�v�������B�L���z6ӟ�93��/g�����	��&��u[ �@����_<��J�Ɔ"߁E�n�G�͋���Gx�&�D�IDR��(u��RB^l�-ï��о�m��kv�z�����_�Ma�Ƃ�<z�b�-0N��]N�pd�f��OVî7�OJ��JSR�-�i�ƛO��o<>�R>��r+9��c�J�i��E-ԡ����w���4��L���ίg}�w[�<���<���PT��2o�(Fd��y� ��a�E�����x1?9��|
��G*���"��_��PC��C���a����\K���%� Y!VHy4m&�˲e����cNSAه�P6½+��Y�p*O���b�k��B����{�#�%��O.�T��k~~24��x��\���gxB�d�߃?jVOϯ���3�5���E�.s<%\o�c�˭_����&�}�p�y,��j�R����E�=x��:���0*� �i	nv�Σ7<~��'��J��5^l��hM�����'A4�_IH[db���gĺ�ɣ̈́,u�Ib	�)7�E@�K�|�׬��O�5�0;ls�Ҫ��{��͙&>&����,�Hk"ۈgid���#��������j+�_�� ������o�n��FZ���}�n ��+�����w�ޡ�q��{�͈v�Y�lc���}��i�=~�[��sPL�!nX�F�U�o�Ѩ�z�}�|�#�-�^ݎǘ���4!z��wz&7h��4���~Wp9�_� g;�˃6
yx����
�(������$}�n�p��h�#��Z=D\��0���S��pX ͹G���_[%��L7xC`�Zsz�^TaI�UXg�c�e�B�P%���Z�ӽn!k�AIMR�s>�%��5�G5�!N�X����fk���+ �>bm?,J����b�5!��'��w,�L��i���X���o�V��S���S{츢W��wx$���Z�^^���g�k�X�ؑ8'�"h��rf��0e�C�R��X�+��p�4�T��'rX�%�l�fh�������C�����G0gʔF<�?�+�,��T?ս��/
�	;�J�-�lט���n>�?>A��Fv=7��!���.�hJ$�m���<��
��^2���R�^���5����a��]���X��ko�G*J@$Z<�ru&	H[�.ڃ��īD�_���.�4a��j�h�Qy�#*9sv?/N�i�\r�\RU��_Lqޓ�ͶM:YAk}ʆʈG�����
��%�rQ�IMt*�څ����ͭjs���bnS�>�t��&�΃�\}fg��|�߾Y���`�z����UR�<���B���&���W�.%�7��ꈅe��y�u����i.�d��
:ѝ��M����
oA�N2���;�q��h�s��*���wFq@�j�;���d�L����y�o�	/�s(<�M�Y��|Ȇ��<�{y;�Ni5]Z��z�Xv�!l.9�c�FH�r�t�z�;o6���Z"����r�l��g�~�G����� ��{R�?��_�Ώ���aR�K�U�1�h}7ie���{��N�����6��&���fvg9�1 �7�U�Y�ɲ^�̼h�z=Sf<��=�ػQ�Ȓ��B!B������V�{�*��Hug�=A�	/��3�gRC���Z[�U������K�<52f��:j0~RU����,��z11	5�ӺŦ���ym��٤o*�R�Ϗ!�LI�b�<v��&\F	�Ҽ�����G��?�V{3�$DϺ7���1[�����rB�dJ�t�#����np��wδy��K}�ߵ%ZB%a�_�!� Q��������PY�J�z�O�P���?�h����0���*?��|[r!u�vi�c>�:�<fo��;.�, V�z¿�f�dOKއ����Y��
r�H�>>-�	`��AǪ��m��:8z[BHL06$�Nf~���r��e
�B,N?RG"U����}j0�ו�/�Z�p��T���;�=��R���-a,=��=�bgMU2���]0T\��+��i�s0�o��6��^��%#n~A��2�i�Ӏ����p���]}t��1��QA��hZс���]GK)y�^2bUO�|�,���G�����Sj׿ӽ��yr�U���I���]���O�&��iź~s����2��&l���`@1?{NR����6�j&ɟ����*�?͜מ��P00�(ZQ�E�A�����I��)�h���u'\����0a�2@Fա��A~��z�c��.�B�a#�'�*L�� ��x���X��(�Nz���ޙ����c^�1;���s�@A�/�1,)������t�c����S/�E����%'�G���<��|�O�����ח���CnE�&��%��B�-�%fzw�2�/:ʸڷTI�X��~�#�ʸ�9/����[���_\����p��`��eƉN��ICB�~H ���P�+�^���6��O��D��
ݧ�6����s>d��[�9?�AC��Lw�F����:p0���,�/	f+&p���+�3��S��qfb�$�|�ll	�^���j�gɬ���0#̓}��a�ZRF��E�7�� {or�~�@�V�W���1����=	�����c�+�1���8_��إt�Y2�g�ZR �f`�C���� D�	�����+��u脢�����]�?�ՙ��l{��@*禈�%�'��ڒ�ב�˫�Y�T˂̭�-IK*N!���VSUa�=zS]�o����A����|Z�i���K(1�JGO<c���B$�C��*�Ii�xw$𶻙q��@����.��#I6��iO.�2����Q�Kbж�T��y�ѱx�0�� Α��V����z�h)/�G�*������ץH�"U�ۧ��h;�������s�~g°���筏&�t���]p��г��R�;�ϐr#��]C�e��U����Lb)�|v���,��F�д{�d ���#3SOH?m��ڠ+L�<�!H~}G�ɾ��(�`����4����s��I��}�������u������:'!�A�� ����o*�鰹��O<�5�7OZ r����_�!x�c�|�ޏ� [�0N�jn�G���fg���{�W,���v�p�L�	��X��]/�T*ڛhl[���Ĥ�M
Ol%�����^��.��zS��q՜\_:����G����4�\WO�GJg�k�i;�JU�.�
�GȃO����U�
d���֗�c��ꯆ�����\�1���=�	�'?��3�a�b�g��.F������0�`@��t�q٩�\�PFG�l�(N�l��`�b�1Gj�[fxO;�"��R�N�6����9�WQU�85��>���^tc��Y��{�'{�l˻K�{���A���v������%��ts��T�PV]_�S,��Aĩ@��=��տQgC�/{�c��w*Q��<~
A�R,�kk��a�`�È��'g��\*8/i�H�$�_H��f�Ŵ�bj�p��bYغYT���t�`֮|���y��캓����n�/��Dfr&-��	=H5�^o���F �e>���yK6`�=���~(�ړw�䖸a� ��x+��3�U��V�-��G��?�t@��+k�:�:�hj����0\��&�n���6���o
EaD�?q�-��4��l��fgw���07_S����ͧWx�Qu{,���r�vk��=m���??��!la��ņ{��J������a�k� �Ⱥp2eK�
�ү�`�9T�F\ -�o���X6)�k�N�U:'���*���s��Y(к��N��H��S���`ߚc�>��È�~�y�������#�&fB�f�f�݋�>E�W����N�~����:�?��#Z��UIM��@͖�[Ҡ���	����v�.�@��MU��2�$�Y[�uS��%.�Q�.��Y~O�2���|,Z���duz�F?�6���)v?�Qk�4Y�3 `nӆ�,���݈N��5��w���oW~�'5��ū Kqə|DR��Đ[�P�r�L�I�ϊ�|�u�ex�*����&��lcFX��^�8gj'�&{{f��-�vQ[��c��HU���J�7����"F�-��Y�e��K�ZQ�@�qnԹE
��U��+R���q�� h�3yK����Nꖗֳ#u��P�7���u��{~����3�A���2�4��m{���jYk����)���L��ȶ^5�r���9@�Ue>��6T�y�ٮ��vU���nZ��@8yE�Dj�;�@�N8������$`D;�[�WU�#|g��=��9���25����d +����`�����f9ly� �=�&�Z'�ʣ:�%޲��F��Q2�=�C�e�gga��V-��q�	�w��sèփF�rֵ�A����u6�qб��q�A�^�OPi����n�ed�8�e�z4�_�,j�h�ԖZ��Қ��e���*��y��is�.h���td1{���$�8eq�۹2���fkZu#�Fa�F�����]2�;�&4
&M7���ŴK��g�71����������Di����P��Ueƃ2�ȩ+ĕ�]`��\?�.���,)�1 ʲHZt�"��h����fO���������q!	���l��iن-�@1}�n�^ 0�$�Ra��紧O�#�OH@���q9��P�+����=�Ub́�e������V&��.W���p4��̲G��ư��v���8M�4���X��
���m�aةO<ueZD��	; ����x\R}85��� �(�I���Q-�*�ç6u��j�������������@@P�ÕX����h����X]��ݔ�#O%���p)��~��:�}�ʢ�at�-fݟ�aU����Tj��m���b�Ze���pʆ���=�e�X�KPI	�{���2��Ǩ�Bw@���v�HI�v���A�^��G��0�@w�	�� б�k�3f��K�m���b~	-:`._,����d�H5 gƺ����?�0�ܝ?���ʚ$Sk���m�E )띉z��I�>�����5�C5�ڜ�lE���Wi����|�y96^��j��=����A>�T��2/����Ϙ&6-�&~� �7v�^�:xe���r��1�M+cv�8 �i�G�vv(j$s1��?�z�h(u0�m.��<�;\�������UDW"�{���R���|�/���F��@�
RS�*�f7OPk�WJ����D�y��0e0�)hĮ�uZ�n��5v�w(ѻ�0X�3S��.]���~m�'��iĊ��E#@t��W>C9�n�1r�bB�%xtR���K���J�d�sE���Nh�XX�l:^���K��p�(b�^�n�OӤ�7��iD��!��ysqDr�[�ޅ� i����?*���,pU�*h�i/�Ps«��R~��	�=�������"2s���P��[ػ��:�$�A,��v?�$@�.�< �����$��[�j-�/�{�d�O�o�<���`t`�خ~p_9\}mbv�~�\~�|��=li�hrn�%FC7^�@vW�a�7S�:�/:��,o}����Ƶ@�����Z�Iw�P��,�X��F���͌���Aw�]�t�7g��ظ����lt��Fr;���)P=�0�}���%|S����Ç����L��I5��v�pf@�ylP��$zy%d��5��=��"�قL��Ӭe�\_3]��ӱ�I����9H/�\k��'�Y|���x���&P{�SQ�GQ�@�Կ����hg\�"�׀h���D�hx�-�kN�]�-��m�������5�<""3toᵾ�)�)����>��L;����%y�|8���26�續'�e���.�'��S��d��� wfj`�u��AFNl0�r�����'�;r�_���5�G��@fxw�
mf/x�T*Œm�<�t��_Y���SѢo��#�it���	n4�z8��ut�&򇠷`�Ӿ�Yvc��3�8Fo�Zt�?��}R��Ф7���{��cr9<���^ }��H�`sZ�G;����]X�c��q��tW�ʡ��y� ��Yf����%�ɧ% 8��쭹	|B�J�غ�Vu�2E-�p�͝|0cׂ�6
�=�t�����_�h�� k�E�F� /�Pt�by���̧C��]WsA�Q.B��}�_:�\e}C!�̿���f-�|HH=�9j�D�2��U!�d����0���^�B�3�K+��U��#i�m�t��,�P��Q%�cSʕ9�����D��E��y��3�u�<��'���P��$�7��&��s�j��KV#�;�ls���6�D���i�-��ؕ#����Z��T u��B���W3G�����(�'�[��~3�����W�R<����i�w���� ;��u�2���x�0�?�O�v5��欇�ݶ+���d����<5A�5�
Q���7U�on��Mk%{�/i���q@m�^/�,B.Fs��䍔�.�N���M��H�J(��Xw*AdKlMiH��S���d˵Z�=t��C��|Wx����q4�٩���>
�� &���v%�)^���n�x(�N�g#����"�^���)7�򆕮X�V�g���5�n�V����@����U�V+�����W�F�S�F�hgL�&��PD��V�?��y�j��_���!�ɡ� �:�V�J�]���l�bן��W�H1'c�l��~#[�W��������b9�$���kL���g��R���j$�=��B�C�k�TJf>=CIp5Ry�����'�{��� =�4�	�&�;��T���$*: u�b���,����H����<�|>��2$��>��]��Od��?�:*Ø�~�i�e�%L�h$3Ue�Z:
<�P��3��J�{�/�.��#�Q���+`�Qe��a�z��s<�u�G�2�`�� ��yOz�S#B�[
]K��%e�@7��8���0�����@�Y*�:9�Qn���:���%2�BbO�E־>�Z��!�a�'��Y�$Җ�o��NsD�I��8�����c�����L�����g=������ �x��/Q����m�|�O�#W�f�Y��BИ�h�j-3�):[�s8i���U�Ez=s�

�I#�S�:��	���"S:l�Ml�Cie�8�H[{r�M/�p@WCA��@�iV���u�f-f�? 1�7�@�������bTE^�S	/��c�c]ȳ��B=������^X�����K���vQ"��V�Q6�k��уNX��;�9��],T.JG��q�g)/ϐ��a5�U
�J��
���!D��ٞC�4�����.**?Cf���t���T[��WSX[1�!�,[��P�Z� y<=� ����3��="��-�/�[*�v|�0#L�&0�[���r�al����Zo�zT�����zr35�'����̗�����:/�Y��,�&`��X@����'LG[ã�đ6 =p����9��N�R�jX�3DuB�)4��ڴ�a�F��z�H"��z�M�Ӯ��]���׌n
��}6��p�����|���hcRң���e�w�B��������@����1X�N7���Mqi��B�1���h��儿,�i깧dW�Ҕ�/�m��lD�=n\�P��n��EuO�EV�p�џ�Z�o��P-x�6Y|嶦����a~���]��z�o�;8��Eׄ5�eU��$��5Si`�ψ}6�����'*MF���g�NV����Gl�n���XE�tѳ��R� ��q��B=�qo u/0��H(d��~�E�/f��W�G�f��^�/� ��z�"��:�#�z�g����!o��t�
��z[4��J�<7%D$ 1K%_B���=�ǃ	 8,�}6>��H[P���\�'h`�m4��ϡ?�K�x�~�j ��T#�+T�-�M�b�F�Ӹ�k�t�#�6U `W<�K��ϋ*7B}{����XZ����!!��E*C-�0��3�v��0��1;MϦ�Eى 
u2�E��{�^^[<�cO��'sjl�����ԥ=@�<�e��|9 X�&9�F���ũ����q<K��HB�1�0�z;yevJ0#�O4B�Ջ^/i��zoV�+��]��V�-+����@ϓk���?-����|�ͥ��+��9&׈=ܢ�^����S"�����^�ؾ'���`!|d�,�����6Mp���rp%���b�;�� ��R�
��c��nz�sy�E�1���������BzK�&��iђ��8sƝC�ܘ�O\�6_����o���"�f�v�~�	� ���8a~��A�Tw��Fsv����n��4ۀ"�����&pY�Ny]Q�O�Oў�C*�?�EX�2����j;���zX}Դ��}������i`�~D�p��l�����]�ј��Q�!>Q>z�bB�t�b��p٪� �����$�$O�� !Uy��p[R�k��&��~���-��p}Z���"���cV,���V��?���{q��B@va�����_G"v��h��1���K�T�g~� �����Ա�ە��0h�9Y���%�#� �#X�E�yr��� ���y?�\R�ާ�^��Vc<����:º`�DG�(H��Jbϊ���߷����f-ʍG�<��-*P�w�Ҩ���mDZL3�_���" :���X���N2�b�e��>��������k��q�=����#Ej�u
�N�l�2�v�9g,�xk�9Qҏ96!tX*;w�9��޾13�~�����n�N|p���Lqmw�6~���������Orԛ���n��mF�з�B w-�*�k(��e�.�z����w���El�(��̆N�N�۪)���ڬ皣0�JaC7B��Hy����⩎���8~G��qÌ����\|��J����},�����Nhvd��=e\�`�(��|#�$Gh0jx�S�2�(XG�5��#�����L
Q=܏���/QB�`�c��!�{d��Y�E��A��!t��+nŖ�kߩ��R=��J� �#r�[qE��0�[��������eʊ�ͨ�Aui3���}h$����-݅�z��������� �g��$�	�cҷ~\�M-\ew0��2kL�wpbLO�춰��|��ۯ8,^�j���mV�$~��&C+	g���f�1\���z��m���;M�JCS�#9~�amM���+�{����"L�x��S�Q^1��r}����E�����c�8�d7A�M��W�e���=ALڠ~7�(�i.��y��E6Ä~$��y��v�Ʃ��];k�o���C_��_+���P�%��=*�Q^qی�&X��h�jMy�ܷ�м]h���D�J%�����O�����ˠA8��C�6�u	;��ilhucJ�&=J�0j��YI���",��6U�+U�^�
���l�̪,l��6���f9������!�'C�i�	��0+e&Ļ��j^�zю���+��U�^��Q[�|@�L�4�7���^F�uK��E̓��8 �L� ɧFP�@,��2��}6�����M�XLܮ������V�/��J���
���?��B$��d�d��R��jve�}����X�ݐ����W�$f��`��)�iTG 3*_E�,��	MŸ��
.QE[a�J�:b8c,�7��]z)4i��z�]�\����5꒧f?����!
08{o�(�_׍U��i}f�b��_>�W��|3HvN�d��{��-��ad.�{+�v-�cB�*o4�,P�==��������9/�IY��O�Q���ռ��j����*�k�VoP	=��qX�B,�䊧�qe�����9�Ʈz�,�w��(V�a�Õw�)~�;5?��h���H�k��j�@�&{��Ҁx�⌃���A�[�r8���r_Jט/���z�d��&|�o��t6W�Fެi�<FN���F���0�]��������k��%^�f��>��و���sn�ť:4p�x/�.��urs�(�uP�V�sf�/z�_:���V�0���i�mkU�����\�nh\�R	xJ�Z���&偽,ߝI�C(�R����2LO�M�ҳ v~$�NG���qB<�E��)�ߏs��t�1�I����B����f��f�=9x
g؀��A?O�M���&�ʿؠ�
�uͱaQ�"��0p��z8T� **��c��J�sp6���R�tA�4Z@؈�kgǵ�o�k"���
l�Z�6�Z�?�(�+�q�>6�:"�V���
��*a��?�'[�3zF(�$V����}���`'�a������0N��@�F�i����p��
V��'�e �H�w�A	�:�����|k_�wn�L�yژǞ��/�J��톀no�&�`u��$�z��|�Ã*�޲r��5T�E ��!S��s���!�V�ks�C_k}t�G+]`H�q���PB��V�̏�f���=��d��ne���AFo� �9�(����WRIj�!L����1�J��3�~�Z�[���!b�jMZ��')O��U^i4���6�u}#���ث+#�����]���N|�ꍡ5��$��֯"�8r�i�N՚�ق>S�Ӱ�z��]�#L����7�/4)�v��Tr���M��4C��Y���AB�����N�G�h&	(�_�|E�gWx[ʡo�- �L��Z�h�`,��Ȋ(��ɥ;�}[�,�"�D��7�YK�<�`(��ӲS|�7�쒑�47^��j$��p'vQ,�[��a�q�+��W�����e^�Ғ��
���;��!i�IJ��Vs%�
M�G4�`��1f�+Րw�[�1��GѹZ��B1��6%L�;̽p#V;7qK�oļn�#��Ƿ��Ԟ�) ��V�)�,�HĽ���>q�s3��R������[I�s=�y�R�s ����@�������T�8�ձp$�@X{Dzv�Z��{�q�S[�d��0*r��5s���������E53d�B��˲�w��&�]*����-�uǠ��s  ��'��M��!Z-���A^���S���������)���h�U�2+�p�R%�\6������|�G�(yZ7����&o6H��A&��ڍ?Y�weR�z�l+�4�?@�����-��LP�	E|�`��0���P9/�$օ����.�c]�R���!L����s���0����(>�9,
�3i'�j�����׈מ�H7WX8Kx-ɬ84|[�S�S�q��k x�Ͳ}��s��}�1�
zt�*˿��$X0zG8G���9��[f;���$��K���(���q��:��ń�o9Y�jE�Q&Y�1�nK sg�4�T�x��"�,ʎ"$3���Q 5�$����Ct �����C
�g/Q�yQ�xn��_�L�ݤ�Ճ��,���t=Q��z.|-pW�D�s��ÿ=�A�]�~��t�dM����TV���/������Xd�$E��ֆ�z#�t$�>|�#�ӳ�=�>�fz��t���ٞ/i�(��R��}I�0�I-x��3�[�%�ëUA爃�Z`� C�Mx���4H�<J��),��@��k6{��[�I�;__r�uߊs4Ps!�0��_9G%���O�1˽� �g:�^�/ڎ�g�v��X��P���8��l�����{\��Lp�����?Qc2&{d܆��Gh$98���&��,η�f���q�(�S�V���R8a<��B\{B8�UFu�?ڪl A�L/F�%s�G�>������Ke�~�k`�b�]��1��s�Ho�a���8=��p K��lׯ���f<:�W�A���J!����[ۦ�F��vS���R�ž���ȕ)	�3�E7��ߵ��v�ji5A�@w�����lW�V��Т4s��q��+�ry��5�H�o���5G�Զz�*�0!GIf��X���A�v�(�����6�ne(	�u�..Jb�L�H=� ��ک:Xz���g����>�׫�~
q�-[�n���է}w1��闠��p����}ID3;�+8�Z#��uw��3u�� �n���-��.�b�N��-<V���'_���9��nP�Q��%(Hv����쯖�>4+�@;���� gH9K�b�g{�n2&���0�����Eo��)�[>t�#�+�f�* ���D��O6V[�g0S��pby1$�i�1ˊ��Ŵ�M(�FK����	��_�>x1ղ���0��)7q_3��L^���O~^�'��vG�]�x�rz�סȌ~^
�mS���^�X�^�<A ܑ@Axo5y�6V�ϛ�8n��s�0�˒��ھ���6��]=f�g�͖���Z�xd����	6��~UFk���µ�v�#
+X������fȢ=1�cz���Ŭ�IP��Ƞ�unv�_m�����3�z�3Y����Ē�V��XN��<�B�SR;�¤e�������"gQ�H�s�Bn���/�vXm �=���c?dI�Ҵkle�}�&�G��b^�� ��lJ0�f���u�k�'?�f7>�p���\H���Y�Nӑ����nIP�<'p�?\J`~9���$x��03#�<:P=O����?�y�3��-.�� �D>��V����ط^��O?��Zȃ��N�zm����Df����>g������ +����@kg&��B���զ;[��?�k���D5���7�Z���5k�ߪ�/{����N��vO[�iX�yxkm���W v�THI��I+� b�6�I��N{8��U�c��	�5���d�zc~0"k�F7��cV�,�F ;6���.�&	���x�e����}�r������z�x�h�m���|�p�V��HB
D���]`�F,���W�/{�>���|�bWlJ�e-���%��ɘ�
��]f hN�F�fyU"���??�4rx�+z���\�s�\<��������Y���?ϻ�*1����5L`�]ig1f�+}f��fz>�'����E:��)]� 4o���d:���E�a�h!�WL���n��B@"r�������2��٬ҖD~2A/T�W�N��x�PS0A��h�M	��aɿ�ʹ��v��'�� !�)];.��9�u�n�9��p�^���#w�ڧ������qJބcn|�7@��_��{�:Ƅh�z1Uܞ;����[� +I�^T�jp��� 3� -�'ٶ �����A�\V�]`�����F��Z_��@8bJ��*Z���l��Ә޵�
�p��6�����o�y���u��5~��i �B������ �n�N�O R�It�Ł�m�f�l}zO��k������*L�7Dt�`��Ë����v�F���ӝh<:9}�Ϡ��Ԭh������^:K�Ո�Аr8�w�,����ܚjb�����;.ҪA��Dad�7զ�x^���B��(pƽ��g=�x�Y@�\&��ږ�yj��O��Կ"uƌw6H���&��h��NNsz���됞�Z�|`}:�(C�դ��CKcY�iϪ��c���y���<{�{���u������fs��|u�#�0PGT���G>b���r�s2Vc}-(�5�E��0����޿��e��r��Fc!����r��f<A=O�ආ�� ���b�\��2z(�:���$�� kd�sَՔ���Ȥ����F݇��WtH���>�D��O���?���N���5�z�i������a�8�hCBG:6թnFk����9'b �rM^n��r�	"c�a���W��#�2�5fG�4H�ً����mNB19!T��5bm�}��O����Ր�����\���3/��O2������*�������
�u�o��_ ���t��A��XB��F���K"5
�����Bd����X��Uw�,����~d�9�K�yw�]r�車�C"?�/�@�\o�8~b-��Buϒ�y������'�O^/����~E�|~�L�h${_�So"��P���~a�+��>�JRy�m����X�`=�ߦCK�>XP1�n��<�����I��FB^Ӛ������b�s
��[*�uHz��k���K*��ek�tO'-��L:�� ���%����H'���ܐ�+�Е8o!a�t&G�J�wY��:�yxT4#�:����J��K�/,����$��P2D��������fЫ.��˺'9���b'y[q��g��IӲk%|&���B�G�����ڿY�@�\{m���2'��e�aaX��#�7۵'ŝ����Ek�Λ���fy�N�H�m�KL����||����S�]ã�Y0)/�c?��&O������S�`Q��e�V�N�y֯1�����2}Ӡ��0CgݕɎ�F��U����>��2���SF�2�u�CqB����R�+nk��AM*����h�s�?�"���
�����$��g�P�����t�ϟ�ζRNcN�Eq /�{� P�M�4�l]}R\ShP6"��}���p�W��Y�[Y���i���pKN0�����}�y�f����:!�2��D��:�C�NWm'�xxʪs�3�hm�N&'�QYd�l� ����I�����-��ذ7}Z�T�RGD�K�g�wB��5FS���%GC��+�l4/�f�P�b?~�]+���'���ct��˱@�|�$�%��$�{'J�؍����[+��i��x�x�T88�$A��%ic�2��35��ɡ%�'���YC3�5�x�!�;;��{!d.�r��hղp�ޞ����"�B׌��&B��!�)�Z�+&v��o��&�����k"���Oc=$(v�Q�^��ѥ'5.[k�[l�r��s�T�3�C��.�wK�ƹ1* �|���� �>$yh/��Sn9D�����)�:�l@H�F}��O,A�X{���=В�f�4��l$�6#?!Z���2��_���1,��Ӭ(�M���:�7yJg�7�q�R7ō�m�ew޽���Kn<^�^�c6��;��fۓ�\#w��3��*�^���	9z��	�n�Sõq�P�g4�(pӝ-ߵA�8���3�r\�X��I��$�0��uo�lY��؁*/_<�Y�=�~�w&������ g܇�)⟴�u�r�F��	��/ m~�;5`c���5
o��c��_3] >�U��J�(qҌ;�턞V~cd�\x ��!�����
P5jISd�f��ȹQ�Y�Չ�ǺOz��I�
t*���Ì�\@�+ğ}�� zzW�h�|f���t ��͊zrsw_+1����r�����ә#V���c��VM�n�z��^��l��q�&6FB�O@F��]��ÿA����+<�ߟ��A�@����Z��[�g�0�,�J
�'[���^�5��/��oA��AMB������u;}�c6�(e�B��U���q�HK�^��č�R,� k$��&4/#�˘+F	�L��ׇ��~��ݽ}���Tl�/j\� �Xs:�)\��r�p�}�����W�Q�r[c����̶|���� ��vM��RíˎEk�(8��5T���Z@���c[��`v�|K?n�X5�+<�3��ͷ;���
!5��9gڤ
L�>�M��v�� ���U�?d�=1�8�����]�p��4�1��Gcb�'41/I�E�:��1E�c��@����Խ���6�L��9uH@_����s^0*��X�� ��*��w�e���{��P�X<~�1\oϮwe���Fw2e*���N�e1ax3r��J�l���p����yиsR�T�FQ[�[oUiZ�{a�;Z�3Vw�o�� ��߯*P&MHj���/����������L#��2ᶺu.�ŀy���2-,�;}6�w�����u��g��w�%1�T&9�]�[S� �i�1����s�Ix���}Js�S�#�G�#�0��4̃T��+���C�J�!�T��"��[�v��ki���R^<v��V�P
J3��uu('���LU�z�������x6�BD�7-���H��t�w���Y&�r�� 9QN�F��S�6f1�¥h_N3��Nq����(��tB�Hb��v��v_�*3�o�"���z&�B���a��V�U�&�����D�����CjGL��$}��}w6�D�TN�:�{]u��"
��ǽ���+�_F�T��2�F�K�sh0���l�j۸q��;�2�F!�Y1��<1��Dq��'���} ��l��o��da�fpT�F�ug:D����x���K�LRM�b�ç˶f;��+��tz�A�Q��������P�A�wVY�S|z�t+ئ}�,l7����[�@��;5H�б��I^)U���F���k��I�Vw���KR6�D�������˳�="+36��#�����iB��R�:o�� ��pU���Y���z�U'���������/Ru�������yHY��I��b�o�1[w
�ĳk�4�Ʒ��>@�Rݤ�Ig���"Ge�N�h4����E,���k6�{^���,02�E��Ai���ݱ�2z�v�0pK.Z�;� 7�����>Z@�I���s���K�~Z�r��d�5g�e���)vD���g:Z���DSW�;T:?�#W�MJSW��i����k�Q��J�w��^��!
@�+^��l�D4^ֲ�%�%�V
ڮn2�d�p����!&p�V���8�|b�{p,5W���I:��FUl��7K���h3�^q>ňKl�L�� �4�X�h���\�7nq���$� ��3�zßI�{��>Jl�B����*9���������QhV��ȵ90�>���p�׻���S��P��&S�e����O*��[�7������z��?���jE �l�|C����j�$�7�$�V���`=��A8��:�_��b�Z%���s�৲\.�>��$�s���T�ܮ�[@�Gx��?{� �>����j�V��8��&U��Ǔ��s�L���#�gi�f]3�o}�M��r'?\>g�����-�D�K�
�E�4�\=�aA&'�҆�3�3hq�R�^Yv�bA�,xܹ�
D��`�Mf��.����5���Xj,;`��26�Ю��H�j|�H\�˛;���.z�s�?|��u�	�|0I05��� ��x�.����ƾ��ՠ]�x��Ғ�q��}96�C=O���h��t��Ӌ��tlSJ��1�i��	�2P�EC�z�k���A
B��ƝЦ!�9��V\��(1��-�L.q1�G��3#���&�f��釖{�o��+�N�Ѩ�� ��(�o�a���t�fAkRU��W9A�!7�vb'�8��;3�5��5���m�Q�""�D8�����d���Wzĵ';�A�=z*_r{���\����q�`�nOG�� �cm�g��5S�>.�]�� ���3;���hEN�Y�Y���@DdY�r7���^@lj���ԇ�S7�C=���d�R�A�� Ũ�4yV �,��g���@e�&�k�Tz�|���ݦ漰cB�&�=w������x��*��_{y)���}�%*R���8�2�-e͠���l:�8�,):�N��@GIZf% �/o]� ��gY��l��f�kp&��<@�ř]^	l7-�c~������DW]Uek��"X�H@��v�xp��G)aX�8 �;���$X�S�1 ��(� ����易&;䌊Z��-3+����2d�\p�XP��l��ݝ7J����[�����sc�b�~�I��X���Nn�y)�cI��0��D��I�#�J�[��7��9�}ϐ<Yk�Lro�-�"�������G��.&4k�6����u�3{���|ǸwA~��C��*��;����7��")����E:���̅�t��Q/i"��Ϳ<�ԗ���^�k2����*���T�{����
vM��{�I�Y�|�q6��65q���,u�1�|y�k-7J���
����s��B�bc���/��w��G�]>z ��R��}w��1܌,^�41M���g�K�:���̕@<	�i����\n�E��@i՛���)�x��y���AK2@��Ir�����"�Z��
+�l����:� ��l�q"�	�����?����Xe�ob<	:�sf.��%y�����dyr�
�5F��ڀq����T���J�=��F�N��cY�����L�ȢL]<cv�,d_�b����/s,O--h �E�t�u�����[�a4"D�KlS[P��߹�o�������$�ۃ���"���]L&��K�E,�U��%4�q3��3�&(�w�w���MH����!��|��!,���j�q�w�j��ď�N\5�b]:ܵ��匒G�{.]��ff��DMUz6熜cpE	�%0nJ�Bw�\e\H.��>����8� ��?��3�h?:N���Q�������������?����&H��b0V 1M���-����IM�M���j����z��`8�9@�P�*4��L�yA����=�R;%��+���4eB3�p�tG"D�r�^f�J$4�	��T�Ҹ�$��E�/Q��׎e�?�M�ʘd/��C������[_�	�G	�]C�.Ь|��
�>�-����R]k���~q(R3��ت��#�K�����u7T�E�se�X,1⎗НO[�^��_�\�@���(�ӿ�[�.�ۻ%�}�����E��6:Yv5�M ����EJ9��Ѫ��x��n����n~w�׻RR5��z�&�W�ek0�5)�+n��z��v|q����3���Z�>���1��umQ���g�w�C�M�s�E|��r��Vy]W�I6�-�2�pL��N����#i�8��e-}�	ǫ6H���q���:2y�����!O2)�8O�܇� ��,Љ�{`us��N��J���"�%/����e�9�tť�!
��StUbN;�å̐0J�]1}N�F����c�)�����w=���TD��-��J1x��{�N�0bBE@&��=�!���l>�{8�r����c�@����l(�`}�U�>.��=*vE�+yZ�C���W�����ÎڿȬ�X�x����wr��M��h������L�n��[��W����G7?7dA_~�J��/�0-<��;=�-���c� ;��p8C�m�k�F?�fZ],���R�C�	�ysݯ�l�N˘=���M�Ls}�
�7M7����%]�G3���=��q�.j�1 r�y���Y�8IH�"V�o��^Q�V>]�HH����:)���ö�) ���^}E��/1�<�����Ɔ���ޘu�y��$Im�PJ���Ȅ���ԩ���R�"ޮ�
Q��'kn�7Ck���zԫq�V���远�?WP����ڈ/�6�Nu�<��Ͱ^�GTN��>zέ�����O$2�ĳy���Z�$ǐ�T�������>]��	G�6�1RC3	�bP�?Ѧ3�d��6�4��1���psY�VBV�u�����w���t�AH�̳-�!{��a���
���=o��))��o{��Ɲ�|P���	��02<^ś&$��p�����U�O}����������<��������y���G��'�tS6E��� ��>`��ہ!��@��㢁�ɿ��X�j�7�>�X�2��;�|��#��@n�жm��ޯ#o	=3"�;�iU�#�ktS������B���-�s�c�X�w G�I''Ʀ ��6Rf&6.g
c��nV�O���:��ŗ����Y/���T?)�9����]g�⤬�d�Bn��_�H�2,�Vr�:�\P�i�ۂ4�AT�^�}hU9���˰���lk����̏C��ޯ�;	tg��*��T���:�l�J��8Y16�k0�Ӏ�+E�;%>[YUT����	}��^��:������l��%K!�w��m�P���b��QL�μ��S�����-�yEk�����p�<�6�54ۚ�V?mL݃���uv8��>t�z�R�=�h�!�LQl�QN|6Cәabi_S$t?���Hr�;�v�c�s6a�]hB���݇���EB��T����m'��uc��a�]��^Nnr�6��W���[�0��}	��ΧY�����/>�6��WB�L_��
� ަ��:��R����n�s��U��wچ���[�S��DB"e�8\5�b3�XʍvIL�����k	£"��d�)��5�$2�e����'���8��6�7@�����!]�nQ��N���칦�KY����sA��d�n�d�h㽙v����Sn4"�k�Vid2���nN/@�}���'��K���;az`�[�[;�Cu~s�t�눒�a��¦'LՋ��?��өt��O��[{���c�Uc�o�{�o�"�-�M�X]��3E����Mf��Nuj�Q�g����{c��
�2�#���<����Z�[�>�@ E����&��
9}�����������|D=+՚�Y�9q�ʚ�қDI{�(�������%řmb@n{t^85|?Wd�/N�Ks�-ʵK���w.�a�U����>��m5Gx�P�����"��t�Yd,K��uͧ����jFON��C��V�|Koɂ��%д.۔e�2����a�ȫ� �$0��y���/��&�����X�`�l���˘ˇ�p2�o}5X��Pцc$�(���u�d�'���+�AB��6s�6�V%�V�w'C���n	,g�����E�l��S�A�Ϻ�k���!$�.A}\N�(4��NYԡ�<<w�Q� 
�&V�_�*�oծ�f�%�ˇ��
���;Bt!�P��e��N�!�W�|wc�'�&�P�h��5a ���U��
 W�D�ޅ�w/U�؆��5I�c�F-����tta5�1ϊd ��pu�l��R~{�ǧ&��2s�.�����Q/�ŦI$�'�t
�w{}C�ۆ7��dH��;>�]6�](|�����O�р%vL�)���30��$6 L�l
��S��^��֬{����6��e���4�=�B9n�G+]A����ɭ��r��Q#�VY�y�(��T3��lB�7>�����+�|­�+��Gq
���e?[��)�_�@������KwY�����#�e�33��L����������7��P2S�y;��Zܼ�B7�A�-[-V/�{È�$�d��3T�X�U�w��-��	��Q��^��"�����5�3)���Zk���3)��i��D��v H��W���$*�ih�����b{�2&��ˠ��hR�0@jLX������1���5`�S]=�3Xʈ��hLS0%Ϯ�4A��
�F�N��E�;�8�fa���+��#�;nm�0u��y�G�N�@A���xS
8�`LL�@Z}�>i�ZW��b��;}፷7�b"5�Df�A/��Ét9+�=��f���g��D+7�t\H����R���7���A���Qf��\��T �fF����ٯ�VO��q�M�_����V���h��U����ɍ��~R��F�J�Kɩم{��g�
��J��o�Mc�3��Ħ�P��Զ�8�8O>�z���
���-��]�.)}���y?�+���I����{@�h4C����4�")��(K�
Fx���3�?f���9RV�O7��d�|@0��0�	�~������ (�Yw��2�V���C!ڼW�v��ޖ��Ġ���pP+{�D�Q��Ũ=�]�yIR�D����?Y܅��s4|l@�HB�ڌ&�Tt�Ew^���0}Mw��a8����A���x�'��_yZ|��ɯ��%ڼ� DPg��k��<!���倫؀�<��ڪ(�L8�Zk7��_[gʓc�=
dSĄ}�8j�����̩�F�|k��b�!2���3�����]��w(\����{Iu�݅��Ѥ�4������d�;�t� ���2|� E��rG p��h&
-�PW����X�M��0#��sJ��?	���-�?�7����1$wP�Mv�g�E:���ቐ��%��S�+�N�G�չ�ڞ���0�9u)t|}�W��]ox^���4��0&T�6��+���[┥���.��C�;������]�ӛ���(ۑ�Bt��5�7�u{�g
���J��G��'����Q��!��0�㘀����qP�P����f��x�aOgb�Hn���i}�����" Q�v0:OǙ/�� n%�g�?U�n�Q���T�;5��&�'5��N5P�8�����9���헍�
@�|D��.*=�xAr"�j�&���(��ဦ��6�hd:<`7�i���j3��Cf�u=tM���G���,h��$x^RZ�\LI�s�3�5M�M���נg�nh�w�d�Da��Л��(Ĩ���%w�"-��~܍�V<}���K�1�]��ϸz�SSF�_ɱ���-��ö�KcǛ,���w�p8G*�ר3G�3&B��39��� g�Θ)�=|#��l!�֤�(*�]m\)I��%.x�ѵA>nB �*C�;�o2D=@}m/m�����1,lmQj�߂�#�P����:P@�g�ύ~�͇����S��Ғ{��T	E�*�J[Z͹�4��;�����6V��)���b0�y�f���_���GR������ɀ*�u��
�6M���O��w�XqM�mm�͢�p��>�?���_�D��-��4�	��_v��h.EO�=m�����?`�~SI;�l��<k%���b�����?��^X�F׶�k8�|T�v�tjߚ,Qw$Dej�\��`a�����~�"�4��Es�5�؜����c#�F骪�}g�ڶ� ,0�bLX���֌�E����T2η��=Ϫ��WϻR�z!�R�x����F����>'ľ�)g��6쉞˴f:�U|����f:��tj@�GyU�#��D���ڨ��K"T[s7t���Pw	�ۓ��^ �����1�`�o5]g����Z�	�!�j�quҜ�+�s��ʲ��b~9��Ł��6kº2���B�@��S�Y�O��)�Z7!4킌r�9�~߸���(P��BԼ\=p?Ecؓ��[�VqS�@ǌ����I��ğ�t[u��m�gX7���$RNo���Y����	l=d�G�� -@�%��-�
q؝A�T���[��5t���3G1�����6x3�b5q����֒�ݳcIl5ڦ���s�F��q<��(��/sb7ؽEY;�>�z:8I���_ݟf���!�q��|�[?;��2�?��Ae���',�R3�:<�o3��lN6P����${g�>/�[Q<�)��|�)�v��]K�2�s���\�a%�q���*�}U���pO��"�#��_#�+|�u@q�X�HM�w�?.��<��;2Sr��g�xP�C�VF�7��w ���^J���2h�k�Z	��hOI�CW�)�O��~�m!�n��8C	�X�Zd�>�f7\y�� �\�x���+"^�?Oa�si�J3	�F��	��E�����ua�ѸX���*���]��ۑ�KŜ�Q^$Y��`�C��'�[d�
3`�$��ݰ�	��I�@#&�T��RH"�2���6/ȭV�~����<��P�s�&,��o	�vݑ2�˩�ߘ������3��)���~A�ӄ��	��1sνcs�l	yƿ��$U��/�8�������[�߭��2.7���R4�1��Q����9�.ݳU��6ٗf���f�