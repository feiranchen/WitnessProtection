��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l��$p�c��U�W^�A�K�I!��(��`�˻�m�q�枒�~���W��uc��^�N�����Ʋ!5;��g�*{�܀]^�m�gB��Y��M��3��P�Ve���tg�)!���{m���j����K�[΃��r4� \ *ХF�:}YǛy�@���d���=
w=�r���.sls{�z6UMѫ�X�Ӂ��[��|�ԥ�I^�5���.z5*�hA#.�T�pm��b<�n<:�� o~�k^o9��x��Vۤ�_����3�,I�	јSkV٪���Q T��+6$
v��{�w�(B��@�����#�b�����Ӷ���|[d���*	$Ҩ.yPU�v&6!�WT~�h��<��g��	�QM޿]�_�2���aЧ��2�t�v�5�_S�[��ؗw���1#�gY��ji�u��M8�y��@Z�L��6K�e�	�����6[��d��w*̯zu�Z�xʬi����n��rE���D1���i�5x9�)4�Gݼ6��|�1lƿs����]�G���r�a���F�}��n}�4�v��g)����U���h�4�J\�EXe�j�I�r��xk5��2!	Q@��j���O��J��ZT��Zhѕn��MOŗS�����8U��@�A�O�|T]&�V�r�~�:QK:ļQ�\�ar�@��
/�>�p U<<�V?�1�+��#�����|����<�@4���P�E��a6�;@����'���o�O;ّ N(A�v���6_�7�X뙉z]�Ǜ�@}�-4�X���<<FPz�}s�`#gk��w�\A\|B��c��7����b/ru|4��eg�lck[�x���,fŸ�~�o�~���;�<���ݐ�;F-�ƈ���|�uH篛���#ƦԸ ��5Qt���NE��\�a4��kSJ.;V��$"�K���`���|�E(ٹ�V���T�C7[r��l�InІ A8�hϻ�,3�`����I�����B���"�<U_I�%`��H����VVw�?QA��Nщw�=T.��>J�iXv�&�e^�u��Uly>�T�u@Q��Bl���w3MSfEz��cI����gm
�jE|= HfP��;�c�֎�>�Ϲ@�w~�)܊|4i��u��'f&o��3�3LA�27�S���^hN���z��l�r���60��-����b�4|�8�.4C��$W��H�fC��u��	X�f�
a@�m��2}+��5�#�C��׽�j�����&�L]�.�rs�y)~��������wt���BJ��7�p����A�=��
�m�'�lZ��F$Sy����??��r!Ʒ4A`{w�WN1�1���5�:nA����S�o��M�y@;)�a�B[�M;'\�l!����O���A|�UF1-��>$����b�,�2<�C�+�&�O]x�M�,�?��w}��؊��K��&O�_���H-/O�վ>��8�I Y#���:�޾`��ק>}8�e�e�[@�$bV�jW��Y1F`���Ԟ��8�ԅv~��};�~4��w �+M[����_R"�Ԇ8��1Z�_��N3&5���Y�HLP��eѫ���)�Q��j�;f>s�����C|�ï�Il�^�o�'z�nN'֫8�/��R�^�5D�hF� +�(�RE{���p�v�!^�����ل�{�[a��;|'wD	��&�$،kLAS�W�=�9VH�� �� w��T�_Ï�C�_��C�F���L�����M;��RW��?�y��
Ϻ�E�ڜ���,Qqͷ���q貘�
�����lgxt>�5�J����:/?���D�gm] �l	��qIE��"<_{ִ0�u��9f�y���.�2ߍ�TPC���T��I���J��lm�i�準��S�U&�H�5.�r�?!u�~W�Kǭ)�BN:�i�نN+��'@�I�[�ji!?k U����2���^O��/N��|+c�c<�«�d�:v5��ka���b/�@<rm�b#��&@���J�����}�O_�´�ω�8{Z�D��`���������/;1��Pٴ�|���(�F$�z��a.���-vY �� T�U�p���͔$�ےkW>[l�L��%9���O-�6	��#"M��"�ߏ�AdE��'ſD^�?�|���E���*E���a�¢��FT�����`7��9Xn�`�"L;3�Vm+9�d��
����9ܰ��aJh��U"��-�~����M&�tǖRA�!�4;�#AI���_��45h��ܳ�F��T(-���ә��wtH��;���A�OA5������@��q�> ��)q+_�3��� u6j..�ڡ��L��� VDwJ����c��o��/�jbd"�f��bW��?N�K'�ݯ��by��ǂ��XZiu��"ܙ��r�����m�
D�S ��wNvx�g%d�O�)^���sA�ҜQ�EJ���f{ݎP9y]H�ai�u~K{��X��K^�=&�h'D��-pDȁ�9�zC+�1���{b���Ź����L���ŭ��P�0K��w�������@emQ�ʅ��v�P�m���>�ldQ:�ԕu���؝�)6f��`�x&�9��u�cK�Ǯ�g��uxH )�'	�䖭%��!�ι0
�є?��R��<�ܪSݲH :oW��)X�08q�y��B"��V�����_p����	8��$4���x��2��t�
��J������b?�Z����s.�5���W���-oz;�No�oR!��9���4%�����y�bZ���
"6}v�V�G��@q��������[�I���>����6-����	7�B�J�GaS０W����Cjcx �;��ɊX��UM���)���=r�-����#un��t0��I�U*s�g�Lr�0�dI��Q��5���N�m�����sDOf���l�������O�h��O*��k����yo�	.DqL�Z]�̿a����Acj(b�[�3���T݇�,�ߚ8�K'��1'mp�(�}���,/���ɡ��,U+a�N���T��M7u�f�sq���%,iN�����W쑌�������-˟�j:j�;�����4"�)rGN���#*�l� � Pa��f�%mTu�Χ��ԳY6CP�z����+�=�xC�	�=��Q���ͰLlt�W4�]�3_�D�
X#�X��GҰ<^�R�����C�����U��3f�OO����HO�Xk4����ctpZ�w�^��8�a��ϡݨA�E��:Q����D!qj�c���u�m<I�&�$܍˨Iͤ]b^��%��d���n�S���w2�(���?/��)����H|�iZ� LMJ,ٮ���mf�0��]���j�k` �Gb�U�ޙx��?_�U�m��"������
��io�_�3P��@�u|d��G��ؑ&Ƌ }�&�;�:����Xv��V�em��\�>͕_�SC3[�&K�^7��-h-�"������!��#�(_�R���M�PB�|u�`n�Vλݕ����Wl���I/��<;�+�B��
��4S��S��Ɂ2GD@�/��0�24���%�^fc�G��7M�t�0).�M�@%8�	A�	�3j�ѤL$�-�W�n^���	J�]��y�c*�p�d�MC`�Չ��
ː>���r���U[n%�P+)��X�|z�j�?�΁�N�f��5n���i���:P�_+��5�c�<�7����ɍ�����x�QX&z�{��a����hdMk6��F8��䥮�ڭ#�>p6�1�8.�2��5��<!!3�2(Rz���d-K��KnDY�]7f�jh&��0w�T�۹/��-���{q�~�@�n�fМ)��gMa!�Sp���9$�p��Pt��Þ�d�	�yP
Z�"�_KVVݱ�3`�k���R^TTo���
��]��B�R��D�A�o�,䞣�fΌ�ܵ�i@qUWl�1:��R��A���=�-�a\$��@��
VZ������w����9Q��D��J|b(��<	ڈe����Q�c��B�G�t&�B���;�D�c)>�h�U���-e������%j^sɍ���s�>F���#�
�,;qm���A[������2�xa���6ű��}g�/�2��2��ԻD��˦��� }yL��&�[@���I6���p=C�>��QIG���A�X:�O���b� X0_Ъr)Hf�{^�N���^�����A��$��ع�Ɯ��{uu8a?6ܱ�zQN-��� ��5*ܻ_3���RJXgD}�v�ͩ`KwƠM�bPXm9�~z,�G1� �Ŕ����y��f��\�%D��Q�'�3!�;������֚�����Ǩ4�./�Ӈ��>av��7�Vf�\�~��i���E����_���(Ewp���a� �%TBN�5 �v��B�n��q��Q�+w6����^�,�/#)1��X�EB[��(��v�y��~�	��{�bnj����g�S���%��(
$d��aa�P���L�p����4�&�XW�������!*�N�J����,���4~��F�l�&lk�9z8��FL�y�#�P�P���z��uĹ��Հ@ �⻼G���M4��Fye�4�v�;U�,��j�$�R�A��=t��h��Z�7]�9n��D򓌹��)r=���OA>���4��	ov�귨�_��r;�aE���]?��|�0����^�Or��͸M	�u������sg�O���';s7�*Ը��