��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>���q=ԓ �AJ�uU��W�i�#*(B�u�S\�mL�9\[}�͖H����F��H=�a(�U��rL�y�^.\d�x�&(�0V��穰��CZOJ Λ�I�z��$V�GVV��oc�z��06�Z*݋�4�ɪ{�BR�M*�=EL"� )eb{dq�X�AO�
�s�Po\r:%ck��y���2Ed�F{5�щ��4Y�ɷJ� ��+�Vk� K��	�4�netg���*��b�o��by{ٞ_J��k�6TH�Q�#ur ���j^	����b##���RN��:���=lt����e/����kcO�e�W�y�R�k#�����뇕
������x��<u�G'%�]�]�.ᮂ����<	E7�#��2^���G�[hi�����	D�RV)���`�����h6��oV���>�D2i��o��>D���O{ۃ�4�"��z���(������ĩi]k�m�Y����q��Q���_R9��,��E�^Z���=elʹ1�ȳ5o�L[�ODp]xchO��m�^���K<��{y�fٻ�qv���&eS=W��V�Ȯz@lN���<�Z���=��k��G ?¿~���g^)$D��"�5E�Ì*'�P!���e��� ��T3
�P��̼���j�����[�p�>ZgE�7�Z6~M��l��TE�$'��s��<���(j�9Ǜ�л=�B��n����|��gV{X�4)�#d�X.�K���؅k��1��\v��,w�\qnx����'�iN����`�ބ��jQ^�W���*���(h6�;���s��uO	�N	���o���M��MېUם�#�~=r��I|�D@�^��Lp��1'W�P
K�&�|�J��HWڐA�xF)����j��ɕWr]_�
^yL���������H٠ߵ�8]�L0�8�ֱ�5mŌ*��61�KE�s���>�U]6���Y7�+����}�Lq��QĢW��ݥ�������Q� ��mӢ���&�P�¤0�s�p���xp.*����� �R�Z�nC����ۑ���x�,uT��I_h���Z_�1,��/o�p:����x����F͕��cw�ط��y:c?e�2��@�L/��6�����FnN꯮"��s� ����AJll��ɮ7�O;��ɰROurK.z�Z+�6c}�Z���]uO��ӽ���@��߷��ѼtnII�7�\ٔ��ez����۵x]Ieƥǚ�Ph�y���T� ��+�sz"�)ߺ�ė�J��.4x~�"�q�s6cM'A#��t��A%�}|i~�4nV������/�;4�Ed>������Ⱥr��.�{HI�]�
��v�B"�w�ß��p��k5qƴ�$�CW�����h�M��i?4�;����^6kZKx"���	atu��HS��ʉ��`�r	��R�؛��J��A06�e/�����I��G�wt4��#��b��Yթ}�W	3�S�gw�tS���>�t�v��B_�HS o��6��¹H�(}��x!6�k�:��`�![C�޾��|�9����|v�e�>A)u�ϧ��X�����Ϧ6t�G[a}�kV°a���Z�����c��:��_1����(�^�Ө��neq+J�{5�	\��CE�Ҥ�.��Z��X>E=q��ˌYI=�E�ms���Հ�A�
�E��	���������O�E�2�������_�E�q,�f������e�d\�u��mZ�uw�kA|���a�����Þ���r�}��2��v[$��w0���+vV0��h��=_ }|����A�<�ED/�2����*�d]�,j0�. �je�h�SU����J	�M�)�T>�6�4P���ov���m_��bE6���m��@����Eg�)�����a���v����I]xX���~;�1|�-���8�C�
sQƨ���}F�����+���ǹ��ȸG֕�\Oϲ/+g���ٻZ�U��h�{$L�ϴp3E�9�fs��z�KI�E �/��5��01REfc�!#D���g� "��|�	��E�m���IV͊��gΔ��u�$� ���^ƍ�$��O���u�@��sD���R�����?YNbJe�$Ɔ��鄯�ϣ�^�kh3�cc������7tF�����c��1�)��4vFǌ�ODb�����!�SVh#��o7�4
}q
�Uj�j�����5�9ecٸz�TJ���(q�cF^��Wy���J��O�{�\9Vn�~ž +��u�b�Ң�ŭ����YO2�9UmGO�`.|��E���!(�M-@�O�PM��Tg������p���K���h�R�%*µ���Kz<��ɉKUg�:J$��i�X3`<>y>��})���#a�щ�U>���韍|�#�̻Q؏3�Ն~���T��8��'o%+�e��m;���{1�XN�E�U"Vlr��1v�����v�>�i_c�K�;������흫?�?��'}&z]z���� 8O�q�f���d&���u\���{9`��4��P:�\+u��8,5G�8c�d�g�ə�ڌ�c�
���N6\��N�ia�u���M^���B�G"�L���|Vy��Ͱ��4�>���a:�x�S����)���uNSXs݄�OI��0�)�U�e掺��lH�$��? ���1g+wǹ>�A+��h�o�s�����=,��t�d�[X7�6�3�[:Re���=�.��>������r���"����v��j?;��3+�t�J0��bw+'��X��y6�憓��;<5��\��`��ێ����4%�3�Q�s�!џx��C�P:���~D�X��/�TY��_�a��_Y���a��)w5UUA^C�a0�JʵP~(ק_೺�q_]�lP�1��L���c�}Q�`t��0p�+`�<��d���'�Q�~���^� ��B$3��������AS��"����7��7v�mJ>��jt\Q��`w/~�ӌ]�j@H72F������9s`�La��OP�<�"���3�J���t'B$�X4��Lj�k�W!�(n���Cb�����*U�_牏*��]@c��#�xuM����	�pZ�|����\e�����xl��]}68�^`I���4�(8F���xP(O��u����=�Lc�r]���uM�%�#F�C�Ó���B T�eҡOLS��H���X_��sD·���S��(47�^���hc�<~�x�0���۾�;������������r���Yf8��a[5�T CBݷw3�Fo��J��w�~kd����}�s;��iٓ��w�^؋�w�jh��4�Z�b�͇sq�R�s�E���"���#RȒ�~�`n�OR��v���n[�H�"�3J_"���?z���S&�O���	�{�L��o3=�#s� -�aY?a�K�� ��̨>.�G��ʌ�J8+�s��x�8���B#!��}�fN�&�u.��D�/,!�����p_yi�c.���:��E�w�0�ߦJ7@���R�}��W�<g�9,�����5�O�e&�4eԲM�-��;X+��VI���;�����8�rg�ް�j=Im5��$V��`s��.v���Z%8|efCp���������h�Q�"���
�u�I$�ݢ(�9!�r�m0߲!d�-o��]�PQ+"�����9�>qp���"�e��ͫWD��7Z���/m��e&�Y���2���9�@)e��z�1��Z�_�djr�d�3���S������.מ�1����Fa��	;ʔ����Ed:�9D���F�