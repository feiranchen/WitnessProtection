��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�ƶ�biA�9F�k��c��A'^@��l�����k��+��4Q���_�1"�9�ц!����7qV�+2E$�m@5B[Mrz���;�Q}�*�4�/��� ���@��PI釋�Vc�r��j�Ƒ�1�h)>)՘m�hwO�ߔ����'����D�!�����*�|�pq�Q�2T]���t��)9x�=����Et)KY�86�R9v�	W\rEV,!p���R�`O�����P�c9�F��-NJLYO������y�J^.S,��_E�^�������hrk����I�e���~Tbݰ�48r�5�����)옦!9[� ~�pb{Кq��)T\��V�4�[_��A �=��`zX;i R<K]y�ch�� ���ԧ�K׶�D�2�&א���.8#yRD�Zm�O\�jiư}��_�o��G������8%�'��%�4�����c�OJ��1���ͧ�]��� ��8G45�e�G�UHT�v����4u&��Q~���<.D�y�a�Ej�1C��jI/;_���6���t�B(��%���쨓�y�Q���o(�#�N�g<����AK�ǂh�X!�͹���s�D"g@Y����:"u�y�)�<� J�&�v�1�ɥ�:Se!���g��I�'��|�k9�M>#~خ��$fYf���4���x�Sg��dIx�R�t. g༏+���ǝ�OE1=dd��9p�ղ�ߥ�&Ԫ�i�9�H]+��*c��9�`�7lǎy�W.�����8��
�������!KjUE�}�T�2f).�'��y�h�n|���ǁ˕���I$C���1~��)9]K9JB���mZ�=U���Zl�p��z�U-xsT�����Au�;�T~�k��R��8���<2�o��uM[�yX��D�~��H}�R��䃃����S
bUw����
�4�7l�y��z�d:�Kf�����-��r�,dB�L�;�s�@������sE{������v�ėT �׸0�k�бb;eMc荷�����"���"SQkmXmCS+xt�w=S�p��Kv�;&
�B��\��شdu��>~nEQ·���^˱�ɷv6���[U��e��l�e��-K*���:��99)�}�w�)��e�OQ�bXt�,lqݟ���'׷/���?PIE��xo���lh��+��:<��V�2?7��9�k1����r��Q���ڹ�G��MFw�2UMW'2b]�,-��BLz�Gs �}4Ͻ�M�'ɰ��/>ӟ���㘺@ں��a��\^���	p��~���z`U�+�n�`f���ı�@���L��>F�SV�d�fE.��%g=̼���IҰL�0�ͽw��8WK�<u��<D҂
Ҟ1ԕ���B�M����G���4�gUF&�7C@ώ`
�@��sG["(T~�ǝ7��Q���ғ��v�7��9>/)�C���(P���@+~����4�]k{��ҩ�V���T��TV1ú�p%:jߕ*�%��F� �Յ��k��{��56�6�0����T{�$g��A��5Th�@��kC�w�._Z��޾�:��ɻ�W���Dx}vR>�ݖ�į:�J�ą��NM�`)���O6�BW��?'M4��Ü�dN_&q��D��2�;��Y'Enj�@as�lͽ��J�z;�FƴZ�����ȒMAt��u��Q/wb�&�_6��St?��B��b��S>F�C8�O�&J��\��s��u�:>J�7V4o� �"3��n����hT��6��d��Vx�K�"p��s�uh*,�#��U��U�r���(Mw�m�����煡H���g�١�螂]H1|!0��b� sI�����
��	���}�ҳr�֣t��8M������+��{{،&q��č�-T5�V�vbK�;���� u�����F�\?���Y�X��?�Q�1����`U�aݡW�1*	�^��d� @`�k@� ���H��W�c��VJ=0c�Z3�����UA"��`n����ꁖu����,��,��?�ËW����pq=��f���Y`��5���v��lǌ�?p�MØ�7�B��V��x+!�y��f��W����a���q������L9cv\�XfS�VWN$qN;DHO6r��5������X�[a<q�z��>��h.,�o��H�9�%l?k���}�~�IW��|NUE�x�����nvv{T�S��~� �q���}�Ȅ�/�$�,!L�"sS�S?�>���[��rV.Z˂7�cr�h�3J<�0h�%՞���+1��T��(�V��f<q�KTnu�2����bx���w�]iJ��a[���Ef��W�ˠD|-|����v$�$��Ӥ~x��HBY�{,s�?���{!"�ZƟ�:�CЉ��>�M���x34�RX>v�(�y�J��dk*�LzkˎF��,����
}�N���D�.>����V��W2�}���e����P�:k{�̸�}�􉍢���&�
J��Y��nFH�˶{������H�����Y�߽�д���&��~R�N��]���l��7��tX�hzur��F�!"��Ğ�����A�Qf¡,�$s=Ȣ~�V���}�k*�).?K΀t\�|�>(.~h,�
��X�儡	��u0���[\ ��$;��ow����lr�aa���7%��d�,!_��[տ�P�&���u~�eɁNu�U�aR�~檎�����P!g��4Y:�Luw�ـ^a_Ѐ,Mx���oLB�P��wͪߊ�����\���Y8p�	�{<��}I�W��(ۻ�ʄqW�iT/P�/�v�ۚH��������_m��,����`�t�����w �y�g@#>��|��s�C�8����Q}�������%�5w��œ�6;�%:q�c��鞦Rʷ����'��Yb6�l��!��W7�
�]e*V|,k�$��)3^n�0�zDz)�r���e=�Y�5k�բ���=�r�þ'S���:M�Z���S�����an�'*1A�
ͱ��v��z�'GZb� $5���u=6��/C��۷C!Of�L�0���3;R��{5�@-���D��4V:`�%���&���Q�ys�J	k�cOu�5��Ӆ��VM��GҌ�U���n�QMTҩ9Fss��W�^lE2��w�NZc�R�,��,�J<�ٹ�@�`O�B\�,P�Nt�����#��x2ɛ�B.M��.��l�U_S9�{t� �&Ʊ�s��))m��K���b��t���{�'T��ٜzR��C����Ⱝ����ax��O�\(�?>~�I��b�]�~ٮ���#k��>:m��:.$TwN����C쥝N�#�k)ng�R�aY���`��K�[�o��z�-
M�Ç�&g�h�y*���w��3�l23�X��_�	�'t�!
�F�I�>�JɄ�T��E ����<&������C�qc��ϓ��cHW���6 ������t�a�Y޹<5�	lp��(�ۛ�_���~i,�9"O�\"��R�̜mu�,�vZ� ubg:jGqi���K�05�E=��e���Sa�O�f7DE����nk������g�zP�C���zԃ������U����<j� U�:^�5գ�.?�	6T��B&���&ύr}�,�4A�'�GR{�t�W)����x9�p��� ����J�=�A�������I�c&(:�qy�4Q&Ϲ�n��7iU�2�B��jRy�c;i�n���r�vL@Y��H֌�Z�D�����1N�W�IVC��0n�yo�ӄ��V|)ʼ�{�J}\Y�$��"��-�p�e��C����;q��ؤ�F�J�)�	��tm�<�xTvif�L��k,��(S3�h�,XTFU������U�8�b���E>/NI�cP.T�[���X�rR��!H?ba�:n��L�יA+��~]��`k�h*�)q��Wb,��x�5a��7�b��=�}���>�V�M�o�T��J����7�����f�����=�S���1�N�S���z�p	6JCfN?�2�e</tms�@8L��X���s{���w6jWV�X<�b��0�+I�>״E
��i����jj�V�hv_���]ۖ"gV,@���"�Z��U�]�3r�+%��8�yl���~��hT-2�t�o�G���XJ��<���^u�_I�ڻ�C';����)��?@�x���E�	�A���Q8��4�^� )&{j[z`:�ۢ��%X~��6W��v;8F49�]4�D�H��]b����n��3��5�C�)sm���R[d��D������̖� �C�Tg���?�Dq�p�nzW�B"�sq��T�#m�<q<�>6����
Ur��{�D��=���|�}ߘb�G�s|9��*�V��N�n3PD�M�S��3�	j��-{#F�vU�ТA+Cy{SYMd�s���z�Voi�$��bq6�4{�B%ܤ���l/�x���X���IY�6�&D���Q[4ENIl��~�p���N?��O��Je�<���A��|<�_Se�>�G���=�D9J�#�bh���Ҵ��s%�0���
"�`��ߞ��`"���vjom��J+dH��3*��uu��a�E�̵-�����<����B�|�� ��`2i���8ᨵHe\h���I�OL�Ͳ�!�Df�P�8��{�6��$�yː�_�����]�1��|�;��v� Y@�)s'�u�Qh�1�mp�Ų�Y|�D,�R:��0�W٤[oҐD�f���\��bxRD�bW��|�qV|�|/���8�� }���o`�,�X�(
�Zi�Z���{S��R�F!)�;k��#��?nj^H0;������N�Yuʱ"�a��:['E�����0C��G��͖�����#R��	���:�h��8�[�z�Ϸ�&>���o��US������;U�*ꤠ� ^�-v��j0/@����' �Lc�!�3R�|�0~Յ��]���H@�Rk9�:r6x[�~B)��p�@��ZdM�aTܔn68�+�\�/J�,\'1>ʌ�����@~��O�kB��O�\�F4n	=���a!�6J|_�G1��Q�R.m��⿚L+���[!�yEl��a�`v��"l�0O�Q�;