module win_lookup(clock, address, win);
input clock;
input [11:0] address;
output [17:0] win;
reg signed [17:0] win;
always@(posedge clock)
begin
    case(address[7:0])
12'd0: win = 18'd0;
12'd1: win = 18'd20;
12'd2: win = 18'd79;
12'd3: win = 18'd178;
12'd4: win = 18'd316;
12'd5: win = 18'd493;
12'd6: win = 18'd709;
12'd7: win = 18'd965;
12'd8: win = 18'd1259;
12'd9: win = 18'd1592;
12'd10: win = 18'd1964;
12'd11: win = 18'd2374;
12'd12: win = 18'd2822;
12'd13: win = 18'd3308;
12'd14: win = 18'd3831;
12'd15: win = 18'd4391;
12'd16: win = 18'd4989;
12'd17: win = 18'd5622;
12'd18: win = 18'd6292;
12'd19: win = 18'd6998;
12'd20: win = 18'd7738;
12'd21: win = 18'd8514;
12'd22: win = 18'd9324;
12'd23: win = 18'd10168;
12'd24: win = 18'd11045;
12'd25: win = 18'd11955;
12'd26: win = 18'd12897;
12'd27: win = 18'd13871;
12'd28: win = 18'd14876;
12'd29: win = 18'd15912;
12'd30: win = 18'd16977;
12'd31: win = 18'd18072;
12'd32: win = 18'd19195;
12'd33: win = 18'd20346;
12'd34: win = 18'd21525;
12'd35: win = 18'd22730;
12'd36: win = 18'd23960;
12'd37: win = 18'd25216;
12'd38: win = 18'd26496;
12'd39: win = 18'd27800;
12'd40: win = 18'd29126;
12'd41: win = 18'd30474;
12'd42: win = 18'd31844;
12'd43: win = 18'd33233;
12'd44: win = 18'd34643;
12'd45: win = 18'd36070;
12'd46: win = 18'd37516;
12'd47: win = 18'd38978;
12'd48: win = 18'd40456;
12'd49: win = 18'd41950;
12'd50: win = 18'd43458;
12'd51: win = 18'd44979;
12'd52: win = 18'd46512;
12'd53: win = 18'd48057;
12'd54: win = 18'd49612;
12'd55: win = 18'd51177;
12'd56: win = 18'd52751;
12'd57: win = 18'd54332;
12'd58: win = 18'd55920;
12'd59: win = 18'd57514;
12'd60: win = 18'd59112;
12'd61: win = 18'd60715;
12'd62: win = 18'd62320;
12'd63: win = 18'd63928;
12'd64: win = 18'd65536;
12'd65: win = 18'd67144;
12'd66: win = 18'd68752;
12'd67: win = 18'd70357;
12'd68: win = 18'd71960;
12'd69: win = 18'd73558;
12'd70: win = 18'd75152;
12'd71: win = 18'd76740;
12'd72: win = 18'd78321;
12'd73: win = 18'd79895;
12'd74: win = 18'd81460;
12'd75: win = 18'd83015;
12'd76: win = 18'd84560;
12'd77: win = 18'd86093;
12'd78: win = 18'd87614;
12'd79: win = 18'd89122;
12'd80: win = 18'd90616;
12'd81: win = 18'd92094;
12'd82: win = 18'd93556;
12'd83: win = 18'd95002;
12'd84: win = 18'd96429;
12'd85: win = 18'd97839;
12'd86: win = 18'd99228;
12'd87: win = 18'd100598;
12'd88: win = 18'd101946;
12'd89: win = 18'd103272;
12'd90: win = 18'd104576;
12'd91: win = 18'd105856;
12'd92: win = 18'd107112;
12'd93: win = 18'd108342;
12'd94: win = 18'd109547;
12'd95: win = 18'd110726;
12'd96: win = 18'd111877;
12'd97: win = 18'd113000;
12'd98: win = 18'd114095;
12'd99: win = 18'd115160;
12'd100: win = 18'd116196;
12'd101: win = 18'd117201;
12'd102: win = 18'd118175;
12'd103: win = 18'd119117;
12'd104: win = 18'd120027;
12'd105: win = 18'd120904;
12'd106: win = 18'd121748;
12'd107: win = 18'd122558;
12'd108: win = 18'd123334;
12'd109: win = 18'd124074;
12'd110: win = 18'd124780;
12'd111: win = 18'd125450;
12'd112: win = 18'd126083;
12'd113: win = 18'd126681;
12'd114: win = 18'd127241;
12'd115: win = 18'd127764;
12'd116: win = 18'd128250;
12'd117: win = 18'd128698;
12'd118: win = 18'd129108;
12'd119: win = 18'd129480;
12'd120: win = 18'd129813;
12'd121: win = 18'd130107;
12'd122: win = 18'd130363;
12'd123: win = 18'd130579;
12'd124: win = 18'd130756;
12'd125: win = 18'd130894;
12'd126: win = 18'd130993;
12'd127: win = 18'd131052;
12'd128: win = 18'd131072;
12'd129: win = 18'd131052;
12'd130: win = 18'd130993;
12'd131: win = 18'd130894;
12'd132: win = 18'd130756;
12'd133: win = 18'd130579;
12'd134: win = 18'd130363;
12'd135: win = 18'd130107;
12'd136: win = 18'd129813;
12'd137: win = 18'd129480;
12'd138: win = 18'd129108;
12'd139: win = 18'd128698;
12'd140: win = 18'd128250;
12'd141: win = 18'd127764;
12'd142: win = 18'd127241;
12'd143: win = 18'd126681;
12'd144: win = 18'd126083;
12'd145: win = 18'd125450;
12'd146: win = 18'd124780;
12'd147: win = 18'd124074;
12'd148: win = 18'd123334;
12'd149: win = 18'd122558;
12'd150: win = 18'd121748;
12'd151: win = 18'd120904;
12'd152: win = 18'd120027;
12'd153: win = 18'd119117;
12'd154: win = 18'd118175;
12'd155: win = 18'd117201;
12'd156: win = 18'd116196;
12'd157: win = 18'd115160;
12'd158: win = 18'd114095;
12'd159: win = 18'd113000;
12'd160: win = 18'd111877;
12'd161: win = 18'd110726;
12'd162: win = 18'd109547;
12'd163: win = 18'd108342;
12'd164: win = 18'd107112;
12'd165: win = 18'd105856;
12'd166: win = 18'd104576;
12'd167: win = 18'd103272;
12'd168: win = 18'd101946;
12'd169: win = 18'd100598;
12'd170: win = 18'd99228;
12'd171: win = 18'd97839;
12'd172: win = 18'd96429;
12'd173: win = 18'd95002;
12'd174: win = 18'd93556;
12'd175: win = 18'd92094;
12'd176: win = 18'd90616;
12'd177: win = 18'd89122;
12'd178: win = 18'd87614;
12'd179: win = 18'd86093;
12'd180: win = 18'd84560;
12'd181: win = 18'd83015;
12'd182: win = 18'd81460;
12'd183: win = 18'd79895;
12'd184: win = 18'd78321;
12'd185: win = 18'd76740;
12'd186: win = 18'd75152;
12'd187: win = 18'd73558;
12'd188: win = 18'd71960;
12'd189: win = 18'd70357;
12'd190: win = 18'd68752;
12'd191: win = 18'd67144;
12'd192: win = 18'd65536;
12'd193: win = 18'd63928;
12'd194: win = 18'd62320;
12'd195: win = 18'd60715;
12'd196: win = 18'd59112;
12'd197: win = 18'd57514;
12'd198: win = 18'd55920;
12'd199: win = 18'd54332;
12'd200: win = 18'd52751;
12'd201: win = 18'd51177;
12'd202: win = 18'd49612;
12'd203: win = 18'd48057;
12'd204: win = 18'd46512;
12'd205: win = 18'd44979;
12'd206: win = 18'd43458;
12'd207: win = 18'd41950;
12'd208: win = 18'd40456;
12'd209: win = 18'd38978;
12'd210: win = 18'd37516;
12'd211: win = 18'd36070;
12'd212: win = 18'd34643;
12'd213: win = 18'd33233;
12'd214: win = 18'd31844;
12'd215: win = 18'd30474;
12'd216: win = 18'd29126;
12'd217: win = 18'd27800;
12'd218: win = 18'd26496;
12'd219: win = 18'd25216;
12'd220: win = 18'd23960;
12'd221: win = 18'd22730;
12'd222: win = 18'd21525;
12'd223: win = 18'd20346;
12'd224: win = 18'd19195;
12'd225: win = 18'd18072;
12'd226: win = 18'd16977;
12'd227: win = 18'd15912;
12'd228: win = 18'd14876;
12'd229: win = 18'd13871;
12'd230: win = 18'd12897;
12'd231: win = 18'd11955;
12'd232: win = 18'd11045;
12'd233: win = 18'd10168;
12'd234: win = 18'd9324;
12'd235: win = 18'd8514;
12'd236: win = 18'd7738;
12'd237: win = 18'd6998;
12'd238: win = 18'd6292;
12'd239: win = 18'd5622;
12'd240: win = 18'd4989;
12'd241: win = 18'd4391;
12'd242: win = 18'd3831;
12'd243: win = 18'd3308;
12'd244: win = 18'd2822;
12'd245: win = 18'd2374;
12'd246: win = 18'd1964;
12'd247: win = 18'd1592;
12'd248: win = 18'd1259;
12'd249: win = 18'd965;
12'd250: win = 18'd709;
12'd251: win = 18'd493;
12'd252: win = 18'd316;
12'd253: win = 18'd178;
12'd254: win = 18'd79;
12'd255: win = 18'd20;

	endcase
end
endmodule