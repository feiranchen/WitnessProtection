��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��x���y�5��mT՚����&���8��������&��!�&(�	�[��W���%J�E<N�K'� ��I� `l��7c�2&�I��z9	��c�G����wL6����҅z�:,?��~3t�˷�p+OX遥�'�l���l� |C*J���{Hox�^'�w��4"[yt�|��>���<L���l���b�����.���>��}�5�C��Z�ʱ��������r�θ�����%6l�f�|,��j�Z���B���������jf�$�.�t�˯�W[���q���� :�v���~}̓ڿKs�dnwD�y�C�N+�o.�0x�#�4������x�NjS�~��,"�	�Z�U�=�F���N㏍��p�ئ��>����@=�rPХPa���"(�7w�i�:�HjB���Y�Ob� �Z}�tB]�R����Q��-���s�� L�������w ��-6�|�G.�����>��wbR,�ϥژ|U����*����T�'�MQ�"�㘭��\j-��=1�L�j�v���N���(�H0�k�V�J_�2��������SM_0��G�^�p�.#G�I.�׋zF��?it+a�F3+b�)0}�՘X��3ޑ¼t�0t�QZ)�t�qmN���W���֖1�� �V%G����KO���+����	���v*!�xG������'����.�Լj�US;�8��s�Jm�JG��b�:	zN��"���u"��10� s3�)�ݘZ�Z���R(��[��l�l�,���x~�e�i˘^"���1~z�Q�s��e�H��qQD2� e(B���B�Y{	ɏ__��7��ˋq��'��Qא�>Q��I���926ŤK�q��E���'_�>'��c��f:;&H�Ȕ��鬊�]n�}:��%�ȐͲZ�	����TO ;�)���6N3Eω���Cd.p΁HB�6w+t���dk�KgR���"ܫ��yb�Ie4%ʀ��4^2���'�ۭ<=��zװ6Y�1����a��A��P��F5���>PzOTݶE�K����,�l�b��D�>�5�7�a�:f���(J�`����0�q���@��/�NR鍕&r��΀�91(���^���U�ג�ЙDӯ����y�>ל�ZrU��T��_�\�HЍFQ�DL�l%+���$Xd|�T5���>��}��W<�^��8Z˲��ͦ��C�݁�#��Vظ$:ޗ��dh�Ņ+�0�l:%�nr��L��Đl���mY���9]�%���7�1�Mݗ����HV�/X�F�b�B!�