��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�AT1k�:����-��kQ�	;�� ����z+�g���ܸ�6�#zx+��*y��IA�=�>��Z�A�����yDS&�\����� %�������))}�>��4Q^Ճ<C��d�%R	�col�A^`�(S�>���^�����o���.3�ڊ�r�r�x�i����ʠ�]v�I��M��u�t�
�[Z�sf-K�X��w�;F
Ā��Q�Y�e����i�5�k�@v�U4k���5�r�6u�;q�!,?�)��M���TwZz
WY�g��}�M!�wų�y$����R���c���4���" ̫��9;��C�-��w*L�����E[��Ӟ+�䘭�Y�Z� �o�����������_�p9|=M������G�C���7Ж���YknE8��+���l��$g�>�Wo�Xˆ\��@�ʹ0�:}�͛~�j�q�y|o
�+�?�v8N���a�O$�;� a4؂�&�v�����<�Yr�a-��p�ǩA`��� ��0����s�R�X��m�:�6*���uO*~!��I<��B#MLK
lG����Q�I��I�XA?�dq��k3�ӵkn���]Z�O�y�=��O�:�{Iё�*( ~�%���A>�g���C瘔hރ���bi�_���^AC�����,��6�qk�w�\�\���lѸ�=�U��?��]�1k�^1��Z���kZ��dQWk6@lA���p*m��!��>u��ɯ��M4�o����;rdA�:l�'�����W�1Aϥ�
�����"��<}��)qA�8��6�G{r�FS���ut6��Vv�<��_�?	�K���~�������e=��ޚ�u�}��o��}S������ҴT��i9H�.BfĖG�����1���� �7�r@�_>JFCvZoJ�T�j�ʺ_�;�s&��w�5��������Qɇ#� .����nK��zS��k����>�Q1�\�8���턔;�է�q�j�H<��T�m�=M���^��*�g�9��f[-���8�97���>�$�6O4��	����\�2l��/�XR�]Wg��ƅ8��.�|q�L��i�[d,�ū�)\��ȅY5�!zW&[�Ж�8l�s�  p���y�w��1~�'c���j�{.7/e!��7�8}�s�J��H�W��p�2�ҥ�`��ǧl�cV�f(i�~<}Z���U$=2�ٮ�H{z���ГhC�.�������_C�?���]C�ONOAr-���.w�,
�)��&��w08??.q8H
��Jw�~qNF�C1�jn,yb�����I�3�-���N��k��#����ng����NG��*�`
��b�\��R��T���Cp���^��h���n��T�?r%yF�)��m(P"Ƥ�.���I�7����C�JA~t(�o��Ĕyr`���h>#��ר��t�b���z���z_����1�����R'!?W�W��V�n@PA���R��k�p�a�^��Ovo���� Ε�3�?	w�N�d��u!ҫ/�r�DSa��q|l�%��w��2��YPJ8��y3�J�.�����D!��!�Bg���9BT�Sl�X}�:_#u��~{���=;^��k���䅤�^�bxQ�Mػ& ��t�B�]z����?�e��Jv��1��$t�	=>�-?/��;W&�X�*b����[(!�.����p��u!�C��]��¢a|��z�ן#��k�7-U�X���/���ái���s��65�����	�&���_��,��=c�Z{U�,��h��c�!efN�s`��ٚ��X�R�Eҩ�U�&O�<�d�7K�M���oD3��L���UO���Hz4�H���ps�4�;�Bo"y�B��E�8<�I�H��YOP]�ЌFi�kL��-��-��F
��S���~=�m���O�*��u�<���@B�Si*��_�z��ы9�Y��?x����&��)��	̦��X8���]��C���
����Au�Z�#�zz��:u�^@;+�l(��=_��>�⇠��ߝ��s�Rr�:�8Dp�ݕ(#���+����rӗh!�6�i��������fF����f���J�����<!y� f�\]>����/6�.��7Kx \�Af��Ȝb?����cQ��~�ۜiv:���c�㹸�->�$���:J�x���&f���9>ܔP倗���[�K��|��Nѡ����m�y�P��j|]J�y=��8@*�KSs�e�t%x�{ĥw�,30�cG�{��®V0��ە���@+�iˋd�;��'�r%5G��q�8���R
1S�'|`CM��J��-+S��&c�)Ɇi��~,�m�P__U�O��*�폙�IJɻ�&x�rm��~�6�}[Wz���)e
�h����H�T쵓2�m���2hm�C��k�T�^�iG����#Vs��U�L�[�^{�BA7ׅ$]�����H-Az��;�8לl-P��l����Y�C���y�|�a5�`���q�-���B�'�NB�"���5���
/2�j���o%��`͐�f��;l�s̊(����:����W�&�-��x�&�,�� �� !6V��C0�����/���xL%�W�Qt,Ez�li����
7��!�tw$�W�'ֳAV��>��e��!�P|~�d	�oggF�� �+<�m,-������4�!L�Lg�\yjK�n�R��-�Z��>���F0%p���%�7.�W>���cN�ϟ���퀊�PW@��ٻ��\���쭢*�%���  (���ζ%��s����g˫ߜ�P_pE�Rb����p(��x�\X��O�M����rh���eC7B�J���Et��NKG���Vw�N��wW�/�;���;��#�L3I�/X��OYU�b�.�jKN�9k�u|�Ϫ�j�E`@�mF�gf���oV�a�_�M�O����6#+�J]��$�[Q�jڳy?�|9�2��҅w�M]��#��+k���<#R��L���0����ŸV�ȣ���U��?!�\�P�*�EP��\�Hx�3dx��`�7��w	pr9;�n��>����)���;R�X6������7�࿦�V�g���2��i�=��	w	g���G���r1w������	��!�*f)�����m�uT�n�y��I�켊((V��e[����K�*��~'/3�j��_^㥔�Ѐ�X-�"U��L�0��>wCfr�#s��,�"�2n-ee'�W[�*E�
�Q��0��D)����w(��۫��,�_�7m8���.SI=�䕹�����,����!��J�I��< +Z�v��}��oxRj��������6b�Jb�Y���.�
A�<�|*$��E��+�������q�a�/��ߕ˅Ī�:���/N8�l3:d�g�K���a�ȓ�����o��D��Ƌ�'u:d�Mv��{d��
�+ǐ�+�=�g��8��0 a]�Y�^�ﲇXf�+6��M��O�cu&:X�8��<�-�n�ł�΅��=�u�B��Յ�|ͅ� \i(��{���e�ycjN���2К���s �&���=�K�y'�>�;]>m�,�����RHyR���r�
�}�ܧm縌�ء�:]��h��:h��X��n� �ߺ��L�~��R����z��
��OId �"!:C�dv�Q�KJ��1��υX\|�����GG;@XԠVm�ӟ:��{܀�F��miZh���_�!�§X���f&�_��3����}��x�8k�>J� �����F��m����c��k!�OYn���A�w/>���(큚Vbg�[^���p$���)4QNQ1��YT���)���J�_���q�U�!��x)���ne��xt�'�2�$��f�c3����;���&u(
���@�c�˩�
��"�Z��x[A$h��Þ�r��2���H��;����P�/���&��Xb����jO��iq��;�.���b���=��eh��&5��\LM�Q������Q�J����������;$-AP���D�t0�d���o�D�Hʢi�Mr�#�Nr��?E�$:�0{�t�E��ϵ��ޤ��xl���)�t����dv>����C�����Ih�q�<eŠFߪ~��}?���,�v�T���/@s�zx��+!����U��9CQ�!@{������:ڧהՔ�O���}�Y����䓓0���w�19�C>�v� �W�v�-��D��qDέ*���bIה�D�i�U��%T�Tr�3a�P��Q^���� [�_�_a ~�]�DYw�PĠ��!"8`������7&�3�G(�-!Ey�x��4(e� 5��O�Y�4�E����悪h���Ȅ)����Z�I�~��nt�,��iԿ\8i��������~�~0|{WwJ��<�QJ5�]�aN��
�D�|
'��կt��ȣ�Ǻ�	$�P��[��������Jjx!�D��\�� Z û7��`�nj�4�>}�}�8��7wA�u�-4�����]kD"��x�ʹ&ژ�]f������=�E[�S�����'g��P�>���xt���#A�y��f��;<Xڨ�l2ȟ�/����y��u�c�h���r�?�z;�i��g�L|�"�)U[��D��1�V��!��|�4�B�@�
�,���)�ɍ��>4���'�D�i܇� w��W|�ۜ�1��M~"�%�m߶���b�O�ؿ��u>e��erz��|�R�<��Oq�^�%�Av-��9�-]�?�������Xe�a-/`Adv������̞�&�x��GT��ƕ�k��dJ� ;j"y�_�؇��cӳ4��X�8K�h���?�a������� ��.�Z�S|�_��4x�j��P��;3E�'^�Z��'�UbR_�_-�z��Hd�ܒu����1�D�	1������ɝת�^b�����P1�c�j6_�!_����{P��pU7�8p��JMM/�߂�����(�����8��E�lw�k_�H����,P�X�[77��t����m��!UP������3+c��޴j���;�0�4B{-~�4h����,�)����v�ߙ��9:�y�J<������6ғ��8��*>������G׸���F���e�gr�xr
6fi(>��Y=��K��9ƣ/�/��S���Xǆ�T�u�$�8�(�)��r�@9��?�#g-�U����xA�{����H��w}��	<�5�`<�~Z�M����3�h㟘��`K^S������Az0k��m���BQ�,�WC�H��
&�u�5�>���#�Fht�� ]�� �w�٣��il�!����[���)_�[�b/ ��;��(�Kg���f��VNc���%f��F 4276:��������O��;�ޅ�S}W��vy2qK��_o�ƈ� ?�|_B�Fl����c�e�DX������nE˒�Ʀ��c'ӏ�y���X�jU�p��*9j�f��miY�w�d���Ȟu������)��8�H5�IfCh^2���早-Y�'���N@�� �������4\-�;x	=I�c�5�1�Q]F�h��B���i} �ӫ!˽U�׉��w>P���ސ	����R��@Zu��au7
���\��W�t�$�ѓ����#���b�  {�в�z#܉�&����� l�G����!:��h$l�Zh0�+�,v���2*�%��s����
Mi��s��ܤ0­i-�	��+
>΁șU� gރ֩���ʥr��d�A�P�����1��r���o�8 ��������(!*O
r9�ę��4�;2&�0����H�;�-�����?��s�I�V���F�$��"�$��r"ʅw�V �XM�?�>%�P8��u��2��ܥ�"��7L|�mdB����C�^|-�/�.B_;=�DA��m���P�,Є�����B1�9rV���Zs������tu��!bug�}ԡ�l�(T7L�&1Pc��;`�\�t�,��Ȃ1��>!����z����#I���ƶ���/A�Wll�Y>G��[���K녌.>��1�p�2	�\|-k�r*���^�HhdK����ðN��vҦ�@�bu��M��;/��W�-��}v+TN����CQUxj�K�9���~2��*.;�[�kXsC��>;�+�HG�G���u��S�,�J6�`ѿ�	2F\d���an�:�o�dSD�Й��t�im�oZ��:��'4(�3�ڿSmw���\ts�
cpH��	�T^_3��&p�cI$����)�:H!ow�
�a���a��v���zW�+�ßR'��^��FHn�u��Y5V�n��j_�M֭݊�C�����VBV1�jy�k�ڻ1����<�/b��� ��w\��Ǚ��j�<E�%�0��	�ל���Çf̀J[��(1��]�Ԡ-�OF/�
��O��=��K���[�YnO��>_����o�n��ٌ�s�@�%���jJ��T���0����b�hb�u�WJ���]�;��~�P�R��=m�����q�k�BͰ����d2��V����J��sIq�"�4g]�v~�"������1ZMZ��~��S	X��"�w& � eb�0��Kna�q�Q��$���X�,װ�c��s�����K-��:EY_�1�S��_�:���XP��F��d4�P�>1}��3e��e��¼|��ZDV$g��f>f�۳����:q4j�G�n6���u\BUh�sU�'Z����fב6|}�F�<n8��ׯv�@�*��4���v��Nǖ���|ey�X�¹DM9/i���(�}?.�~�s���ӳ�Ǯ���B�)��6O��`8�)	��)C�<�y�߱ϰ�j�gȺ}��e�ĕ(�b��G�i^<��Õ�hS�yݡd�eފ�D�0�1t��g����@~#�P�,}�=�c�	��Ɓ4S�����3Z-��1@4�B�'�(���l�U��FN��]�s�^d1�Q:��R�WRj�R����)�>ƒ�(H�|L/M��I�a&�Y��}��4L��۠&8�C�D���+u����c]d�Kb��-*��Y�h�kdМ��%�1&��a�s�%w9lЬ1�;y�qK�V�+��5+�=	������jFvO�Lԏe������C�X���i���B�ˇ[g�6*~��v�Oq��I>��Uu�4������&Jɹ��+#%�I�����H;Tj�61��tA�o�J?n�f�/� ���$`*J��kG�L��H�!�R0'������;4Rx��=)�{��o��y%;�{�Y��ÒL6Oʪhj��;q��k��mG��ʏcr�G�7��i��G���4�))1�;�{�D�,8ts�����4g�go�9��!V--6�R	�X��\�x�ޓcU����r�bS[��8E�߈E�X��aiH28�$>�r�I��(o�:�7��-���Q��kʄ��
�=�2*�nUS�H��ȵnl�ۏ�	]���
�f�	$)��&�T�b��|V(5R�<~}���Ƽ8�M?j���'į�g�ƨ�J'V�B��zV��?ɂ}���u.�Z���6����g�G�+Q�Q!`j�2���K���[��8A��=_�/��Vy�6�
b\��8ȶj��J(��������i�aa��=���|*�����Yҽ!���/�I��^c���1T@��b^O%]I�d#g�2���F2��$�)\��,�:��Ddx Dp���p������w:��ӿPB8�4�6�]��T��aaOn����Hgl��m{E����>�����R��/ĖY�\� ?Dٺ�Bt���Y�,(�������h^��UX�--:����h���?�OH�Y���iJ�BG��
U�u�*[V��Ђ�/�4�	���_��o��гT�Z�<�B i``v"�9y�$:�w�Q�F���,M<1X�\=��qF���.S��� E��7�b�34�/���W���P����J�
�
�@u�gQ4���4\f�}�OU^8��[��a�j1D���Ҿ�����C�C�΃y�!?ɵ�����yU��-�f1���M���K��@P��� {�̗�j�I��Y�;��TB��w[/�#��k&WP�z���؁s>>�2�聽q��&���`�o7�g->"y(�Hý�-<���
�O�lJ8������))}:�	Y"��[���N�����qG�)����4�đ8��b����DIY��!�lZ$�z��r��T+J��AB�Ҽi�߾�.�cViW-�_o:j��83�����b*�������H�l�{��s�kF���>�'�0t�4�;eS��=*i��z�����"7�48}M&0p�2�+��e�Q��W:W���@^�^1D�˳�Ui%�G���3�;���'eL!�H)ǭ�P���~F��ap���.�@�m�y�xc)?�<�J�yU�um�ل�ȿ��ԑ��/z�[��[.��3��
�V�yn�o��=�����V"�� Q��d��dעV���S��=uE��09�Vj������0]�����|Ӎ��C��7|s,^x�lkKY�^�6׉�=�;6ma�&�NR/'!te����-u%���MaW�(���Ѥ��5�C�[V3�,��r]��<��b_2S�9�x3��ξ����p��C���myH�)�[������N~���g\��v�~��!8�P[�$Z#{?Z�ٽ{�&0��z&w��0���%�4։�$-޶����:�^����:��ǀ�(����P�{[���0��L�4��a�>~9����1֐�xZ��7�j�A��l�~	��g2D�Bh5pc�/�.P��3��圪��p���d&��u�����>L�sa�х �<8���#��J�q�!��ˇ����]���v�C�oE���.���ea�S�@�`΁Q+|@���P��c$���gh!��J�M6��b���=K�x���m�fz��N&�g9�Y�'=cj��X1�%ǳ���T�2�=/�x��OCb��[p�c�x�a��P��xY�-��J���@'��\A"��4-�l8Z�(�`�|��:R���~�IB!51���@�/.�e���Mh��md��oD9�&hk�m�Bz[���a.�b�3	�V�0��f�l��#Ir	4z���<�u��U�倀S��ߪ�dC�K�ITV�)�/)L W�}���d�w	\��چyJr4d0M��,[�[���y����[��Xu��t$��wi'��$�qu ���}�%��n��ۖL�u�>aP����<l�Af�ʎ��D)2l��,!����"$�G�BD�����cTd��~E1]ݎJx�����j�B{
��-�:�_�	�q�W�UJ�Y��TL�G����{����?f�,|\�Q(h��i��1nG�(u��{Þb�N{��'�����w���O��m�W��-
����A0�	�`
��`�/#��~�� ���$,�*�f���IQ����������*�18���!�o�_1�7%t��w��2Z�o��3J�S����M��
��ϕ��l1��Ҋ�����$���=_��h"RPR�D��&`���1'�ec:W��qn1<�9L��m@0=���E��Q^����?��PA����O���� ���p�-WZ?C���e!�s��8��U,MY�Pj�e�f�W�sr�t�������׈��1�=�`�kM��ϱzQ��U&%��v�.�T������ŬA�.��Y	Eރ���W��beյ�@]$9ƩvsC��a���U_�.Z$���T�q��,ڷؕH�MNv��;�VF��Z��H�^(֯�X�c��>�?N���"{���4~�bO�{h�qbk+6X� ����/���Å�?�X�6��֐L@/�>ΰM$۫��b����>�-a�H�0�^ݫ"�I��B4��l����{H��ZV���� �Ex��>eĕVR��Ƹ��M���D�R�?�X^����:T��[*f��3g+0H�̆�y��!>
��$����G3:+�A�����U���[5��_�7'�&����aP�R���,t�k�`��
<3kڎu�)��}��_���1��M����G�K�������� j�?��hXH���'�;�2~���z|G����� �ߺBjj:G�W�IbuShٸ��D��oaI��O4�vi���R����p]s�=<ϭ��#���I2me��&��vL��f�/	��s�/�M�����_Ų\`3��2�e�)����A�!>r�a-��3l���s�rh�d��F����p������RS�)T^D�s�"q�^���P���5T�
L�������9@yTn�qZ]����|���IIk`1]�Ŏ=��Qj���˴��v�y�U�me���h��5M�m�j��C%�JOZ�B���Q���tm��{���@������3���=��ǈ��kÐ�� ��Ӛ3�x��K�h��K�]��������P�-�l��0�S��ׁ`�e���&��J�p�/��thE�Ne�8Ո�G��	^(~�����!'(5�4�OO�2��Y��t2G�O��a��(�x�5�V��i*+�{���?�ɜ�?���� '��=U���s��cm
��բT�p��,D��/.=���U\������������u�q1WD4eɾY;|��_���$`d��Sأ�i��%:,:�1� ��m(i�V��ߵ�ĕ���1��l	��yD4�v�x}��ɾQن��x���2�h�:��8�봮�^݂�-�GDE�X4ܲR�I�{޴��)��u\����(�[���{{��řJ�Xz�-���ߊa��|���#�
©X��)�?����9��p
O9<���z#38�bݡ?�E��^��#j_�Ȑ�>P1�*
�&eW�b��x�w6J[�v���\<�Q-���U&4i�}�w'���)�ϯ!���#��U~8)U��{rA���aC!�[k���>B+��4'�G��2>���ʦ�4#�:I��y�?�V1xF��.���ť�޷�m�5�U��Bו��֔#�c	oj6�9E�i1�@w�n:����7�J�a�fD֢^0��Ly,�ؓ�,k�
�q1��mN��j�m��ש�hE3	�8'"?�$]��ܖS�`],{�X+�#O*��rw�k�W��,��d,���qL�Y�����;�8�Sb�J���$��f�2K�2�ٹ	�w���#��r��`i':��I�R6"S\��GĀ�
O0���@�f�0+�z��Q�p�o�H���LUk��!
.�
l�1�^\�mNq���^�����Jݬ`��np�.��~��_�(�ƍ\#�%�m4��ډ����x���m��렸��.0n�v�%��d��"��V:bw#�+�t���ࢷ�\�ZU��*�������+���U����gKi��8S���eD�cPq�֜F���_��w[d��V���U���CwY쏪 \e"�^� �{*rެ�b�`�j�K@C��ĉI����%�בA��{�+  f=�w�12��."���ƕ�{!��r�z��3����6J=-���Dƺ4��R���w��@���c
y[�u��61y�������Ź��l���.%R+2`�@))��F����*��>7��82��2��+h�&��U�.s5�@�BS�'t��w�K��Mρ����n{7yS�%����,w��1��\�*��K� !�$���#P�u��(0�c"���#�i;[?�zD=��OT�{���i����K@��Nw�t
�> �VP�v`����X��;�B� K2��r?zk	1Z���G3�@8�����SH�k�B��M_���̶�=�O�������bF��9
��$ѓs��v����4g)�Q��ݽ�Rsy��VKH�%2�u�?�}����Cthm�v'�l`�V�|4�@		�����V?[�3�wx'+I��'��/o����TƵJ�.1hT��hȾU�G\x������<%�[�!�֌*�LK�w��������Ք���_�H���׻��W�:���,��ȼ8��A h�M��N�]j��P�8�J����z�7��Ӻ�T8�O��c���tl�y�]Ts�@�����f�jÌ���>��>��zR�����8� ���;C8ߧ~_J��0�o�e��ׯz��b%�Uq�76#�� �_�п��X}����s��b@�qS�P��}���I�NZL�;�4 C���']A	�h�����w�IҰ��t��[Y��
}���B�riD�'��凜 F�Y�R&�ȠͮE�<0v��C��-�;�4��N�0�j��h��#")KS��Y��1�m���6,�<&N�f�
R�����"|�=���G'&[��X�ʣ�ڹ��Cq�'韼����@f3T��V6m�9Sq����~�7��z�]�R�����M�f��XV�c0aX�J��2&d����*aɮkvq��VA�K�y���
���lC�m[��ܢV�FТ�i�.B˝xw��#�~�Z���������z܈V�`"GUwa�Fmq*R=������16�v
Y���,o,��Ⱉ2�EU��l����{�Mc�j�`n�}/G�ۃdZQ��Q,�~�a�ʉ���g��/!'�1h��.�.Y�bRf���G�4���a� �c|>�� ���^�Ew�kZ�:��m;KcI��"E�7Gس�f M�ξ?{�vsz2���������辗-MB�r��P��ʄe��q����,�w���L�*f,LJ�&�,����T��l��3_Z�-kZc��Fz���^l���{�4l\?�Y�_�K{N���y���������_������j�d�թ��>�R}crpUs��O�uMq�J�
��RPs��'_�8�����P�WKtcis�p�iq�`�{vv�9x�K��g)�Qu=V�����f��N�J�F�z�f�X��!��Wr�:|K>����"捨�<�y�)������p§J9^�t��	���mN-OsvEI�/�[�2�ǹۅ�K���;��ƨ7�&�?��Å���j+��2�s-���HAw��A�(b5̻�v�͆�Ȝ�h���R
�{b�9�� � �梅�{�㙋���TT/�-ҭ.QЉ��?	�$=z&ɊC'��SP�k�GfT�=[�͙��,�Ec���5E@å�h�S<+�o-���5c����Q��ܭ��o���C��/��m�6�u���b�S������������)��
T�&M���à���P���ֆ�.'�Ur���f]HT:��r� ���pAh��N�M
҄vzB�,�6�<��k=�K��1=�9 2��0 u��1!�4i�i�Z��.��6@]$�t^��)�r�mF�z�:~�-2��TB;JM�y�Ĥ��*��;N�E���Hkt\�p���T6�cONY�*��IO}�_�35;���'�Z	&;vH�D�m®_r�g
2�[@]G�l!עX9dٓBC����Ac�Q=m��z���@r 4q��j�4P��A�
�E>�ў���c�7Z�d
��="���O��K�>-��7b�)S,(���j�
P^q��;V���z$u�3���o�RĎSY�z�?��n,����u��P���~�UN�f�T����}��uD�6D�i+f���l�Co���iŬ-�6����Xv	���$�ҟ��[�	�L\�`��N�]��[� PB����,W�j/.E+"�ӝ��a4h�0�I�3$�^�����6�;����x�{�ͤ6�H�Nc�ۦ'�ϖ8������������;�V��]�?�c��*<��G�J���fA��������͓'���|��'f��!E����n���]��;Q!����av�U���R�x@ �GF�x}�'��������9��	�	�%�κ��0q z<���/cP��Mmv���a��]0��F��B7T��)Qj��X�K)]��gn��\��&��>s�9������+�9��}f�,�
�܅;Z=_�6a��[��^o[��md�e8�%�d(|n�r��F��?�ҝ������Xs��t�\s�@k�����8U���7�G&�أP�A^�|��V+�#Ya�}@=t��S���M:�9��k��]�~�����wt�@�ׇ�=@J�	f�}"���;������Jn���H�2~����ed���l�$.��݈�)�j(���ZB	߃0,��Ɵ�0A~y���E��#.���|e�k��<\O��a���#�d�z4|�0)<�i�Eskp�,�ѣ~�TƠ6��I��G��O��G��K���|1�V�pמ��H����f��P�@���*��^����"Џ�ħj�=���p���C��Y��J���$[�X0���QV��]�u<q���[��p.��)�:Y��"��]����sy2I���b���/ls�j��#[� ��x�*q!
zY�B`]�O�v�5U<�W���A���{��X �"���B��K�&x�Ӻ3�	t�����h���qc��+7���o��1���3�)(�"�>�3?Pƾ��l���-��.&w��ۿ�W���T4L}&e�{Ú~��A-���;�.HS��#��}����P�0<��!y������M�.qj�*���N��/&T��7�'G4�`6��p� �b��C-�����BmmHUz��[�YB/m!0d����`ĸ�xW�l�6,�f��̉UK��c�}���%����Y����E�ITZ�q�7��M�T��91�^���z�x0� ��$}��f�X�4�!���`�ϋ���`)�dBokpwU�*n������>�|��x�/R�b�PӔ7��3�v_�res�W���v��Z�D[�)*�&R����-LW	s��iv�{�wCJXIr1=��FcU�j��~+'W����'#'�Pd��i�0��Uߠ����(�`�f�z5���W��S�*��2~�uՑ��b����V�JX���l�2�}H��T�e<ϼ��������A,K��r�A&��~�h���c�FKf�>W�2�ĥ�nM'<,6��$��baԱ�9��f(eF5^�C���!��a���V�C�ͻQcu��d�"��ɷۜr�춣�_'����m���v�tKҤ>9;���W�p��Ӧ)I�;��ZuWȭ��D�c�q���Cu&۠����F��|��4l��C*��h��wx޸�K��{G����:��<��C�Jk�~զ�##N:	(֢L�n��f]Fx�T���M��!IH�/��xL��?F:���N�aH�/�G��d��0'�5�e_r�'�� �X1vY���es{�wEnI�����P܇�B�oK;/�J��P+�	�e(P��k��78Ẏ�PԬ���<q= ��f��L�yK���R�u�U�������|�2R/�;������l5}��㕴����D�J�,b�*�.��?MA���2N�=ŗ��5���u���g"��1, ���x���^��X"�� g9�"� ��SKB�L�%�q���Ʒ��C�Xd�C��8j�y���~,)��S���
��h&f�&� �|_J2�s�vv��g���W��[b,d2���q�'u��)T!ޗW�r��:Ǐ]@��T����iI_У�^7���:ݦޓ�rcC.�@�1{^�H��)�{�m���:/�׊��V����%�;��ɒ�+>Ձ���>$9�K�t1^�ڻ�1�6��M�R�;ܶ�E�+AmT����vn�#�PEDmr���
�[�� ^���XdJ.�0.��-I�����{tF7Y�U�ӭ:j��Qnen~G#����;���ps�xu&9U�eD�}��b�U�	���jU����f�4����e˯���G�Sٽev~1J������vo��و0%�������K���
<6�,ޠ����ݰ�.�q��*��r
�z;b��T@�A���r�ł��0��to4��J�T%7�&��i�W��s�� �e��A4+1�xZ^1�}�Ri9Ͱ�ܜ7VE�.��. x��X<�Z	�Nvr�u��)�T��o�Cw�9H���̈����l�^.š���XB�ݐ����~O����M[�� g�@�"[7�x��4M�c��a%E����0�L�,��c���,�-�����7�����5-�|2J�c��8t��ߒ����ڈ (5|�:�~2+	�i����R��2e��I��U��ǋ���c;(�@�����P�]d]��z��}ܖ��|gdZ���ȅH&@�8]�E�Oic�l�ʮ8�4> /rW*1GW�C�N`�[So��팃��cp)m���Ò�*'�u���D��ϊ7�t!!�ꖁ2���.��">� P���q���R}L�{~V�N���l�C�"A��w��Pz�p�S�w
����~��̐0hXc�{h�����~��X�6�v���i^ÁLf��e��C>i��\ܢ��`��:P�ց�Y�����Ɲ�|�r�uW,{�ͣ���N�`~���L�����[Wb��͡(D��B"�/J)���[s(�4n��>���D6\ň$��d��_�Y7/��������p�c$h|��OT$Qx�p���p{oε��v\R��� "�w�)�S�&%rM�r}S��i�Є���0iZ�����u{�'r��)�]8�Z�jz�G:'�o��r��od���x��ZSi0��lQץ�/���1D;��`���G�p��TB�Gž �� �	����-3�#ג栗!{Q�|�HJ�R��?�����Y�u�/���gb4�z�}�жܚ=���6Ik���'���)�;zʜp�v�j.6�H�D��e���F[w����G�+'�;&qR���'��bL�ָ�Q{���x�<�ҧ@nb���h�%G�T_�.�{2�ˢ=��2[��>y��z��U�S��޼]5�S`̻\�|u�����������kŵ&�5�D"�P���X�`Fn~^:Ɛ��_��z9�O��?���=@v��o��_>X�g`ۅg����e���9t̖E���^�K�
��P�esgkg*�~ϩ��ѫ$��L�y���P�� v�/�12�Z�����o+����F�D�(�^N��pl��$�D@��"���Ć[����a�Omj߲��o"�>�i!wU0%�s�\D��9�4�Y'v~/Q^O[�Κ)�Y&��{[���7�O�O�4��3�/�T�A����s�'/���^Գ�[�@��M�	���t�n�m��e����)�'5�G�^�����S6�v�N�n��id?R��G?�]jy��@7uQ1�t�j�4�+W�D��e�������8�!����7B	�G��Z#��a�_�hP|��)���4�	�_KJ��8*�2\�T�^(��7f��R�gF�J���F�߻�.��j���26��ʯ���.F�;3 �A(�m�#�T�3��� �n�X�;3��?�����O�2��U�<�5Vt{��D����\��'5W~��R�ޤ�y:�?y=��<�<1����Άz�	Q\���|�$+g!J�|��=���+�
HdJ~n���4� nB���Ix��|��6��3��g6Ҍn�^��;�� ��w��f ��Ҁ%�\�u�}Q�|Qb���Ԭ
��xi����g�j�Ncg�+�l
�Z�p�V=�qj�aKT+ٍ��iy�=��4��Y�����O� %c�[m�\A�=(y�ٴ�E�wr���,=�Qa�$�<��m����:���g��T���l��c�&H���Ե�09Z��B	6�47��v$����=|�3�\ ,�6o��u�:�������.�"�G���� ��Vl��L|��'B�mQ,\| l��g���d$��1����lJ��H� &��sY5� y�$��0.n)��o�D�?��_.Γ؛	����N�CW���UJW�uQof�>IN�-��9n�hY��,�I���r9	�/^ì�@�;!Z�04"*W��ˣ��5�`>���1sw��a#�f�1~�`c���S��q�{~�p��y�t�`��:����S�γ��@۩�FL�n�XC��{չz�}�~���-_؇�[݋GN�4����S"E5=Y/� ��"�G�х��w��bI��[-�!����i]h������O������5�(�*c��tX+%���G��fu�s���[s'���D����\5�Sn�X���-L~zC	v� ��zgm�Q���i!y�rW�o;�5�81�%R }%Rcg+��{�R��SE�)��K����7�f�Qߦ���>q���)���Pk�I������1$��_�,�ZWI���k�G���o��1����nwY�ߓ�1�VW{��)�o0�U����a9BOՂ�[���2x�t/=)��P?'ə�0��MI��ty������4�2�0��� �y`��=��d�Q�S�� ��cK�W�Wpg� ��h#��[��N�w ��c�s��+��fj��_E�Q=�p�\��f�r���m�J���F5������Y�n�Xb�a�Ϋ�G�B��a����'��g��Ե��4�6�@�OK��r�(_���+h�Ӫ XEOp���L%�:���Oo�Ή�d�B_zeC��[�ڃ��T ��S4x��F����{���V��`�u9�=?�3������*�	�ƍtlYP�ߺ$���ݕ�m2�\U�;�بk�Q�
?�������0FW�4s�p�}o}�*�x`��DP�/R��%P)�����1�I0���y�sm�\@<��|��ˎx<:�˸�{���ҟ�Z�y��R���5���Q|'�ְ(���}%֌~_�5;���PrWSH��"-�/PS��<Ƈ(|Hi�g�b�~�_Q�K$5�~b����Q��^���J!����8o�C������W�SEIf��Y��rH\;�+pc��.��eѬrx%�˨��Gb<�o��c�?�@��^dN�rcF�aIM3\��@��믈L2�S��8'+�3��G�T\�E�өN�p
у)Z�$���о��'�w���I�����FD�FG>��V��,�#Fd��UK���0,*$k��F���/�%��M���FQ����A�J�Y[,��×S�VԦ���1���z	�Lt����Yڧ�r:���1A5Az5$�{-�����s�����	�^�b��-տ�{�$Xt6�*�	�;.󲞸CO���6H��y�[����H�p�
��"cI���L�~�F;BC��;���X��9#���#����ą6�(s@ޥo��a����\�?�b�ء��-�K����RP��t d���?����|�	y�	�쎔O�&>�c?��>8���Aw�����^��I��g�1�c�e���h�Ĺ�2�F���j8v���ed���{�,�-EB<��i
�{ 
/z1 ����j�.����j0TN2�x�� m����	�-r1,��K{�[�:�i�S��W�+������f���:���sw�R
6�$��(k�Yjީ��z	S��?.��䚊�sd�u`��xfC��x2;@O�s�XK%d�1����?���Y�?�����J�h�KǑ�� ��d��/�b	�Վ���2T�����@*��z
#zEìY�+���=�	;��uJ�]���U����x��=H� �<o����J�W��4��HV�'�!��r���A�M8c���������m񷀯�s����c�	�\|o�yLoL��}Q���$	��U�B~$�Ƨ<�o)#wLuƖ�OU�cKe
G�����t�~��ɪ�Y����,�CX�
q+�]P3����B����BA��Ʈ�=���H��^������:�Q�f`ք�W@�:��ez���U��_�*�C, |��F�֥~�X��ܟ)�Ə�P-�C�h�ʼʦ
}Z���T��S�^��3��F'�Ă�If;u���0�/|�ǣ��/d��la�M����
bCYg�����;؟ ���7���y��&oU����R�D_u?C��V�ǻ.}"��,�І��f�P�%~�>|)l���!��͚�S�Ȅ���K�ގ���Oͧ� ܶ!#wj��X'brJ�
f�G	_@8L��F]�j��so��i��e��R�(���e	{)��Y�6�%f^�ڐV$���Ρ,.�����yR�{Px��gJ�����i/9�*�"!�"��$~��#���@ �r2�\@�W��α(FE�&����M�����Wb3�������A�����o6�.x��0]]`X믱�CI�������G5Ӱ�vՁG����h����<ð�"Y�7����H	� 2E���oA��4HN�<k�:#�p��#;oD_�!o�TF�>�.��ಞF��9�ɥ��:�D���]��̞&"��*�;u�4d	GJ�'�r��gISV��`�cZ�Il�D���7���$خN9�BӋ�p��΢��i4?�R�Y:ľE��}��*L�ߦ�D�I}~h���䰉 {��,��Ȏl��J��M���#l����`�Z%c
�܃�J�"Ι���wDO)�L����!bݕA�|���5ʶ8cZ'��Z�.���q��PQ9^oϻ(�냪�E�T^\g��7D�e������3(���ѸkZl��Z�xb<�rP���&�zv٢��Y^�4��?T�?��\;)>%���64��V���@�G��Iґ{�����
��:D�"�T,!��Iv�Jݭ�jv5²\��qz[X��}��L�H�����ʍwtϴ �T� |l��b��2�m]p�@����8��Le��2�eBi'JI�i�$(o����F�r�|G7f�`i
p}�������kP����@5�����B��8e��L����̕�71�������**,G� �G��Y�&Kf'�5Ȱz�#;�媏EOy?��r�V���D2j���f����4����U����p�k#5>J��2(�)������H~�~��ؒ7q��DS'�M�ۥ+���μ�i}jT~|(���8�����]������m�;�Q����R�%b3������1[��1�����$��J\Zci�׻p�DZ٪�ڡ#鈒W��zU]I����J�ent��r�.���Կ3��D^�)aQ�i�x\D����`�+�G���"�=�W(/95��۬-��۰D�y �û�F#�S'���rȗ
��q�,�˝jc�@�g���"D���$#q�Kq'zo��5"�J�c�gL{K�#��KC�56��z�jݰC�eH�ٍ����y�O�κ�:���N{H��v8����ok�ݝ\�>3�B���&�'T�����9m��i������ �[�V�g�~��w�B�������A�)Lް�p���$*;�M Y�x��lw��PZ'=߳jA~+h1ms���gtg�+�'2��zY�j5�bQAo�����*)kX8[g*F��|9�W��[Z]�%����fe��cF��|04ߩJYk+�?c}s��9��)O<[��~oz�b��t�H��̉�Pd�&+dW$�D��x���ap}O�cz��kX���ѡ_�9�*��V9��NZVP�X�YQ�!�wQ��%��X�������"�m"ue7�*?��Ю6��Z�̵b�'�z"m��X���c�%��?���6ٻ�7��*S?��Fr
yx���h}���B��MHu�	il�Fr�B����Pdɫ����>IL�9�q���S�Ř�]�#N6�˧��O���n��kC+���ǳ~����C�Z�j%�䑈�
�z�\ς��k�V�r~��1�%?����X/y�aϒ�-���V�vm�s��2
��6m�U{��TP��8n��#�QX��,����=I��/�x�q����� ����ĺ�����q�0���i��H�ez+s�h��������&:'��w��v�X�)�K����������G�NwP�	L-�l^f�ӆK6����������J��/8�Q�{��;-��*+�,�"�V���.�j���%�U:��,�r���J���"���}��������v^�/��{�iI�4~_�f��ط�C��&��*ybo>c���D�2&@�����LN/��K���\S���j�f����� ;���!�ѷ��	�q�*��q���:/2p�%������?iA��17�Qe��4�����K���J��E\��:$"�kѺ�2�Մ�|ګ���o>IL1Ja�NW-)��+O'a�oC��L=?Gt�7�G��Rh�N=R���.��.v�Y�����<����s.�/�Ø}ό�tR˸k��\���/Π᧍���?ĸ��W�]��C��r���}]����>s�ʶޅ'h6���'�M�pmk�ߜ�%�w$U�5(3���(%͘A:p\~y�:������e9,u_oDav��ᣈb��l蛑��� �=�=�b4!p?�KΨ��D��Pr�skz/�;��Ai~J�gϪ�D��ؔ�h5��O*O4sr�#�'�e�:��r���B6aX��N?�x���͛��r�{�ReY:AR�Z�q�K�e_�C��9�^��6cі�;��Q(Z��ri� Gp�WP��1ؿ�!���Vm%�����p-������;<�F�D@�ʱ����Y?��RGP����49�{�1���U�É��-�
]�zD��R��i������Ǖ̴G/��#�ѹ�+ A��M8B�&c�G��ʼR4o�	IP@��x��y����ƕ�%"����xDu������]������4��9Z2����7l,���T
��_�X�txɸ�q��~�����㥶�k��X8^/ҷϹwL!X7�xҕ}�Llr��'�h��-wi��݉����y�91����l_���&��]�*{L��6Uy_��AJ2K}��������)�k������n�r���~p���jfu,���1����e"��2)Ε�O�t�J��}+�1:����ykK��
.1c�J{G���sdgw���η%��4)��u�[�:C�cps��p�АQ[��'�,���~���B�1uA�ZݩN�dx��j����-g����4�-v$�4�6�V�T�������/˳�iRl(�K� ^'$����v��m����߸I�pQ�k�������!�����c9\>�8�Ju�/�-6�sQ�H��f���2׈T;b�3&S4�Ǖ�~���>�9�Q��X�i�ܿ5�Np����c�}y��dGY8��2_��8��̦'.�֔�D�g��᙮��n#��s��57��̳I�
�S�ٚ=�S�5cN�)%���4�j��W�4�;�a�]�T��e����k�+FZ���ܦ9�����D�K����P٠Y�1����D4��|k��8����+�;�IcW���C��98����8��{#��"x˖;�7hR0��g]~O�zn�����ӹ\<��l���&m�v�=��UY?�_U��e���`q=e5�	��R@H�L��ϔ��� |�^}r���M��� \%u�+�uDp���KQ� >�LCdMd�=[g����-��x�,���������b�#�rja�'��,�p���|�9d�YM��pU��kx�s[J�8���X�0�2�ҍ�͚�^�5s|�ENA��"J��=��O��l�ҕh&�h�y��[/�6����sUf�1A"�I�[�9���8�k7���8�Y��#��o9�L�D$���^L��hE!��*�N�kU�}����? Ѕ��n����
��+�z�([��4l?�d����,e��|Yg�4��]!�eQ���ԇGK�T#5N�Y
q)b��]q^x�	@��]�����'�����B�����A_�+����X�ݻ܅>��W@���迺�T�xW��8��[�'�-�3Ԙ�Ulj��KJ��Z��)�s�:��:��%�Vش��1MY�)����8�yg�^��ȹ��h9���G��E�~ͺo>�ؘ���ב�����g��!N�Σ�m5UKV��)ң�z���s_���4��@�<	�GO��~�næq��T�G@��	<ⴹ�A�0�z�I�`�<Ndh!^���Tu	Mf�mқ�3)�w�b��X'��M
P 	�t��0���{ur@�\�����W�>8�Ұ�j�Uu[��?h�^~���{�o��^$g,��$�l�Q%�|A��Z_��r: ��Z6�cv1K��QU����`�ÿq���\P ���/���Y�Ll�N	
�����}7D�J��Mg�eE��W�0��^oW��'Ry��`�K9L��`�F����"kY"�A�5>�Y�o�K$P�aH�=7Г4�QOܥd�����2L/�BئP�ﭔ}�|}���]}������ڿ��� ��0+�氙2�[�a2�z����5�i|s�n�O`U�r��p0K^r�<�r���@{X��JK�D�)(�sQ�w4@��Ij�[��R�'H0g+|\+��K��[.<����*�C���K��Ʋ���*�ұ�#\������55H$W5nuv�&���K��<��@��Օ[�졸6���	�,"��M��bE:*LN8��ވ�|,�bhf�N�ic��������vk
~��	2U�j*Fp|J�	��=���UZ�k�G�ֺ��;ct��x�3��y%���pm�㤊ab���cO�N�N��������gm�ˎv��J��^�s�k�V�i��x��0]z�iO ����ofo�������~��sN.U�(?ҕe�K�`�!"�?4��_2�\~�;�S���ӚH��D�d��*��F�&�YT�|ӛ�&���m/K��¦����4)��B�;4���{��:��.�:)[#�|K�( ��ַ�E����^*�T:���w���V��w��H�r��+8 ��E���-a��m��M2���g3�ћ,����:�xKfJNa u�'^aǤ�W(Mձ`�ʀ@�7q��R�C����vD��Xr�V���<\�4'����@��-H�mO��� ��L�=���M�'9���'	W��7��j��PG�:�D�����mR�w���s0����Tl��gfиOl�E�ĕ߰�SYTv��}a���l���j{�$����o`��76��T%Df+�a��I.�񞶠Y6}���׆j@� G�Q�A+�]�m�!aM>-�G����{
��k��W�?�h�*��3vuNB��mՀ=p�I5�A��;�]�#��cz΋�_����6�����:��K��M*<e�fuFyS�r橺��X37�!%Y��#,k��|ԡ�������ݶ�'���C��
6���� �ܜ��Z��nZӝQ�l��+�@�;Nv1��Ɵ�V-Y���B�X�x�	���DW>f`%�Ѯ��,̇��ˈ��9��F��2Į���8Y�Y�1z��oj�o�g�[���(���U�)��o�cO��2%f)v�Ő.EiN�T�ߏ�R��������_�Y�?r�Mǽ�Q>����7��葺+�����t�{�t<w�\5�SYA�#�����PN��z¢����C0����������!>((~����O��tl��{�)U�aS�Yd�h$Z�%���`GC��ro%�̀,~�)�����/NC�8Q���v��a��P�(.�fՊi�
��7�'	}���M�����R��3O�rh+}T�u�d���6{�	����)�L�Ŧ[�u�j\8�Q�ò�ߘ��z@�_#�P�������_ZD��5�WN������1w�ڗ��u9h��:dNQ���%ww�f�G5�|ӌ>x'��q�+�_���Y� 5%r�t2�,����$���c�1_\@�'����'��o0*�u�l�w�e��z�W.©��1���7vjg~�C�+�]Ll_FJo;��q"���	J�F��Π%
�>�<^�+�yd�lT��ś���>zz���M�oXRj+�7�����R�����M� ށ䆛S���va�Y�
qmC�lZ�v��\�e��R|��e��糇���*�۵��*V��Eƴ*����n����_W+<�fm�rBz�x��j�j�f[�1j����D�5`6/"�|�D�U�3��pwz�I��s���Dk&o�]M1������~�J@6W���,g,A: {Q��?چ�}��y �82c��S�ZZOH!h&����\���#4�m�*�3�B���_������SfX@�#�.�18�P��x����!������ZW>����*�����۞3H�L�o&���N��s��K���P{�(k�.s4����HZ"��z��2?esjJ�<�ʗ�"Gݎ�?�(qZWvۚ"7�PP�8����&e�W�K��#P�{���9�����4�t�z�]�c��2����UW� q����K��8Ч��(��w���p(�Qdߞ�F%�����n�)��wǤh8EuY������3_9x���M�|�=FJ�r=40�=~�l�,��"��RB��a'om7r%������.�y$����5�#��l�������P��m���_�e���?Bf^�ŗ�Ck���5n0��� �%��¸��g+_�{����g�n7����]MqV����Ec�&S*��!$FΙ y��tSm�Ő�(A8Y���!!�~FHI������(�����j2/:)��
Ө��(7�d�a@��1��I�:�`@�N7Q#�ِd�탈�)U�+��Q��.�]��/�����͝ MA���ҥ�n=#3ƙ�F��W����>�}�)͹��_HS�e�q��D^�g�P�V��=��e͠��q9��i+��lH��?�>��﻾U6�gu����h~�$��\vKv��~��*m{@ty��d�@�NEP#�\�MgXR�a�t%��f�q�;j��sr�����4]Ϥ�k`|�|SKÛ>�܌@���zd.p-��F`s��N_�Z��SS����,�&�&��k�ً(���"R�\�$��x�F�+$��U���!�4y�Q�~! M��4�)���^c��C4��)�#�<kBV��L:�wv�"�$z$����].�
�ۃ���ĤvML���
��Zd%N:X�$Y/���m�|C�f�(�'F8�hZ�u����&��H�s
0���.Ζ�4���֐<����E� @�i.{��#��_9���I�����is�;���>�p�Px)�H�`�����[�k����wc�s[��[j��l��)rK��/����9#h.�8f��n_��>��Z�5�rZ���PB�y������F-��^Ih^j�CƝɸ�Sl�d+��.���/��0\�~Ε�"��N�	,�o��N�� q5��T�Q�鹋swgҋzi^�匄0�"+�e[4��ې�ң�G���������|y�C���@����Ow��\��ы�Ϳ1F.%1ll��N�k�z�0^2�,�Ol�� ��{���{��)9w%\�?�7���4!Q�F6`:X΅���&R�� �K ��b`hr�r��������a^l�*ڲD+�V�a`Y��M7r����G�P5����t[78c�5Gǘ%�<w�Z]CU�b*�%��k6�.�`��yf���x^&�>\��w��Z.���B;�7q8pg>�I�b� S�nE��|��"'ג-��С�2Yi�ί *�0q��/F2B�<�������B��7��!�Q�tCR�(ca\G�t�t�G��7т����x>�I���3��o�&�-tgf��7�h��k0�@M�$��τ��f�G�tI��Ɉ��b'� ����`~��G��~z�r(D���G��JNi@�$ޓ?��L����]vLx�aȹV��ׇ���eG�< ��)N�Dr�R`+`z�J-/�ΎO��)����/)�ݮ���N��bfgg �s���pFXNg�k< a���� �(�&��F��"C�m�Bt�~���y0��H�7�7� 
�)������?��.�����y�fսg�)s�I��w��������g�8�K"-�&B�U,����zq�c~4�r�<�=~	)2ieU[�������[�q��9\  �ՆX�ܪ������>1����
g4��Te�c����-�b(y�	�*p/G]�����e��&�{L9�-q\P�	��[�MU^�&�un3[����?��ZŴ��\��ȧԽrM�zFG�IM+ݜ'�r(�
�r S���OR���Ni1���L�+���-��`*="?��fcY3_ϲ��P�U,��Nn�7�o�#�tb�����R �iq���|������qa�.�v�q�e��v�F�qt}���F�����
�p�</����p��fJf��ó�u�*L'�:yʍ�_������]�J����c��V1����d(D�*��Q��h����C��pW��T�	����6a.�W��22�-�w1!�]%a�m��1��<2���������H�]z�����3I+lq���kEK=���p&@G���v:�@���~�H#��(v�	5��c��}��o?������epoj�%.���_7�.��7�'O^���Z"
i��D����v]�2�u��7�a�е��F��y�t���Os�Y�Jv���gYf1v�m �I9��[1V/:˥��y)~G���2���x�\�E������d�8���?�[!t䋌k�Dt�S����F�}-vV�C�cF5t�������X.s{.ǷX�̩hm]��(�8$qE	~;}U�̽]JY��%O9�K$�����Ǿ�[r�@�I�9Έ��$�~�r2��N��.A�9�
`d�d�]L�*�b,��_;�*5��P�_.�#b�be��@"h���nvr#3�����ΑZ�:�.�*Т����Y���J~E���޶ڇ{N��\>��m�S���:t��R]~ �k��&?�c��z=���1OI������ƈ�o?�{��������-aþ�	��ڟ
�W�Ǭ3�|݆���2���]���,j��b8������'�/�v������4r�I�����tb���5ɯ���:u�I���E���2� �RF��V���q�0j��3�k�_��T'W>�;��f��h;�{.(�-���4�P�(���2�ra0*C¨s~��o��K"j��yN�����
�`��@�ѐ����((�ӎY�f�y�"aw?�~�H�(#J#�򘭘�B���!U� ��D�^��$��@���_.a�y��7ܚ����2���bp��Ey����������#�n��md��3'Wg�@naQG ��8��ٸU� b�4�q��X�h\�i� �p�	5�Fnm�b����2Ƶ	��f�;��s���¿�@G��V��^KQ@Ӱ��'��(~�8����c�qCd��	�ջ?�O7!��C�+�T�s��3_^?>��D����R�g�n���k��V�"�8݇
S{�n��u�6���AH8q��N���nAp�3�恌N'F_��2'+BZ}nHKx����b(X���W�-"���3�)P��T����4�<Î����������L%x�̑�k���pq�v�x2�\7U��C̋z'��w���{]��%-.�k�Ky8��
�\�ah�W>��%������2`�k��wS�s�-粵?/��Z`�x�5�Wp��(��(xc���Nٓ*�L� }0�l�N���tUn�-�V�C���jH��Ed�,~R��>�y�1�N��^p���]a*��[�g~�XQ�|Z����1�:�0�B�g(�?���|��Ȳ-:Ҕ��w�M�a��=}U{A���!`�e�A�$'qXV�_�y�Ƙ�3�A��yW��^�SG�4��p���>�����..�<�R!��g�Z��Q�F!/���V�iT��_w��؁4��̼��n~�1Zߛh���4Z<`�s��
G_��U	I]~�?���|�_�/�倦�v��/�oF#�h%�q�,�˟!�f�C�l1���yQq|H�x�aں������b����JZ3��)c�߯�k� �%�-�Ѕ�Q<��5�w�����%E�
��'	D��Z����0=��f�s��)X<%7�h��� ?�0ca�� ZZ�`��� @�aW��+)}i�Rm������u��l:��.�W${��p��SR�'��I�-$�����q�W��-�!�^ډ��=�뤐�?�ɇ� s\�mƲN6�?���^�[�
��Y����I�_�2l��O���;����$�˯[Oz�f�p��`��WU���.�d#��0F��<lF�"��(`�Y�~�C��Q��[7K峛]�V�D�KP�Gz��$�4u�����8ߩwC��f�c����漆p�W�s@�X@v�^��ő)�y��لU�,�؟�3�svU�rD�:��蕬*sr>b�&���y��.�F
��4Cϙ\�;�^��-A-q^X��h9#���
kM���x��$1�7���7��Z��{��;Qu{��f��ϴ�q�ά����.�X.��ȇ^r�s���^u������&q�jy?k��ykA(ؑ������I��cGC5 M�z�z�<��b)=�1�Q��-����LtڧO�8�0WA��)4��/wA���k���7�~	4$���Ʀp��t��~���Ye�Y)}
\Q���n�a����;��3�U_�P�����7�CGOH��� �02��Am9��d׈	�d�45�&����6�ٸ`�E�UI�����V9ꔮ}a�S���"�C&ٻ�ǈ
NW�x��K�&L�{�!H%�I�E��4�l'��aȧ���XՉv=LaÄ���D��S6��IP!��ei艶@�c=�L#3��VC(x��
���	���%�"��{Zt�H�{�.��CX�o��D�h�k8�]������1B<s")�)�Ϻ����W^���i��C�2�<��ku�N=�����*��Y�Õ�5M�V C�k�'D��Z��(�9k���[��K�����X��ġvMZ��{%�(P�@*�#�>���$ݸ���pr������d���/`����6+�P��+��ܯx�a9t�����!Y�����F�^�[F
LO뉟��	g>р\\�������Ĉ��K��Kx��޷vE��Y��qb��������>�	\�)�Mt5Z_w�V������G��L�^�p��t��N��w$86�s���t����Ϫ�8cN
�4t]<���O�`_�����)R?N���Nt��ew����p꫚F�A�YlvrS����,Ѓ.�'Z�� �Lw\��.��ˬ��K۰+wF���4P=���ҏRH���*���TMpvZD�I-���2��#�{3d�:����|�Vo�I��Y��w���e
~�u�;�a��NJZܦkh�"�(,K*�ޔ~G:$5R<�4���p������nD�����ۥ���vE� )�j��	u���������}�����3:~�%1���rc�`s`����L�-�-y��j/~���s�QS�N���9�٬�ʪ�f�Q|
�$���U���vb�G���0�Pd��ig_y_�n���\P��j�Y��!EBČڢ�P��X���������И,D�h��PV�ײ^��dǟ��v{h�Fx����ZT��r�NK�
��r�5�x�pq��C����D�z育>�(;p�b�;6f��u����ƺ6 6$8�J�l����j(;�)�A��O}������"�s��HK㖮�h�A��ĸ�����vVG'��.%�-N�tHþ�N�%%ęu���<U�}��Ċ���s=D�^o��VQr�"Ò� ��φ��W���ő��躒��|�mx�C�܂� ���t�>����e���"1UY�1�G����&�b��*�Qx�O�	/Ku'MJY.n�?gFތBR@��.䥐�m���$ҕ��~O0����V��}+� S���
�E�J3W@��zhPJ;�Fϥ��� Q�d�c�,�B��%{]l����U����D5��Fg�L8��n�1FD�5\�,�w�,jk�Ρ�i�o\�{mD�>]�%��"��2 O/d䝹(�x�U�r���|��ь`P�������[�j�<VBD`"�?��a��Z��5D�^�r�os}��5�����k;+i�U�;q�<���sn�������oԨ)v+�k1�J��L��G�|��Og��jԙ��֠ݺVeG��Q����P��3Z<ǰҿ�󯳺Gr#�mX���0h	��4�A��ޒNYB@0,9Ѕ݆�:��oo�����A�m�k��|#o��m�spU1U������SAs���D�D����"!��լ��E��(O�0��fYS�%H�� >::�����_dX�m\�nFC�5X��ޭ
��'ցC(�h�7�	\kE�8�-���B��{P�W!� �m��a=�X�'�0��D��=A�4�RfBr��U0���ӳr,x��&�mH/��5��#�꼤;��G�*��~�����+���"��l���$����Nn�������zGS��M���s��� ���g@bV�<,a��?G��ė�@9�`����!8�n��!uJ�ǿ\R�b@�(�lk#H��^��fL�V��k�7��`+���(�0����ɒ��`d��%�s�pl���8G��F��B-E0gH�XM�����Yl�C�� �b��+��ܳ^%���ju�Z�����~�l=4��^�H���lp2^�-H��:`�yw�e\8>zDp�A����1�H�������˭T�V@��.�(9*%-����՞fI�2��*�~������_6M?V>{RUq�p����ŭ�+i�D3S��fe`��3s���mx��H���@�����&K���}�r�	��ڶ7�����/��_W�ދ&ߘ�߶��P�	��{x��*�*�bf76��@��-�"��n�x$H�+���j����CX`���b���K|�z�Q.̼�A&.�u���D�^���wYN >^P�^���$mL�kZ���h�4�|9+���=��>z�̄�Y�M,�����+t���F+!; U�?����.�I�:<�U�\����	,����[��1�}O�tK�i���*���:6Pfl�L}��Gk�c�a��b8�1��C��e[�j[�ar&V��`^>�8�+�.�[Ʃ�ֈ�<Q~Ea��F:wP�sh��-�� ̑n�߷ч��#�%�pu���ACa' S~�`]������}�E� 6�A!N��U����qi�ն{b&�NUs�U���{N��.S���G/K��gбlr{d<�[%�@}��[&@a�Υ83IP+Uz\��?-7U�oE���ȒFO�1Ģ y��$�X��B���, 	���/���~kV��N��>��D��v�L�\R2�7~+]MY��wh���Ώ �f8-㭩=N{����}I�Fe�B0��s��A���I.��RW1��ȯr3�4�L��D���.-��o�ip�WmR��R8�
�n
�h���fZ��{g��ݢ��1@�����+�=�U6�Y�Y���0I5�MV���УQ��\1�P� ��1tC"ʌVLy���-�.t>�(��m����Kng5�)�p��.Ol�QT�/l��ρ?�"P'u��z/唖_C�0{D(|cQ��Y��e/��Mk?Z�~�0*AXgm&�#%uZTx�>?��A��_,$�~W��$*�D<�N�P� ����&�ۓbH.a��fw3�ƃ��� �>�4��eZE���2�a�b����ΒcS��ݦG����-#�W�^&"��u�h븫��a�w���"�k�V�%�i���_�Ȝ�+E�|%t���:�!BB�l~7)V�<�?� �'�\�	o	O����G�"\O�V_P��(9m�`�5��M/lա�-�xWL���3�7x���Ծ��aRf]��o�Cd��{.�f`Ƃ����H(�A����~G8��O�/��G��Vq1��=X0"?�Q^/��K�7���fqJ���~8�\� n" 9UW!X��a$�$P��Yp�`�#��;G$�?��8E����Ɏ����i��L���Z����h��IL�OT��[W�2����iTN�V
-Z[��X�;Ѭ 	�ţP�;"_����םeI�6tہ� ��ڞ�� ���W�����A����[*i���4G����ף�`d�U��&(��R������+�Ѕ�`--����H��/45��|�77���1'��m� �Kuy���k{U�+_��&=Z`��X�1G��S�v�I�Q��O�FV�T�ݙ~\(����Hñ��� ��g��}� �l��ʏ�1���GO�Vkp�w�T�XJ�������Vj���޿��'�^�NΓO:���%�oeWFb}�՞7����ټ���})�WN�Է��а|w:��ʋ�����ɢ~��?�{c5���H�MwF"�%��6�ֆx"u=�n����s�Mio="���b�ق�z�.�Ĺ����G������ag��{Dw����i4�rn�� ��E�#��%\B��NB�H��Oz�CVH?�%�q7fԖLY`������k�͡PmH?�Zr�%F��fP��pD�l��e���n'ڡ�\ίW��3�l��A[�lЙ���^-9�n���]N����%�h�h��V�t��-�~����4��{�}���/�
dM�㨜�e[�[s+�M�F�e����z;(�I*`"����-�	���k��a� <'M]j(��d]��Q1��=�G�W���VH'�!J8 >��=x�ܫsQ�'��k�m9�tđ�_(��\����֢�X*(0�w$���?���/����q�l�<�pT���"&n1����G�^0� `�T���L[�׏�C~�:���KM1�?mی �����g�1��N����|x�������a�����oF��$�4g���)�j�6���م���r�r���[��p(}�n�+�F*��o�����V�K���?J/�� z��^ Θj��}��bg����ߜ��;��i����q9g͉�*t"<���U"��ierǮ�ow��I(+�!�
��(B�0����𶄁 ��zՈE�\MQ �	7pl�؄�-�%������"j�S�w�u�8��c<,\R�����+����V2�,�.���I	������D�Ю�aMJϻ�!��l��Ļ2_��RKoyN%lD��Y�~	���bp'�!X5��cϨ7ڻX%��xOj�e.�j�������e�C�@q�	Sʍ�f��4Q�����x�n��x��jgTI�X�:Q뺌�G�dfAjGI���7�0N��Nʴ�]����޿|��[;�@r���"���)�[���`����=�n-���¤��x�X��i� ������f�����E��z.S?��{?3�}�W����_�Zo8�'��S&{��������ۈ��5�`� \����l�_�������w��(H2}T�/��B�/OK��C�d�k�2Ru,7����'v�vA�}�X��k���prr� � ��e�2m��&�Seޢ���lc���-��
W#�Vb���5p{f9�\��CIiO��x������+�m��Qt��6Z�e%ĐA�%8�N���v�����J�$�i�łq �ۑp�㜼e.�s5��f"�>"C_�6����(��*%Ɓen�S�@L?�?�Ӹ�M���[[x���:�ٵ4��]�ɒ�����߰_V�KGʿV��&�$~�YN�����]��0U)	 9�5+�&�k�TQ���&5�p�9�Y��;����͈�-�.jn�� �}=
I�y����2D�=8�����5�e7PCs,t{�n��j����ȧ��#�^[l�mFŧ��j��~G�0c��/�s�V�g9���1JdO�)�u�t���e-)��ۨy�\m}�|�F�>\c�9��ƅ���Ʒmӂ��~_Kώ7���sN�֤�K��'�'�E���#�fgT�L��ိ��d�&�Dxރ! ���SǬ�̋O	^.
�S�����.���<۵�	p���[�)�mҥ&��0� ;�j#����[=NDp):���3|5�Q
/Mi���xj�"�s{�M5�,Np,�Os��5���Ωc�И@�¦�5�/�KN�/BS5(���MX�!�C'X�/����Y�4��;�N������RG�b>�D���F��;�x����#xp�9�0�r���}��� 7u��o��>�#���ol?}*����b��2|Q,���>�t��/�+(�;��P�ѿo����n G�>ބ�"��Has7t�+G2KCcm�����7���A\����qz���]�nM��kвVϥr�P�8�����7˒^I��uk(A�6m	la�F�x�+���ǌn�;w��2I�U��P�|
.H�_�3�p0%����_#)��I*^Ռ|�BØjJ�N�#d��"�/GO��%����Unr�{��|��f}wb�a��j�q�(�G'�ߡϧ��LF$�W�죥K�N[.�����@�\zl���z���)���� ��)���5˥�nu���a���|NQ�[#�d��;�2��m��gn�����3AlQ\d����f��ݳ���I����y��`Sk8v"�0ͨ����lR	�F���Y��Zt�FX ^��3n��Ģi�Bh�sF�aV��i�q�N�ݢ��u/����Av���EV7'�Lb���}�@��;?�g-Z�R�C"���
N�K �
ͽ�/�)��R�
��H��.~�Y��:��JF�Y*Y���%P��-�h[����mlo��r[�})n��������cؘY�5�r����~���V����h~�b��xE5Uc��'p��kx	f�� ���C �9_���Ɨ����u��r��ir�[�J�3~��)������gN�ԮBtݿ7P���7�;���Dm�N-l������I��/Ţ�SFJ��L;|"�1�$%YX��+h�CiC�:3͐.���9EiI�3�k���Q׎����������":�b��,}�����l[k�1���i챭w�D�տ�>4چ	
�J#�TMv&R����Gc�!P�����{�;Q ��X��gW������<@8Jб�AۭA�]����R�J@�Z'�x��8Ǧ�f���r���h1��VU��T*W�KB3V�<C�U�9V@kg���P�
��nZ?��E�D[�uK.�1K�LbH����d�6L@_q�9������FB7�A~��c��@�%gQ�x[Z���PZ��J�Z�Z��8�7�S����	w98sJ�Y&q{�1�~Kdk�`m���\wt��� �4��H-1e�Wz
��Oo�۶���Ӫ-��04��Q(q=i
7��y!��,�����}���r]�����lS��7�Ԙ�vH�c��'��(���t�&Pk��+�Fu����"~�as�ÙT8��b�*�?MV��F,�'�q�Q�|�Fl�������j�>�=8�؍�]�z]��z�DÚ>oeP%�U�m5��:C��<2�N�t���o��pU��@:�NL��fw�G9��;1M���s� �̀���&���I�����i�p�J� ���]<?����� \-�9K��g�oy}`3ZAj�z繦��V�¡6R��T}]�)_�kY�� {��.y�t���37�:� jmr�nw@�	���Ǡ�ӧ�"��z����p���O�'Ͳ�m*H��T�J�+�E��=�V3�m��a]0:�Q~a�8�:�q�%ww,ٶ��.G���j�5J��Mѱ�@V>�F7��_r%�Q.�V�vTs��:�N��w��cuP�Q�þ���;��$Bc�̈́�w�W]�ؘ��|+Xͽ���C7פAL�� ���gW��°�f��:7�,ԛ�yy��N����4n�^\ΞCs��V�g���0�v21����[x֬�:RM P��ԩ�Oz������͌���m��X���R���.��F�$w�;�?U#V���T��Ԏ-'*`�� n|3h{p�l�]���g�A��d�(��b�Y���ķ9>$b�������o�|V6.��$,����
��j{w46��T5-�����
,:瞎��"�W�+�o�S}x�$,��'N��������E�s����r�?ꊥ�pKE�4M���x6����Q�H�b<IB�Uq�͆Q1��-�oqߘ�e���0?}"w�/���]۵=wnM��q�ؑ��	xV#p)e���W�C޷Qj�U��� �-�����_�����J��ޔ��&����lTա�p��E�A���e{n�gP���R}��;@����Y��<���	Q�z�:56�b���}��W��:q����3��T� ;4`'���0#�f,Ԍel��s�<���\J��ͷ�U'lgi����ȗr�o�0LBW`#�"S܎�xΠU�&PۓI��tT-�U���yf�9���xx�?�B&�%�)y9
"Q��}���5x�fr��e�T��Q�TE1�H8NY�v�����p�k1�����b����#��h&
27�ܧ��$	ڻ5TI�ɵ�h�R���oϮpgg��ǍS�nn���*��Oj&�v4�{7��������N�p���(��̕���@t��g[|#���@�4G����WXP�f9v/�}����EDfя��-�0BF�m��GR3_�OohI-��m�ux^�p2`f��-�S&#�Ny��k�(���q��P��u�� e+QY��x�i�H\�V��&�[�T,Mk%�u�{H:��~�R]M��6Ӯy�c�?���4Γ%ߙ�z�k�D�N;��𦪡��+�Z�d�fpg����%��O��~p�AZ��ψ����@�����ʮMʻk�'wT8��_Y�l?�Rn$O��/�=����8��p�a(=S�ͅ_T��Pr�8����}�J�,�1���&����SN���B�K�oPc�@R-��Ⱥ���Un�0
G�bP��A/�쁠w�B@C�)Q�Pb��F�849��/Ji���[�,��m<d"�$CS�	��
UN40A�j{��7�tZ�y�������#�`5�*�����y�'2�����U[����#9v4�����M���I��6�<����KsQ�qV֚H��L2�"�0���VӸ�p� ��dn��%pSo�t��r��ڋyԣ����|쎀�۷���c%�!2�ƁJF1dZ]��cW�o�}���k�!
���J��܌�����s����o.��+ �˗6�P�J��}Ǝ)�B��@S�Z}���-���38s���Ug�@�(�,��&���o+��e�a�u?Z������NW"�H�3m�Z�cT]j���l�ޥ�-��z�'s���g��-�P&/7��A��ߣ��Hd�AQ��tS��R�ΐ��" .�J!�_�k��pS�	��1��	d��ާeu82w[�)�╟7���m`U��+�#NUp^��L�I�""W{�v�q�+�?�9.&өJ�'��wW����+@z��QW�N�V[Jz�*s�FKAx^��$��ӳ��7�Ϟ�1އ`��9CfJ�ϕ���͐���u�Ʃ�lTf!r��.ȏM�@/ܐQ��V���;W��Y�`-Q-�;i�reԤ+�VZ9 �}����c�k��tc}6���\�W6��bQ�#4��ؔ_]3�{v��fpY�o�$t�	�"����41��������
�a�^��~��Ɠ+{Mȣ}�G���v�X�l
/}z����oN����'/(�Xk!��e���E����ߩT�߲f��;�b;�f�#
�2�_�_�-?Ͳ��X�;�b�>rl�6�t��n�W��<�d�j�1�dђq��4����"݈$N3��<eT�ɤ��R��P��--NK]:���G��ր]��WF���M�P+�ٹ_J&"`�#�>�L��kۋ������`I�s$Q�C.��]5��h}����{�(���?
�V�A�����
Q�h��큡sA�"X�g,q����TX*~��x,̕��)&�lvZ7�l��Iܛ�U�F	�S^�Y�EP��GZ�'�;>�F�d TQ{�GUš�0D�����Ģ�d0W9�4`�EV=�F��G�V�NQ�r�zq�	�m��P������:i!�hj�׬ǞڰP�Ku7a�w��5܀�2�H�^�y���G}A�]����Sr�-^f�溠i�o<d���hjm���pV��<��}�v�l��~����k�GZ<���R���������J_���|����Ս�4���d�%����Z0��Gx.�8_b���v݀��l�XSX�b �6`~t��_���������ύ��w�Mb������y#��3�o�����4�0"���J�����랋��A����+�y�֘J��s�ϴ3]`��/�/���&C�6]��C�)=�q�Ҟ�k1��GX�ӑw.� C/j o9���D1��Y�.��4�ld����}`9m����Z����Rh�r������F�z�p�|sIk�a��h������6�U�>\�*g����k?	�`�?��s	���q��G�8���������7Ibفy�� ��	1b�FXDq�	�?���=��;Z�������'�s�Y\���}>)�u��l$i�v�:�MYj�no���9S\���hrE�r:]Y�֖�i��jBV�E`:�$�#���d}|&T�1|��A�����a*�4�6o��sQ�Gm�0�Sn����#�׊b�\)q#G�%�?9��}����ݿ����.N�Uoue��3�~���6%Y��%�c��}Jͳ;�bZ�o[�[8�4^�X�t�K-y#Z�AZa�v�kmI�����zJ��ǌ�z]&���Jo��j�B�94p턓��F�*B���J��`&C**U��������m��ޖ�^�Z��DUP6m�����@b�c�A�ή�r��O@�\�k��뀪z7gW�w�^�* |p��H�'?��Edr�,n�ֈ"x�r��~s�s�b��$��
 ��zR�A��������Jgr��)�4K�ga�Ԅ�j�\Y�Yƺ��3Z�PT{�����ZM���h0z�yX��ٞ��Q�T������XP��|�1�3���r��z�P羍irU�5�eYkׁ�%]�qu�W_o�Bt&-�c�Qk�mk�I�ؼ��Ky2?�[X��z���գs"B^D�o�(8��ԣZȨ�\-5��.u�6X��W�E!`t��l�m�[��ķ�G�%Ԍ�E���v`)@��n�s��u	 ��.#�u>�m8̢�3���;�c$�4�@?�S��k�j�a����4��u��@��Q��o�!qQ��F�v��k~	���/5;j�j9�G{���fCw�nN�s���)Qh��.�QF_L��S��	��R��f~��5�Y��6�З��;k���C�wK�S�� �a@�1�S��:\G��T��TWr��c+e;�?�0���M<�^:�4�"&�q�S�8sv�U�w���sR$�i><4�k�9��Kج�e:MP�{�z*��J~�͙w�ηJ���gJo~�����k+n>(��� �#r|��p�$k�2-Z���Zz������c�����q��r>[���שr0N��G���FI3�����5�d�ΜAO���*<�+�������p� ,9/������'L36K"�TZ3~v�[hM�FL_U�=�����-����
�`q�����Lh5�[�-K��:i�(�օMM��)Y���G�O��,"� �o(�By��*Y�.bP�z��R���ԭ�Tk�AV7�T7�\}���KIˁ����W�V�i�z��+פ߱�.[����� `�G0�I�V.�D��e�V�����Z:�G�/BuؐŠ8��5z�1\,�C�p���t.cI&����)5�������t�Mxr- �����|еC�.1���2X�L���H��A{B��cEw���\�ic>�jN��V�"`����?N�2�TDZ��~߈߆[mǹ��|Kz2�+��7���O*x+��a��e����"�q��G���ᜃ��uv���~'�#���(�4�Rzʿo���Ύ��R�^�l`��FW̯v"~@�ڿ��̧D���B��
gu�c�Ъ.Gk�Ӑ �s��J,�M��_Y����&5'��0���ɞ��T��_���&ӈ&�I�~;����6�叒4��*\n�W�������� ǘ���N��d5�ؓ�h�y'��^'Ǫ@�8�Śݿ��uQ��R+}�o50j�R��Tg�1��.h�A�3���d��B��}�As.&%(9���.r�1����*�X��8a�]���IM�m��É�3@��y4���+P�
��w���r�`��e�q9j����D�A0!��J��R����I�W���A@�g�
^�
��!������n��<ZN��?��Og�ǀ@w5�����	���� 9��'�`�1땽�\y��e����wn3��ǉ�X����;�� ���O[�i|Nn���N^���ঊ��Z?d.t��*l�mߤ�W�S�oE���C*���F
L���	e�BF1�����S��/z������!RAKa٨�jJm�H�K?��9��|fV<Z/�*�#6?����ᓽ������L�Fu���^IZO����
J[�k�]G�����WW�A�����t�$�q�4�d<��:p1�������*�f M?w^X�E���� �X��W0��{�B�7G��͍|��'	��ƛ�c)ۼ�m�Z�k�i���
IU�ؑԞ���mC�ں?:�/j���)	w�zE�&����%���.²j��*B�h[���6N00����*\-�|����x^�
l����;���ޭ�0Du,�=���9�~��'T0���Oe�N����4�κ�p�[;Xw^�Ҕ%�bD�������K4�5"�"FVQ���ڋef%[�����~�*�9>4|�L�}d4ow^�v�K�[*����q��A*=7�m��f���^���ٛT���؝��v����]�65�P�#��K"X���;ү�w���p���%ѐ:3�<�Z��)m��Nꐍf��tS�J ��|l�mf�x)�*.ӹ:�KSJs��8�?�����h��z�,�k��u,���c�^�@�^��� �a4��c)9�}.s�9Ŋ���n��@9�i �n�q�<��6�����'΄�p%��*�мV�����+�w�t�����"����Feb��� ��Z�OR�]�1�%�z,pP��Ҋ9���YC��	:� �1�O,�sҁ�$�~���]p��o1C�J��"�LW�_�[�����ﾞ�:�|	�)��;�i��r�M+���~2��|e�k�J{�����3ָL�IݨI���f �@#f��I���W��
`��,�INȟ�b�%�=,���~�Z fO��zy��l;Atq�����mɁR��7�cD[Վ5�Cm ��Tq�)�I֝��O��K�p�(�v@�Tg���/FK*�8L�Xֹ�����[I���l�m�'�ԧn��SxbYυ�u�i�r�h0�[������ bU�_���6���D�ؕk@ݥ-M��	��>����˚�'���V{�"�y�t���ۣNx0���w�(92��G����E���̪���ٳf�2��T��_�p,A������ܘ=���eښ�|�Ws-]���Fly�\CW�W=�h��WWkB8F���!�8��E�i��8G��&P�C�qC�(f��/d�#��(���I�U�H��1�u�Uޯ�Z����,q.؆�w��X��e��+�++�A\O@6�`b��0+ͳ	L�����I2��nUDosF 9e#-��;1=
f���ν+��K�E1�3`oѪ�}9���`�WSar6�^��"�ߴ�m�g@���M����X#�0@G���������x����>l�>�Mu��]l�����f,��B@վ�)��m����0�kH��.Ƿw�!g\�=��b�r��!�p���2IcZ�a	F��l_��o��rV���tPy�ͳ����s�@�Y����H,���U"�( �Gަ���cFt��{4\*���w���Da��̸H
U{RS�����o�bmؽuz�@���u�u�z>!�=\�����!�e����Z����n-�4�"svH����\.��[��y������ltKm}yD�̍�PG�~aM�Zi��*�qF��^ ]цlSw�B#,�RJ����+Lޤe<�\w�$Wʀk��o�+�88������h�U��o�c�����!��4�4����5���:�<��y���O=5APZ��3A^��+�}��,��>���J���jFSja�M�ų���;�ؽ7�$j.��-��r�%\U��ؐ����� d�I���`oiҭ*�P��y��|gi�ā{#D�,��U[ί�h��k���ݒ@�����f�-�}Y�o�0zُ,�AXF#��%�����C��ܧ��V�?/LX��u���Xf�JI���x�B��4앍�Gԗ��6�l*�]�����<�Zrf������-��	F"�Ţ7��2���H�K�~9�;��6��$1����5�Go�#��p&�f�ObvMV5������i��sp����VN^%U+p �a5���<��>�`�ə99�)C�!�\Xb������;2���u���LH��b��t��H�����E��wzu$�K�}�W ��6��d�+����V�>`���i+P(����ot��9�}y7���e0-��쒒�'��U�SE��&p8������˫���\�o�B�ۈ��c����� ��.:����E�V1���VQg�M�0�k�Q�6���G���\b7�WQGQ3��_Gډv�T�F��FbT���oϑaPHP6�L��N��Rd��ف��mB�i��4؞�����0z@�%|sD��#3P��&<!�on�{W+����P���>���KJv9��8m�я;�K�RE��N��Ap�B��L&��r�ZF���tL%�C\�A�iЏ2k 7[c��*m�%_��]Ih��B2GR�H��ߖ�djdN�,K�O���w^��R3��5��j���7�������ٻ)�+w��Kb��H"?Ӱ�N�z�Ҹ��u�.�?prĆk4 ��'�)B���Oob����^8����1��B�����Yp�HX
aG��+��\��9�{��͜2;��[d�����9��[��>κ���Ѷc���Ǻ��˾\^9�ﲐ��2�(���y����Q��H�`�Ĉ��r+˕=Zl�aݧ�e�uγ��|k\6
�Rl�(�ϓ�#��О�z����0���9g�x�����@��jƫ�������� ����$����dǁdhZDn0��*�d��e�OZه)�s�.���}z��e������d��'Ųe�n�Uc�A����p� ��[EJt����< ;��\x2�!;�� �VZ��9�`�y�wm�����M1�����M�d���حrE�(��l�e��6�J��ts�e�4�	%�.���VS�A�&S��Ύ��O鵫�i(��9���k�7�4�����F���3�G;�����ᄟ�t�ja��6�އ���F��T�a��:�Bh:�LK�{���~f���V�"J��s.lf.w��@�`��6ܕJ��J5Ժ�)�����ܷj��`evZ�U xeLM�d(�G�G9g���&���҂�Y(��lo;E���}m�P�~�'�0�ug4���ۻ˅����90��}]�m�"og���\X~ 3�����b2�~����-�sG��յ-��;�{��^u.\EP"���O�6��:L`���g������W�F<�d�a�96*#��w���MFw�A�ٽ;��r0}%��lx��o���N)�0e퇪rǷ*I9�G|��GM��'}������`��k]�M�K/;*͞�D����,�Rb^zS F}$�]�z"2uc�K��t�D�iI
�zo���ؖ�o��{������猑/��Y�4�2�M�$��3�q8�=.z�w7Ln�JJtNr�x�8/��hB���.�'?F�i�4DApH�3^�$7A�	��l�'�|���'��8͟�9�����BU3w2��<� ?g�ٽ(d�q~WQC�kޭc��eZ>��O�"��Cd����"�ܝ^�=��b}�xP���a�y�ЇL}@9܁���Y�>B��6;��Kq��"#��]9��ɕ��ը�.���0~y��G�O}�ٔ��%35)�{��n�x$s%47�tF@|�9��yp\�#�_ր�m��R�к!Dduj"�=���FH�>Z��-g�4A�r�uVM`(x9P!��g�!��O���dY�q$��RI;�|�
��֞�G�M�m]��J��zkI��GV~5q�X5A��r,G�X*�疞̣��	B«�
D�{��� 0.������
�fS���cȺ�Y_V�^q���Cų����q��A�'z%3B3�_���e������%��.���|���|���?x��)دՊ�j�+��ZO�Ҹ�S�E)��B�s��N�0�Jel6�2M��O�:�I ��(z\տP��G<"���t58������-�Rq����
`�$�}:t�{�4�Us���Wy��qo�0T1���^S����B?�,�5��`�����"D�2ߨk�1y���ka</+}uk�c�fO^���a���[��D�/bp�TN��L7WqP�)Wh�]��:����q3�RP���D4�2�y�i���Gv��*�����myS�sK��;�$��_���Ӭ���A�*W!'�]�lu�n�������[��6j�Y���:r�axnE���Kr�$���턟�@�m[��Nw�M���=C��]{�ȃ�K�=�V3���K^�q�1 �k�n�7���H�~��@'̜m|e����b��J��4��&�y��`��q���gקg+vU߅�އ�ynoc
fz#��(v�^�*6��"#[��Tl5j]o�?��k.�Y=����k�i���~��@��"�zZ�1ݗ%9d"��=`�{պ�3��O��y��7���?*" �Zr�H�(V�Gϲ�VX�Έg|�^��mh��Ў�3b}9���l�����e�V;������0ḯZf�Nm�t���]�
Qo�W85Jǹi����0�
x�b�5���M9Jf���	�.���\�����Nj��X��?���"u���O&���S��{��V�(ju�����E�e�8tC �xXq���(7���ZOj!W3S�����9��a�pO�T񛄆6l�S-��'i)�}%��_@�(xG}-jZ�g1��:s��l�P�T P�7��tc?6 �~��#[��c��T