��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�
y>F�Gϋ� 
��*�4QK(��7$[M3�E �N����,/mY���n~���M�ȸ��� �i�ӗ�3h�`D#����V'���F8����i(bʭgU��1�".���x�Dc��*bn��Ջʖ��љ��@Iz�eQ.��uS�<|�������y��狍9}�r�6c�(�D���gG�����+}�Q
�o(p��#n���)�lgK,��\.�<�����	 ݛ^�A%�%�w<^��Dc$��k��?��h�WN"�&����O����.����¾X�Ϋ����ul�o,v�����H�T���ů���k��\ie�a���p�ƴ?&Ni~R�J;�/���]�ڡ2x0f��T�aS�s�0�a���1�[�tM����f��TaH^���7�8�Fq��w�R��2�Q96L#�#���쁎��3�X8�/Rk�Y�J}��\�~��C2d-Na�Q������e+�-��^����8cgaǣj��4-��U��zu���YO�v�}�NAP���_���������GNշ�9IX��?<cY-%�k��ar[�p�
����	ݜ����&"���P�o%rh�Z��*�")�N��B�t��Q��`j`�٧�����8S�ňJo��!��� b~�{EԭR�A�y�!DN�v����h�B�`<�� �#�6��6·�t�?�~�}��>x�u�L8��3.�:1i�z�q�H��8s�L�+;�~���J ��;'���䘫ݳ��@f~�@��>S������
Csp/B�= 5��y�p��N7�?sp��;1ˁ�Q� Q��AoE�\z���gg�Z/�eD�^ul�������-Xwv8,�lQ~�QX�������=N���	��M�_���n-��fPB{u�g̡�C���a��j�TT09>�7��Hz�c�k�(�E�"�0�lw�ͮ�g�r��)ܦ?th�SӁX/�m3��
�W���1�7�`9�?�F�Q庤HXOB�.r�2Yh�O�Ŏ�������Mi��| �5p��w��zwA\��RI??~�u��S����`�L�T]�6���[����ǳ�kՍ6����C�N��;�W�OE��z��yK���~9�����@5�>|JN�%g�,1@�-�U�즞䬶<��h�v���>l{Ėk�C�{� h�2#�,9�T|��(���܏'=��D�Yw�;�������ҕ�CG�j�yrg���p_ �g�)��w���Z�-�$$W���2���HӨKn�x��0k�ZU��?�]�"�:���j���-�9���q����*��5�����x�L�����OT�0�K� &��v-��ӆ��eޠL���8A{w��*������>qɘd#t��j�<�S1�!�é�~]yB���� �b*q���W�0#^��V����-,����FѸO!R>U���e� �����)�Ǝ4��R�c!�H@��� ���E4''y%9���QW��> �tfU(H�rᅵ����R�o�Ѓ� |�@#�x�Ρ2�!u�W4��^����.�i	�19s+�,���Q������h2>E!���4dG!O��[u�L�$`����U�w]�����t47X�⪍s��`��Nٝ\-��7�E2��0�<�G���8��un���u_\QZ���k�J�F�y-
�1���̃��3�XG�C��/r@Rw��p�2����*L��'��J7��Ӄ��x�*Q�|�FX�M/��OU�2�Dy�[3`�}G�T#F�����&/у��W0)g|��+m;ֆh��7�x=�A�۲^�6�6�4�蚆����p9a0S�2&��l���d�+`�,�Ƒzo$�ՠ7�m��eT�Rl�DO�9�y�6�W��`,Z�z
:ͮ`߭��$`7e�Fuĝ����$���	�.G@��Տ)�U<�w�+ӝ�~��`�v}r�����j����Q|�\������ԁ���[��ի�=���rO�֟fP!����]�ԭq��4ۖR9�W�}��?��CK��,f>
j�O"�$d͑:�@9%��m"W���Q:^��	\���>sUOn��,�1uV�{�\��4,���ch�����ƞX-*D��`K�}9O4��J��@��q`��I��i3Bo{C������[����n;���y��[���J��7|��=�j���0�yN)2I7�Y�ݦ��A'�S>c�aj�z��tNK޹�%u(`C��{�̑Q��w��V��A�?����Ȼ�q�UT#��2<xx�z�JxY�t�	=tɹX�l�a�<�&�Z����Csr������r�K��mZ��x��B%�/�t�$�aƜ����K��i�?�H����nz���(�7�&���6�@)���r��؄uL�st"'O�bi8=k�E��r9�6ޓ������J����-������BD7��5+X)"��fI��$���(D˕��+ �g?�!�[�H��d�8��#%�iD�W��)����7�Ҹ�Q�k�"{U3���F:��Rɩ�/��W<'M��c�{Eǉ`\<���T] a]�m�+!���D�]���6Y�NmEU9AA���-���N½T�1�G�f�w�h�db)|f���^�]���3�����zf�b?�[wW*8�Lⰺxt,S��
҅�"���T
�'������n��-�F��ՄOkk��V.`�K�Qɢ�|���Au�d����;�SB��f�w&/�<&�4ؐ�E��ϫOE�vv6PW	IH(S&_�ɪ/c���,�5y��C���ۗ��D���&P��H��$v���!�z������^����,^�x����Y��T6��l9m(��wg�N��S���i�6��EU��[T��a��������|�����*��Ƴ�d�wzo��В�3!��	q8S�{Z��&�&B�H�.>>8DIm��3.��+��u��R.�5b��(}@����}�(98z��3�I��D�����LH9!���(d�<�	�z�{2+��o�ހ��
]����c�6�X�,�,3��"=�@�S2�i�L}_{���h7����#��|a��7���5<hi%��i= !˷��ܮ�1sܘ)h�U ]���π��إɢTYд��wN��W��ME��uM>�r�&��2�8nH(�n`����� �;��t��k��?����Ӷ���w�ܼӨ�"�����v�oaT�#��q4����{l^�Af����:�p�&�l�a�����,-g�+�[)��R�@!;@��!�k�St6�#��k#3e=�����y��4������l5s�q���$z����{�=:|���5�vN�D��P�����yO�S=�����x0������Ճ�j�*ޏV�:�H"@��U67_D`�Z=�*N������`~�j�7*pd��xu�|u��W��b���&B����Cr8�4�p./U���S���������14kJ=�x֕�?��ۇ�������q/5�K�zı ����l�bS#�ip��T���eQ�6��L��$��o���Kx.�@OUs���J�����FBJR����E��V���H��ㅗ8�r�: S0�e���;����
�W9_��Z6W�K"y��ذ���<PQʘg�����}�.�]觮z�l�#�#��ӉM1�H����_Q���Wul1e�O��5� y,���|�Ϥ��Q�+t�����h2�ܱN)�-n���2K?��I@�MӋe^4���K-��ʠՇ���{�Y��1x��@��*�N�+�P^�y�����Wh�&
�>;w'�aT�g��j�TDQ�����fo�����+_�h�����F���̸=�$��=�ܜ��D�22�:��'���"���F�8�FRp�|�7�boD���eN~�8�8��Z��/-����6�M)PXCb��,��v�p�0Mz�)�TÈ�)8��E��q/k�� �4؏�O���[�G�g��4 �JJ�v岺�NX� p ��=G��w���p���
4g� ��[`hG7d�݂�ގ���Jl��;F�t"I�(��veD[��������Q�x����b�T�4\*��XB�A��ܯX��9oԦâ1�]A�34b]�>9/��nwL0���u.֚`�V��(T�j�Y�ڦ�d��U:�JZ�ز��s��Q�$��9hUc�ӂc��"��Yͱ���8�BıG�Y`��Zғ��v7�\F��Zr� �?�#���m�� ��c�����·)��'/�"�c1h�j/�J�,O�O~ �Y>�$�Q��h	���A���JtJW�H�R�j6c�tJS�����U��j�@_x�IS�C8�+��@P���*��/��Ա�i6���B
v�����pGde��n��k��T�:���x!�M@a)@�\�e�.k�J5���EdT�7��zw  |��� v�1�[p�.��!a�k\��ܣS���ʶoK�zZt�h�\�	nS�%#��=���4�sBD�>fs��8g��4�T�0�'����`r�aT3(��J��-�	svǼb��F��%�]�o���H��Bν6v+[� �`K�L^$Ý�;d�9Kl0$)���^����aוpw�@E���4z�y�ݚ\�Ep:7@a�B�����'�ϒ�M�Z���S��n[�3_�dw�"0�T�q����D��H2?�T��r\In��-_�y��`��̟}|��qJuוp�4�$��yR9KRX>.�R��ޯ#(p��@~W�At�*�h��F��ɂu_��$�s��C�W��w�v@��惹�dW0:�8�q���!愚�f��DHi��U�/�2E �3%�6��G9&�Ұ-�hKo���-&C�b�m"����A�(�x��n�N��7DI�n9��`���+"��̾�˵��ZN���o�����(�m�>�⎹�etM�� �����5G���h͖�=`̾8��^��rTEy\�OL)�X���gs;=��� �;8|n �y<v�1��������Ys�c��#,M��b!Ţ�.�����tL"3��.$��n���v����	�z� ��Nѧ�.C|H�r�ܽ�R��n�ˇ��jq�C���USZ^��T�Y?s94�~ r�0��r5�X�	&��}�P��s�g]�e2�rѲ*)$L����sZ�G���>Gt���z�ay|�{�T�4?�$*��`D`z#QBJ!Q��NZ'O1��I��Ò����FL��ң���R�����{��Z�R3�.��g�U����` M�m�0`Eh�T�(6���fyQ�O0Y�^�K�͋�,q��)�c��/i�kv����>��Z�D���'�A���Q�o��c�n�l�S�~�n���'����\��R�Ģ-�OY���iG�S�6�X��ȕ?���ɕZ6��\hS�# 4g�)Q��B@�@�ֹ�C� ��IV�@M�����V��셴˳@�=��� �N��j
EC1��SҮ'R�	��2��;�J�A2�1��pVGw�A�99��!�[nM���'bʖ��p���wV@��2�(��`���RZo�w�E��q����p'�q�>.�[Y�#����u�F�dJD��]ĠQ�p���<�s�4�a%
��Q#b���'�,��[���k�/��s�-��2P��R}�S�?�����e�t		#Gn������n�&�zA��5��g�D0C�%��%)�
+���"�u�Dс8�I#��}���$Vq�h<�7�:�i2�."?�*9�Y8d��M�Vg�z��@��mc����}x��������q��$�L�E��HsR<;��`Md*��ۮ���ݟܿ��D��@�賃�,wH��,�z��򾩈��O�S�|�D~�����\�1���㕸�!yB��m�j�: l�7|N���"$���R��A4)�D����{���oP��ԍ�N�>Ww1j����ز�d��~�Kgoq"��|�4���T'�z� {��#k�ad��/ZZ��AB�j��1�P����P �����B؞T�$�o%�U�;F?`���-XfR�R�D�1m+	��}�_���4ȡЈi��2n�;e��%��0�؄x�������y`�0`95�Șt�%��u�#���5����4{�_����Q��)��<��]_����ь��n���ēQ�6X�c�$�ɬ�'0Šw��w�)O�8�0;x#��07��ߒ0�복9n��$F��D�̂��V���F�Y�E/��=��-���H�h�礷s��$B�F3�j��B� �:)�LT�A���$�'7��Y�����D�aU���W.�H��6i��7ɫ^S��Sg�7�s4�H����7e瘄��0�Z��^�z�H��yy+�(�Pw6�(w�"�f���yIj��XLh ��12��.Q�-3�����D#�E����Za�����!���_Ya��LZ� Nh�j����{���o��ҡ�I]���ƪO��m!=f-M���4�S�P&��c��z����ķ�O��G��;i^�ʮ�!�;gh����Q-=EdC�w�2�Ou�S�r�8��c��:Ut���L'=�-�
V [�2QAV��P�c�6$���
�Jb�.*���@��Y�*٧�e�)�s�g�c�EQ���0n��ߑ��[��*?Iq��џ�E,����rl@�n3p�囤�h0�d��07�d��(�碫E�g��u����H� �J�/���:�z�����!�׬�$�]ې���F�ڭT���
˙��if��תTsM=��(���x{��QSj2��ش��*�;���0�	)�	��GTÌ��HPP2U�A@��a4�$�*��A68�D�/\~Z>z�����!�-O�ҕ�ψ�E�P^Е~x��`@g��
���Y;%ˊ�=��_��6�t�]�$�.AlRw�k�'|�O�8���d^��«=�I-W0F<چ;��X03��r۱Q ��@���]g�Z.M���^��^���a,�T6_ѺJx�4>.��q@���!Qe�
Yu6�*�죫��3�d�$�:�n��7Qs0[��r7�����[c΢A�8�1�<��z�b`��ȃS�⮥w�f=6�h&]�h�J�>ɻRY���N�� ݷx)�ݡ���W��C�n��_�m�T�E?33�a�k^P�rt��Sp81����'85����+�;����X��G���c������J�)�Y�h��~&�]X@��J�3���\O��H���	���h'�P;���8�D�E.��tB��J�3�I d��bc����wCŞ��_�"�-`���{&�+7����ܾ�6Y��F�pQج5��.Ei'��|��Xe�ߋ e�t���d������>��<3m&��B�s��+x��q2��ԁB�תF縓��ds�Qn[�{you5�`�YY���ƌ�x� 8��O��1�_Sk�wE9k���Ԡ
g���m���\i�� �`$ؔ�L6��q��T��V��$ko{@��H�
���]���;�AB���<I2�����ֲ�h��C�*�ߡ6�%��Y��魫#�J�NV����/Dbc�C�?�m��۽}q�Y�4���k+�L�V5�����*Pߊ�*��3A��s|��4�jAA�gHG�\	y��zG�Dk̷Ka��Ľ����f_p#&n���%�����@�E�B�f �BjO����-�DX� �(�u���xT�Ea��!:��2`Q�R���J���� �����Qg�@��H;WZ����q�W^Gx����z�$��/��O��f��d�����me��2'��dR��/#�fI�P�b��c���V2�[7i$F/c���E@@�Z��_w���&���+^Ӫ%s'k�����ιI_+ 5<��B�		���M��E�zq��@��e��4{��Fz�M湩���i!����kڬ�[�}�§��m�(0��)���?�z��_SM�R�~r5f*"Sh���/�;�g/Q��vMai�������D��}�Nz[!G�^ܹ\��_�km��#3I�uo���z;��6H�1*Ѝ&ȓJ�&փ�^�*���p�H���\_�j/[g�')���w�di�H1H�Z�BBA*%iv]���<�"�5��l�r�)�NU�U=�����ˉDa;�!�ۘ��=WQa�H���<�h�3�/-������@���H�� m�;M��Qq����U|�ҀG3	ŭ�ʤ�?�����B�%�ХX�Gkݨ{ʈ�+�}D`�@i��v���.���c�U�BF�O���K�}�a�|M���ο�M�o�=��kx�iU+0�j7����5�i:�i��J$1޷�4�5������K����D[Y�!Ҧ-��p�~�"
�ǣ"��цa��lob�N���r$�
�� �q���>��B_?�0F�vv�L��%V~�s�!&�i)f�"�*���V�؃3A�/�=d��7�Ԁ{j�p<}L���iS�/�q�)k���� ֞�����@if�o�&�q�	$VI`,��&o_���� o�>d9	��C�:�o���5��渠��S�b~��3�b}�K����D�=5�σ#w<�Xk���t�Vmg(�B=b�o)ˆڋ����Z���'~�۷���U9�2�Q�t*yfMp|���@���	S�H/W5q7�No�{J�ֺ�U,��v����YN0�d�(�	��.��hmAQ̄�u�2��7Zz�l(�_ ;���G�g|A�	�{��~z7�Բ[7z�-Ľ���qC�5�c�ɗ=�IY�8����K�o��rP���T$�����@;�Q���$��?r��چ�m�b@�Y�f�z
�@uc�'÷��k����%<�92p�����T�F�=�����%�M�ޚ���B�˄�{�x�XE��� ��R�<Z.�ڞt�)l�n����e�/�ߵs���5P��\L\[i��Ge���r;�d�#~��%�n��Ee~�F8���:�)#��U��Й����R�H����Ok<�x�9G����O�
^/P��C�?^��/m6��yP��6U�8�E[��s�.K�/��" �YWQ�v�Z��F5�zu목�����pI�Lun��a\�̆��I-��n���ǟ_˰����Fr_&儳_В�	�N_&\q�e�'x�CQ�$�bż�=,ԏ��y��d:�y�1;i���<<(�=e���� ��>����F7Ru����RJj]�������F��˼�m�f_|Ф{�?��4Z�� ����1��g�I��i�Y2��Puڃ�d����4��?���qXyڔ,�Aڌ䚆@��r�4�Uf���'7�aD 0��si�^���=�IuW��si�^��#2�i�(���l����o�U��+ɂ2�(q���´�$�wf1�����vN���ɼ�����%kM:&����_ib_�п���**�$�u)/�Q^��, �t��}�ݢ����Ա[��ۗN�Æ��0�1_&�Ŭ�1�\��RjuӠX�si�՘�;�Gp�/̀dvc8�r6�!}j?�3��E����u�)/<1��j�Fق�?���$eCr��]�=���6GdT����?C$�s4jFq�l���U��%U_7O�P�~�e���n�@/�J8CΌ�Ɓ՚)��9$�Շ���\�u'��GkR[��ұq�)G#Ht��9iA@�w'Xm:n���b��4[E���Yi��o�Y����椧��n��A�Q5Ga ����{vX)��D��"�y��F�x��#��|
�fـ˾#��k�L�V��"Uw״�*��,�<���Q+h�}���DJ4�T6VSF[�22�v�1qB�F�`Ω��f��,�kE�s1�Xp=�^9Y���~�*�
�� ��Li@��L����UF*�?{Pb��&��' 
D��3��|cF]�h A��hM1��*p�>R�Znp%sV�Wۣ&؆||ꂹ՛�V^.P��;`�p��q����&��"�Br?Hd.ד�(�\�"y������ɠ��z��)Ár��
�:�u��N��
����g�W�.FsbߡMŁQT:�<�����T�T��E`Q��Ѥ�[�g!V�(�X���u�奇-�K���M�����BCF;:�;1	L�TV����4����߃�Uݬ�3������h����d�t��&9��A��Ek�gF�@�Q@���K���v�]k�N���Z|�9��t��ݪ@M�u���,�׏_qx����h�$:�&6�����i���
ك+��v���lSm�^��I��V	���۾]r_B�A���&�fD6K�<��u�y�n��oCn����4~h_C�����;+M/�*M�{{���N`fv7�EAU:Ģ����d}���
�{�?�XF$ ��e'/끁���2��� �~��"����q�����s�F����F"
��a�{y��8����&-i��׶Z��aai�����������+��%��t�E,;a~π�%0$`hRJ�%�z�-܇+������64*^�4J��4����3?�����<I�������w��M
R��ڑ����!Y;.XȽ�5��B��֪'�4��=�k���x2�4��|łWd2� ���cK�W �&T�nϮ�(d��)���
�T2���5��{��7VĐĻ�9��1qND���w {�������(������3LK,~�L��˒�8[�F�gU�0-���eJq����B����k�����+���� ����IR@Th��s��K7
�*��<k"��2z!��.������*h'^��,PL��G��P�(�}��{s�����:��1m���8��"��F.)oX>��$�+�k�_{�I|,xrM[��Rx�,7��^j��R�8�	x#g�c	���+���Ѓ�O�xB_%�aM*ݩ��{̽vU��OH��S�Mܱ���
?ܪ�ו�l��/����0g(^�ZQ<W�*�Ǫyx�#�� ���'��8O�-��[��ṁF��X��gR @c�f:�c���F�hBW�Ta��rZ2â������vWO�:��������cl�bN�
�Q�)BK!`�-*��aK�U���m��Y
,hz�%��vi|5fk��P�8�����t�f=c �Ԯsͭ���t���iv��Ÿ[ʔ˺<���,m��0+�%�گ�[؍���S�g�)R,@�q"�E�����;��UTvulU��? �W"'��k���A��ǂ�=҃�J3�^EKx��]�E��5�,�2�b�H�ǽ�>���
��;�Ɖ@V|��7�Þ6C�BLB�f�f}�˝
���
~	XW��6o>��){����Cs`8QC ���