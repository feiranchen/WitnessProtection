��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX����q:�}�p����5'��S���=�(�G��X�~x2�M�����#����?���-�K� O��VB���y�W/�_��8?�bQ��Sn��2+�Do��~߲o�ӡ.]z�k>ڠI=Rߙ[��T�@c͝ɼ)ݧ^��k�\�V�Q��G�6f�-v-R̩QBJ�t�G[
{�#��L�]��Ů�w�W�s�w�Ic#e�PЦ��^���IM2[�ѹ�d��� �p�9 ��R�=wLr�"�қ�+7����#�O���N���e��TŚ)���K�Χ�6��2�@G����[ؚu�o������`�*���'V���7Ȓ�OQ�! j��r���ץ'!�<�)�X+�ev���n�Sp3q��\�N�La��t*b�Q{!��aK��+�£�~Xy�B���j�iW�/JcЊ|�BFnC&Fٛ��]1���
�2)JPw��xQ'�����"�R���.����K�8g{$�瀵��|���*�Ԙ��9��:|����^o��CqKs�\Q�)M�Ŭҏ���m!S��)V%�jv�"���>�맯��hd�-�#�`u��\~�%́'��j@vف4�h,M^����(��+ej�ҴP8Q�W���k`�'�y�=@e\�6�U	�{�Ϩ�2��S�l��n�[~G�US�p�;����&�����/3/ov��ݔ=^��e_�������������Q��s�2rD���F�9�+f! �=M�O�'5E�@��'>�^��e���=d ���Z�MJ��\JU3G�D�v-�(�V���F�$I���]���33�3P����V�lK��1_S<�S���Z7Ţ�7���޺�s/ք����V�����\R�,W�-�:I��H����t�@����e��D�)Y5�.�(�,2�S��[CX�	���Mc��/h�*"�;B�>b�\o3����VAn�Ƌ�D�9�kĘ�w<���2�!��-(Gټ�e�`�'�:ƒ��t��R~e��H�_���xFM�pZ�i����g��
�Ul��<�l
�VٗD'97�Iŗ��o��F�-T�P T�ĔN�P��4���@-6.��4
��C��)��n�7*��wr|��~�?F�qF�%S��Y����J%[����&�yC��ز"?1=��?ؕ�4�=�����GD>�Xr�,o%����f�"%~f����ΛyIav���5��ʵPn��)gl�LM�w�P_$��S;�x"��
��x�~�4]˓Iа��t��Ct`- j:9{�1���s��:?�@eui���h<F���TZ���D��_
�������j6ψ�{>�\z�
V�$hz@8��P�26�T�+��^Kj^�p��E��KR͹9֟W#^��:�]z��z-����(�#������b�P>�g����S!I�Lp���A�.�J�\Ů�÷Z#G"[ׁr�9�v���l��%wJ�q��?&:y�c��hE���ꋾ�h��i�1%�-.V�aC���^��?B��V���H��:�T�n��+���Ϳ�g�~s���K����S���O��!Y�*��l,�,:l�����o�@O)d(��G�&��a\�:��4�{�#�?����l��Y�25Hzi�̗��Ǚ��x:J�67�pe�  ������}<6DA�&���#��*�~��9-u�f|y�Q0���f����	�yS���/]�/���E�!r��]�F.�3��%Ȍ��Β"��S�����Y�*��j+<�X�B�����ޗ����R>%e�w_�V�{'��d�v���5��^0�?�8��܇�&u�,]�?�C*�<-�AVfH�}Q`�
>]|[�"�造%�Tmw�����<��sn�n0qTIʧ�6Dc�����8�&�N��x+E��ރ�v�li߰��`j�fQ��iz����F1�Üo(R�N��D`�럴�O^��38��1D�}u~���4���v� �+W�B_E���P����F&��]gB�$܉���kͷR�(j�"#0w���\)'Lq�I���%qܿV��VO�d�Z:Z��Ka���XM��9�ԭ:����
#��j�~&���~�>CE��B,%�m7��}���e��uO��84�zÿ���m�n�!�[\xt��nÒ+�̡��M�$m��d},Wd��o{(VqL�4O����l=�qZ��:�T��Pd��]�)dOD�sE����ҷ(bJQSE\�@A[QX�`������/՗ʖ��b^l
����i �ķI��N95˖�O�E����5���yk�ҔS���|�~�,Sl{8"��{�p�h�������YxI�������ܑ�#ɕ�B��DQQ�;p�]|[}Xи��͸%Ԯ��E���\}Y��G���2��ӭ����h��G[��`3hF��|�v��3(Ɏ;\Ȝ�$�����S������f�I0 ٭i*��r�yV,˻����o�%t�CH�p���Kn��`u������;�}���\Ɨ��vY�Q�L�=���4@YΚ���=�Zl/6����F����V&�����z�8���i`�ԵEQ�L!�npN���#��.�e1�L	E~ �o������䬡J���Iꌫ!������+Gw�_�O//�����F���=��m���ۗr����`������y0�fbE{O�f��YuIű���Ps�6iʇ��?�Y�z#��_V7^��7�rd`����9SL��M]�<t*j�U8�~Vd>i~@�c� LH�L�����c�%ZL���5�K��-7�+vq�=.O�E\�{,�`@���fAq��ү&|�g.%fe�����᭻K��L�Z�{�L1�v@��lDy6��'��Bm�&��`l`�ԯ��(5ы����:�2s�tP�_�����=�������A�4����6t�_�^���Pf\V⼊i~k�OZY�d�� �r(�\����P?�٪n.uL�ڃ&,<C�y��_B��|/[��[���';��?��D�*�͡ia�v�Mc[c7�>�w&�ge����b�)�Kee�2Y����w��#D�J���&���*����?/be��zS1CH8��$���3�L��!8d�����t�s�*�8�Q-�»&�|�uX�,V�$���	&�J�LswƬ0 H*�2�b�v�o�1[��S����C
" �p�� �\�|ƴŐ��B��$�q(�h��'�A�3�pҋ�ɟ��ȥ�`)T6����픔�Y�*�%.':�S�j�@�ј�a1�tP��˃�z�ڷ�"cΫ�@���'J��:���D��u!A��hh��f+����CHݤY3\��x��	w����)�E`4��z�;Jx
��m��m�a��5��1M7�Da}�:�_�r��ēC��;�4���>ߕ
Pq���e#!�\���Y)kbߣϯ�xke2��a-e�2�I�	S��i��X�!j$���1��~�G�dt횾�.xR���6��0�),Ŵ-z����o�_���l�Q��τ=���Vw�����>rT�� 
*��؃��3�i�5X�w0뽈u���}�"�n'�	�BP5�F]zS5�`p���'���/���\���Y�ޛ�	��8���4����4�Y�J���f��Ȟ(?.������z�b.���K�A�dȉ�{�0�~�s�Y��L�f��cx@(l}������י� ��X�L} �����o��}	�C18Yz]M�s7��?_~hN��pP��]��[6��s-����ܘ)2u��uac{x�k�����)dT����G�t� �-�]hAU����S���������6���R6pUV��W]WQU^ӟG��#���o=�Nnm�	(I�c���e�f�z�R�%`<_G�(��Z�f�U4�a��������yO�0�1 �;ٳ���_y�/Oq����}�m�	$�����I��#1��k��T�ox^�F�j"�A���dӅ���p�s�+���6�?��1˅�P�n��a������1�ey�Nx�JO��Re�U$�,� U�[�ʱ��§wi�5COE��;q+�,�#�:#CjZ���g��OD�S/L��&՚&|;6jƿv�8�3V����ځW���|�� #?k\7�bN����E�A��.P�k�L�'��v6/PB[L�ʤ�og�0�2@d��o��}Y:����(x������ށ`L͆`TE����(���Ҫ�ď(�A��Ea�5u%<wu���C/�ǬA����E�i���6p�Rh��������ɘ=7�����/�3z��ҫ�Y��>@Cʩj�i�ǻ��I��
_�c��$n-���ʨ����+��a:П�0Q�*�D&`%������9�A�b(h�S$s[���k� i�ѳ# L�C�"�o§nq!e!�iOΔ�s�;J����EC��)��T���t[TkM�dW�0	ω�+c6E�	�Ş�g# �e��2`֤-*sp�U��sI4�5?�W�У�����������3	[���bR�	�A;�Ǿn̝$�"RYZ崇��$$�Y�V��m��`����>���	m�v��L�]�.^���H� U��o��7Qdh��4�waE�������}�9�E>��rm�Q5����;ܔ�Q�5��ŭ�-�Xl4�������+]�݂�IF�	��@��h,l��a�B6>5����چ��:�֛o5����~ǡn�����}��P�|��Ў���83��2�'a�D��#�@��>�ۧetK�Y�o�F��Y��[�a��c���^ET�܉yG�D���o�G�j7��.Y:0��ϫ#5��O��2��X=3�Z�G7o�(=����f{��r���kl���bKgs}�)4��݈<�%3��?%�D%7%fH��^��\�9gڡj�N�v���>��*��CE�
CҶ���םR�S0!�o�o�������~���a��m��r 1AԹ�y�]Ff�I=�>�Q�㶣z���E�/}�e>���q����r�q������#�x��
j��ˮ\�*O��:��@�!�I!�`{�XV-N%RM��t�|�ٔ���jYt!�$�G���}��Dv��Fк�0J۴��F���y�o���&:��f=���G� 	��6��G�IB��p�:�k��>Ad�����MI�/zsXؗ�C��.���� b<��a��13�e�)��=Y����|�KgL�	��!.�,��ՀR���I��ZN~��~t��5�A娷/����:�^��/����c1u������Ͽ����o�y���SH5����7F�k�З�so1��y?"t3���q���;l���P��KQ�aF�
��Z]:[�^�@����m�F2���S
g�d�Z���3�)�`��f�CHcm���&�qA X7�Vh�3�2���S��A�X�_י���f^N�fP��Y���~\,.�B�<SM}�p"�G"(�"Ӄ��9�W����/���)OB`%{c����J�{��x��"Wwl�t�pN��)�Q7�D��/W���U=2&��v�
b�-y[>�ELwog0H�̭�[}i.mcg���Kg"��B���Ja�!Ȩ��×*�"%��>�*(���3P�fn\���H��E�
�g��,u��&�c��3Iv59�n�f��at�m<a#.A�J�)�^7���󡗩M���K�0�9�#W�њ��<����g�*#�AH�_S���������Ec�.�|�?[���z�����Yq�p���$�R���/��ƨqA��=�P��7TV�ײ;K��li�f$���.*�A}�}㳕���dM�(9`�����Y)��Ɇ�Z�Ͷ"�^Q��t
�L����{�j�J��su�X���sw;�l�:�
��mf�d��8����$;�y/���#M�\���GtV�����]��ňʽ�@^���GWCF���h�g�%u����fՄ~	�ڡ�&�Ι(8�<�=��:)��lw���{qo�7�d	f|�a�����7�n��\MW�Q�pʔC�.�󱶨�#/ƔS> ���bXH���:����~�=^�����`Z��1����o�v�~����i(���yew9U)�z޹���2F�Ct[��lO�ncN��03sr��*��Xѧssw����348nuߨ�;䖴��v��갑l4�~�߄<1��4
�t@�;�7�Ry;��(�%����Ò��B��T�c}�ژ�6��?>s>��F����\+ۺ�F*�l��?p�H��&_�Er! >�!�K�篮�}�_�,���rm0,j�S �	 ��t"�ba�FXg�����Y��2�*B{)O�Ͳ^��Z���~<:Z��Y����Di��@����I�aD
Rв��f�6ݤ�������ec���b��y�H�����1x�ʔ�-���������U��p��%g��U��K>7��	U� �	�D�����C@Wb�\I\x ���^�D�='<^&OG�W�B�66<�_e���耲	 Vf�������!%
2��>�%�Q�a-M\��$�/R�`a�}���k��
���|>m�b G���HX�8p$��PD�FYnC|�;�h�M��QA-�C���3f�R�~;�%a[ʅ���lm^��ߟwt�5G�7���X������vS�g��I�����ynή�&�"�q�&�%�ص�o�/gc�]^�q���ԡ�p��#S������{��F/$P@"�`��Wl �JsP���8�!'4eG�%�Y%��䢫�B%�(�,,��	�����F��My�h���j��CdB-b~��JX; �\"V
2��7�I�J��G�K
�����6%o����c,�c�A"&%G��d�;M^[�!�V��oZ"x4u SW"ǸF��2Ȕ��l����� �����L��{pUY�d��ҳ����\�tV4"3�&uޠ���rf|���P���9�2�p��"�?ފ�~w�2�b��]'�%�Z!N�l���;��i��8E9�<�7�ʯ'3*Y(8ۍ�#�{��"R��9%ΉP 
�����j��C纘���qk����պٓ�Dw���	A.X��������JQ6�VU�[`���F��]`�q�n�M��(��˼��>6f�����?A�.��P�/�oJ�|������(�',l�D��i��I���\2��w���,���ɹЏ0�g�Rb�Ehʞ��u������a��������j)�!}`t�T�BB�z�j��kO�z����&�9Q7i�~I��	�B�Y_��Ã��q�y�����vL�ZfF+SN��,ϭ��Q��&�Ta1�P�u�����e��PF�z?D�l?�eZo5޺�@�7�I4�|̮_p��	)����l�j�S�ut#ax���鸍��F����i?�z��UzWB�V ��e!ܸx�]�"jY�2�!��
������O��������Y�?#�E{7�j�����f�]���.�o�/�Q���݈����{Sڳ���V��a�M���<����UA]̥ՠҥi�TFpiSI
�l0����=gʗ`o}a�#ly(��`�y��E�����Z�p��cQ��3@ن�]�/\0л��(3|I��'`�(Y���(�ʁq������Ӛ��A�JI��\�6����"��B�3�f�,S[(;4kQ�,逼�qc���1Vՠ3��D���@z�,l��@ %�fIy
&3�R$U��j����f�h:J�.U=��]K�j���;��#�e�1��
�Uƙ7����Th�Qq_nW}i9)�z���|�L�r)'�@p3;�q&�9^3�@]��9���K��Y�������Cui�,�;T�JWr�a-6�v<�z��Z(D�ᠱȨ���K"Q,�t��fAo��P�-ċN��s�