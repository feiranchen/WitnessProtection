��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��g�߃�`Ɯ�����ڢj�U٭�HD�s4eH����h���F���+�9~���qp>�0`����y~�~J�.�J��^��q\!��=$N�����3G�ψάV�#\ʅx� w��پ�n`L��,
ۓ�D[�qiA�SVڡM����-��2�M= f�\̻�:7�:ǧv^O�'��,�ā?��q�{+ɂ�Xz��$�+e�1<S;���tK �x���@xź;�y#v��IB]�7?�n^��O�1d]I��Ğ�껽��ܜ[��M�U2|��u4S�~��k��~�zH=4Jm9-N��7�����	A���w����%8	[c�a��%���t�"�pcs�-���ŜB�@.�W��]T�?l/�N�cO�`��8�奕��G�0֩8;����ݽ��@|�7%���HF0�Y|33��´�Trm��P/C�?����n"
PVR.|ﰰ��ypu�e���n��8�S�P]�v�'��"����\����`�\���'K�M�rp/���M[:����10�N�-�k�q�yCD���QE�ƾ��-�D����WD`3�\7����k��@��Jޖ<<��#����|�>�E�D���ޢ����L�0+� ����e�}-���­4;7Dw��6U��Ù.���I��uf=,*;K#n)�����EˎS��D����O��Z�Ј��͝.V��>��,����^\�`La������N�\�͛�򈱇�u5ڎ�����OX�B�WVꋎ�!��ƃ��fM�9wY�Z"S`�k#�NsV+�*_ʅ�ʃ��˚�`�9���CN�z5��u2�k��e���������ҹ��Ѿ����l��?�I�dx+��hl"���8͗��J�~���];�i���6R��Pl�|d�0�'S�hk�WIE��-(dx�k衔��$�����屼�>n�R�٭3�Z"��K�ܳb��%������=Q�I����t,o���<�$0Y�:�6ߞY�E"~)��"YF	Nk^������M�kK�_;��q��GH�����ȕXi�Ug�;�6��ܔ7�YeIB��G�1�~��\����:��"&�j����ǩ�/�r6TbW�9�B����?*�:o�D<��ַB;���W��V���H����?hX�ػ�`�4�Q�*�Ƽeev���v�-�w|�����oq(�h���I�k�����o���tqt���_��br߮�p*��XZ��h]՚��u�i�-�Q=��i�$4����%>�A�L艚y�����u[φ""'~^~���9!ە�,�G�@){�tV��&u��kF{,q���FM��9]��g>v1.@F��`�x(�L#��<�`��fc!��[~[ħC�vC�Oz��seWJ�.Q��_ԂjN�H4W���i���n���(w����}�X0�,��h�Co:��*`,��4^�%jL&����	ĠNZ�6J���p���o�n�[��%9��jD8��B���2U���mX662,�`�@����R�d���a��D�61���S>R]��JH�o�3��˷�G�h��9��}�ѐ����N�Y4�,���.��� ݌��Ofnfpr?� �Q�=���z���@�R!;�T���S���K(չO��)�QZ�g�`���Ao>C@���i��h�[�2a�m�����U�������WiZ��r�����JN���!ؑi�$V�k)�{d� Ԃw�O������d�V\��BJ�3��h&C�Ď�5��m0 j���y��V��P);8mAsl�6VӹT{~��b�k�a����@�Rk�J[D^h�2�Xu����hy,�xb��Da�O�k��M�g�7)��E_��I�i@�� &D���q��~�έ��3���8Fm�a,v��C�+EqR�ut8:~@K�㱳� ̷5���T�l����m.�W��}5+��X �~����	�1qR'@:q.g���q;j�Z��:3u� 2n͑���?��>�����eo����k��@SyR?��p�Py�&�;���d�^��M������:5�5�H]L����a��5;��d�p�"o�`K�1����g]�3=Y�\x��[�ސ��E����7���['����K��k9zOI!��n�oL�����?M����5v���;3�>p$!�i
�oe��wp��l���D\��e������N ���wh�_�|�� �S�g1]�hz����x�T!�5�rhi߽uB G�O�!�3�-M� ��N��nV<I�B��BGUAh��������g�����ȱ�0����Y�G''�30;%�؞E�L �`�q�v &A��3�&@&|���C�֩����ޭ����#���Yge鍬����]�s�?#�e���/�PlZH��Oj�!8�u���C��!՜��Sd������]�H���	�]Y*��e��!�^���WNb��Hog�QU��8u���"o /}�K�Q��O=�ʵ|�LWbt�$�o	���g � ����?�=bb�`d��rJ�ze����8a=9�R�N4�z���9%�nD&\�b�M��+�;콆(��`���yǛ��*���Y�17�[w%��)�R�!���g��������i�\5H�+��L�N�q찯�`��36;\S5��B�*�65w�e�E_Y[�4��1!���$����e�z��B���0m�Ette�]DH����m7�I�n�`%���L���+�%xk�D��o�ħ����d�{u!K�h�h��%r��(q�3��KpS��C��V0^gdA.-Oo,�
1\�S�'wI�ޮL]͟�Ī��"m�^����ŅD��lW�uQE#(�4�E)b�1�/�R��ʋ��+�9�*D�i�$���F �~ƭX�6��";e�N�h�h�3��R���>�o
�60��(	gs�|�u�r)~7"m�_{k�w��O�P;C��ڈ���=����u�t4��7}J�v�xHk�BY�ƪ_t���i��..�,�)nPí9S��x���ӊ�!�stYt���#:�}|PMWz���}F���qgWF&8���Y���Dqej�O��ˎ!�<���u�����ĭ��!Tʨ3��]M\CA�Z\6^� EOkW�R��� ��h���c��� �`֫ ��ݪ[8�C%�E�;L�+O<i����)jM�d~TB���^�rL:��n���CJ4W��P˜�PH�B[ȯ�[��jO�b1�%�:����[=Օ=�w��[;���8<ix|��^�v$a��ԧ	:ܽ����֮d��UЉپ%k���ϸ�fk�&F	����)L�)�p]HR"���	��l���y�j��v>�Ї��` $_ٖ8u�n�3Mt��Ϻ���< �ވ���[���)LKsu��ĨvE�IR9I�a=�����l����d
l����Kc)p�*׼:\z�Kj ^��n��nO�!s��K&�=�T�2��QL��
^b��`���� %��G�]#���xn�j�L��u�-K
���� r��E��^�<�v ���.�n�e�sO�ф6`��^;�^@�j��ヌߝ#��%����ɐz��b�^���oͩ��/�k��X�\,bb�����5��c�r�Ur��?v��\ 7���`�%��I\˼���(/{�<�g�᫨2Q���J0�M��u���/5�����B-d����&�(����PAӎ�l��Xl-�Rݚ�C�z	kq�)�Ͱ�a���V2P4�~��?�P4�+���[O�3Z�ZPD��.;')�A�A�+Y"�x�"sc,K�6\U����-&��<��ԫ���Kiܭ��b��k�3Z��)��h?�t����4M�t`T5� M=H������c^C�v��6$6��c��@����G��L�Hh	h5�c/y]:�˪�������j�-7��L%���S�C��˸W� 5/���V¶����H�t-���r�C$+��b��0׻��{Q&^k]� �&Z�T!�^A�L�'Ԡ�
��K�J�����W��V�W���B����	��
�,�n�5�{�/t�M�/%`U��0m���]#\�%H�����|D�.��q��;�՚�s/�C���ث�*���Ci��W��p�?P:�R$�RJ��.}'����ŀ\3�e�s M�
=�gF��^b�U�8@�%��>k��H��"��ē�G�����F�V��}��
��Y��?xK����T�M�z�al$�1�$e�3�͖��Y�te���?��7��-)Fw&�^ IP_����E�b�EFܠ4�{��00�j�Y
Y�%�Jw-��v�R���$��/���Bώ/���h��-]?������Cg����1]Lă¿؞b܏P{�[4�}Ě/��i��u�~��|��\����z�M
���m����&����v�`!C�{O= �B&����3Rɀ�y+ � W3]\9�2:z�D�_�צ��MZ�q:��I6�\���	��n�J��嶎����`��x�f��˜t0-��B]������䵻	ǌ�AD���X��ˇ
^�
t`�zi1���_�oм���!i���%p
	S�������4������K3��{��#� 7[aM�#/���)�ZC�}�8��u����HP ?�hL*:~��۾P����mG�j�[w���/�.����a�P$�����!S'�D�Ft$���Ng��*tIޠ�x�{���:rv�CTͦ��H���P���Ǖw"PH6�=*�8��و�6�U��a�ֹ@[��f�6($yk�(��!��{D<����>�:!j�~Q�%�a�z#n��jn����
��ݻȦ����@���y�߰�ڒ��_��n���[6N,@H;�R*ȍX�)@�u�W����N�΅A�4���@�Ԍl���S��z*d�]3)]�X"���YH:�-e��rA� ����=q:{�l�i���r��(�b�%�6P]%�a*2��ٜ.�%�z�P�lhA�.��g�?,O+�:���KOj��L�[�Bs������O��N�6�Vr���`�$�G#�/���1��d�݉�H͹˸�a?��'+���^�*��U�R�9@��b���FJ��M��x�q�( ؽ���n�	��r9�Z1q6�`S�0f��EY	^n�2⪽�.�� N:�3^;��]�7DJĥ�ԅ���cih4U�C�&� �2�ֆV�j��/��χ��T��PT��?�r���ؑ�i�5�z�ե ����aX6�}+���g(e�����[G�tQ\��X�.��C�Zc���	uV�s��lr�6۞|1��G��i��\���s�\I�7KB!���䝽y��C3y�G���`�h3�����`��O`4�i��:����	��:�w�5�W�*���A4iK�i=�ѓ�`K��Luə�j�}*����N'�=�Z��u3e��Z���6	t�a�^Z�8?Z���keL�����Т��A��|)Sv�T�6h$�)0E���L�_����B�	<�������2#��e2��żx��E�]�=���}	y��@��h���[�s�D��c��ᓱ�%�D�6���*���bY�m�>@�$�炊���`4Ճu2 W����	�L3��U�>B���>�Z�h��eD8�H$�(���[=�<oU�EM���&�酝��0~�TC�o��F}�{���u<��N��j�W�y�����x�8y�%����KZ�0F�X��V`��}ō� ;@c�g/��<2�%ˠ�#����8VT���@;��Y�y{����@\�`5�t�K�"
8E��##�@{37�3��eJ���?��cV���F�d����Sʨ�|# ��4�Y�d�M���. _�Jr��r�[:z�<�C�!��H�&�r�d0��P�6�R�קƇ�$�h'�Wy,kz��oL���U���r�É-.6�ā�C,!�^VV�T[��D,�ca�:�hl������#�H.i�����N��͓�aOf����d7KmП[�a^c'���<H�W#<���ؽ���ǙE$��D�# �&����g�A�Kf$z�q�|s� P:��Z=L��̓�K��� �Mx/c�3���h��6r��6�`ґ ̃�m����T_�a9K.�{��"�_�nVb�p�b.i���������%:���i�4 y��K��4�#:�M��Ĝqc^�R۠sŨ��_��!!CW�WT�ɶ�I����iҳ�g�ƠR���
FRV��gz|YQG�fb"��КVC5ۼ'N��h8�޵;�׭X����o������2J��m(�Ė��R㲬XB�榔�r&(��4�h%dţ���S@ '#��D�j�h���g����=-���g_R4��Ōdk�i<X�"{�S:[֝����]���8p�6�%TͨsM��A�tn����/��Q�_�� k��5T������K��$�=�Q4��� r��}��PJ��чm�=��Ï�����&������N�'����U �@e�}M���ק��}��}_�:Wњ�;��Ye�ku���f������b�f�ڇ��1��2f�i�~����R�H%�;�
#>���#�S�%����я.�Y�;��C���Z�����fg�'Lb�6�	}[r��)��P�T���ⷥ����w���uT�%�L���j7����,�ӣ�O�Ė þu�����-9=�Z{� ��/�$�73����ߵ�W�Q�%Y��]���w�Rqw�I��J%�x�=�Ә��v� 7, �g��m�|�SCKDW]��YB�π;f9�Tg.�Ex$���Z�����)�^
n�_���������<���U�1q������X�7����d����5ܣr`�:{ 	�Ze�)�\	n��'iI���y�����)���h4��^o����;��(C��(���G��.p��F�H{��W�8ds*��,W�PW�I�&� �2�Ԭ@X.�pe� ~`���i�2�Tjk�3�$g��#���%�E7��3����a��_y틸!E�s��C�\yD4�F�9�c��*Cd������g�d�@�C�L��{�h2 Ȳ��ЋV҅�T\y
F@}�-����В
Yf�.&����gj�n�~<��*��P&�cLt��X�:����r0��}��5��ͭ��p�J㴦,ܮ���Z�m�G�o^樭�j��i����/���Gz�ki\ %�:�� i�@�u�`^�y؉&."4 ��B.9Ó��V��Y���t$�2c����|���J]o'�on�0=�2@���������ű�Ch.�����q-�:V({��@�P�
�v�@^SƄ���c��/��9�f+��T��[i��(�}�JA6�i��O"Q}��5�jUȄ�嵞�0���nQd�jJ�U9��aa�6���_?����/�m{.ö/G��=?����L�m�M�.A*���]#��xk�z�����IY��%�v7Q��h9^�^a$�	��[xҰZ{v8W`�>���^�k��!��ڰ��<E��Ɋ̣?�o,*�N��I�Я�Bo���/�ɮ^��r� <�Qї%��X<�@�D�t��`�Bg!�&��A��¤�z�2S�1���4�Ļ�Z��z^58��t��
SS�Hs>�f�ү���1�	�A����g�|w�e�@�7����4���W�c��Q��&�3��"�DhS�����BС���.�ᑴ��3s�����U@ɉ4�� eQ���@�{qĳF����J�W���iTj>r��^�0����@��;�s�V,H��[��+�k��~�T��W�5��T8�)~T���q&M*s��ݼ�F��%޻d�y�*�_��xEv�c�������r���J�<�;0�YXXi�<ׄS��rHZo�	n��{O8~�XsL4@�^���HG����U(��!�����p���~b��Q9�e
̽{� ��l;�:
���e��9� ��=3�9ߛ�z$�m$�0slS �[�|(c���?���#�C�!ohP����J?��kڛn\����A�I��RA 0�Oc;~!�$vM7�	��~��\AB���?�Ń طMVt�Af!���76�����8T��n�PǠ��,�t��)�G,�T9��L��� :&�Y�=I�"c�F��|�d?S�jc��fO��+�W��.GW��=w�ff���B�P 1��]m@���֯��Z�k�|;l�K��5:���_��15Y[~�K:|ꡮ�x�ga��p�Cl6.�lak�M�
�%��վ��҃o������B�9�4�7qWxTi���z������R��͆�Y.c̓���|1Y<P���vu6�%�2|3�mF2�]����)���R��-��Ƕ0�h��:>����'Ӂ�V`�u~H/�T��d���)Ap%��z��䡊X�wx������O�_��V=�_z�jP����iƧ�,Ȳ�� 4ֺ_�I#�Q D��Jұ������u:�`�W���_�!t$n[��� �P�Fa/�f�d��r�����z�K���cu�C@ yI}F���ӕc�j�Q���R���6Q����_�Wܵ	���h
�5M��V��{qc��n�����Qu�J��T�G��>��[D��8������õ�"��?c�:��j�=&�ծA5�\�qO�>p�G�q�d��ښX�R��P� �W����f�%������7Y���7�>�pԭ)�~+���>ߝ*��'j���?��KV�0���9�9�y��s����@[u��Ru��1@�Z{��y�#P�0駴ion�|+��(�3��c�G�	b�k�1�v��is(��)@�tYC'���9b`�a� ����Y�G�#�`OAd�'�Bm�Ի+�ϰ죍�kSS���2����l�(=fm��`�NJ��Y��(a1�C?��,���356 �'�N6s��5[Uǲ��cY�������ꬥ�N64?�����̹�b��w�x{Ǫ@���Ǎ��s�$6�߉6�h ��:֘���������Z�ᙣoH�յ��T��r��-Vov��`K�q�"H}��
|Æ�ۀ;6H=|������2%{; ao��Ж)3�zH�#�`��5n�-l����(���l{�}An�U�3�V r;f+���<��/�5� u�~Lu�g!��ŷ���d�r�v��I��DM+�gb���e����S4S��`�=>RG�y����H�I��]����˻�5{���=4R��	��"�o*���3*�*h���	�=�M�[�{Do޳�wp��$gM�dQ,7�6ؿD�����~�Īn78��Q ڋ��M�Hd;�%?��R�~ Ʊ����e�Q�����"8s��e���`gt
ˋ_G�3u��2�G���-��|�iI�D��S�9�Κd[y�z�k��1��Ԟ��;Ǆ#�ȷ|�fꄳD���i�L��PL��ǀʑ-��y2�oP����Bk;��U��
z�P�/��)k���M۝!�?xF���fUG���� ae٪��3�CQ�+�˪ӣ�`F��:��J�Crn?��_{$�S��7������0�-G|ܗ��u��7=���x��=�N0��󭹈�q{^d�b�M;/ @�Jl D3��- �`��B<gb�LE�V$^�x��o%�Ƌ�]��Nn�I��晞�=���������Ыj��W�4O�',;��^�6ԧ��7R�`�7���3��q@1(0\���Ip�$^J�^��"x'=�����Kct��H��h�%|���̠?�%�^�w��ܫ�	�\$43	���1�@���{���-eL����J�8o���`Z~|�`R�+�{'��6J ��2()��H�0�����N����J�$Q��@���7UMW�B���yS��z>�T��:�ך޿�U\B��
-n�a�w3�ާ��=gq>������eVF�u� �S�����E�G���^�'�2�B �O�܆!�'b��Em�Om	�����Q"B��Fd%uz�<�gxVaʢN�\J���n�=�~��gD�˝T"Ե�|�xTf�\��A_KRh\�0�㷼��j�݉�1s�]khC��Ҫ~�,���Ù����|��C�̽�ӻi���R�Nc�S%�GSRXTg������Ԇ�������4o����E.cxP}����,ε$ɩǐ����mtNC�<T{�E��%��(�/�t$��ɟ���m�Ԋ���>{�a
d�~~��?�r$�vEa�t�����ĈD����5]�^�h���^���g}�Q�`.�i7��0ͼ�o� ߷�ٖ7ǰ5>�����Jeߝ�{���l�<���E� ��f<���,[���z.��:�^�)~e�#��D��Ny��2U���bA(d�D�Ҏm��E�˿0��x���r*�HDR&��Q�)W��,�J�����E'���������"h�B��1)ZK%�Ճ��L��)�0|ξ��o0���������w��̉e�r�A�3���*%��5�Q'���m���c0�5�)Fc0��6�.��hN!�'�κ��ʾ?��k���<)9_��QZe�@�Ӭn���!��s��r�~`�Y�lB�O�g�EKR���g�}8�7��my�ǿ3�7�AW���V)�=�����O��:ƃ�5'-�qg��P��)4D�>Y{�8�n�[��Y��'$�=@T���h�1����יִ����b�3��C@R���8�]��;�V�S���i�bX�M�b{r)S��JQ�,R�Y�"ӆύL�z*LK^�/���OZL㭇7�q�$�{iQw�޲j������
�S[�k�GI��/�cK
6��5Ƶ��� ��08KhV뷆٠=ٖ�ԓ�xmq�僀���F��]�+�Q?��䅼gNW��G�doa��D����'��A�v���D�jh'0�	P�*�[��y���'����i�1��I�,��$��@ }�y���)v�'�H���P��hx+'э��`TkL�nu�َ��JAcI�n�v�B07�4��rpB�gMA�a�W�,�(�T#σ!�
�J\���|(wV<0���Sj��2e��&1z0�+s�l�ĸV�
����_��wOs9t�l��d}�;p�\��)+"��3�M�%���Ԧ.q����8fBA�`U����@r�+��K�'�x��I��⇭R�� ��P�����0�2uy���<�Á��%)�o+s	�o�Ã��7֥����^��_�y�`�[	n�ַ���v
�|<�C V�>�ʁ�����E��f������`��o��:y�lL�����u�&����x��_�t�8\W�@W��m����	���y$Z�&�0��Z�HA��@��>|:�����gd>di���t��؟�F1ʩ�k����1p���<�J����	�ZmJ�J3�\�^wf���Ԇ	F��c*���W�	��� CN����>��n=n���ˡM�A�d���.�j�$����?��t�M#X�}�u��a8��E�]xNZ\��w��9D�fy��1���n�	�YW{�ܛ��&��,XZ�WD��w0m1W6=织ϸ���Ar}���X�"kq� -��bh��0�xi7ҝ����`@��c���ط"S
�`�	�/gR����_���g��� =�,�ƒ(�'`)?�$ܢ�'�������B��l��4 �n"tٽ������C8��&�o���7���f�&Q��2N��ڰ�6���Y������'��@Z���1yX�y���ܲ��Fn��U��w��6anv]%,���iY�� ���������X���$�(n��H{���ţ'<��X?ms����c�s��O"͢��Q5���cB�^�t�p]H�@#,���f)1��?�o���Y����36�Wg�����/O�4I�"���6�sk�����Ocn\�t�C�ʜ���o�A���j���)3�5�*- oL$�b]?��g4?�/��8�{ sɻ;�"�v�x�w�*q����?ξ1{�y<�A=�iф0���}�e�� �V�镛�a�C� ��~:p��ʖɰ̣�K�����Z�ph�(��]�5�1�ݳ� [	n�n�(��HOcY .�-x��{��Pm�kq����Pmwy*�IQ�D��p�P|�����7�R����Q�
��2K�y���G�Z��I�7Q�ZY�Q[�Wь�q� _s��4 ��!�>���y7��(�v�VgH>���꛷�����r�!U�6��x�m?�%I������r��k���-����{������.�d��+�W�0��-�Խ�h�j�]H�\L�	�7C���l����Y���FlD[;�����	;Ls-�}k;~�߻Q6�9G@���%�j�C��Y�@��R��0�*�C�I
 �?��ց1��Ԧ�kO7�j�C���y�F'��Y��ݗ,X�
�0 G�]ᑥW�95�f�h��xnA�΃�p�)ü���H��I�7~(��~9��F,��Vv� ���C���8���C�a�䓶�Í�	yv��a `̘�e�]�����:,g�$����B��azpG(pI�����ټ0"��S8 o�+N���f�<}͏��P&��ñ�ELF�'#���?��3
�P���?ڷ̜.z�@ԉ̦k}H^�Ĉ���g������7��b�;,����e|�s���@1��v���2�}*К��0�X���*A�`��X%���(�C�|<�l ̇
��W��I�K�x�{��o����� ��Xcz�Ñn��� �N���gGX<�A�*ya�vS&Emy������A�Ȯ!�_GHס�����j^�M��A�A�"�p|�eP��)PMsdnN6�m�d�bc�!i�v�ۜ�}A^X��`��}���%�;��?&�ڳ*;�cA�������h1&+�c����_�d���Q��XƟ0���BiD�Mv*���g��l��tO�1Jpgj��Z�`W��L��'BO�ȏ�t�ʒ��<|���6#�\�S�3v7G�
��:H_?��Σ�H���?�K�A���֋�=f���>V~W}�p��4kn��'2�[�WH...tz��(�u�� �~�}:Pcͮ�\m"jS{�%�N��C�o��gXꌆ�J|rd�FMd"�h)+�Ȉ��8��8��b�}�k��v���-�c�@���I�M��ZsI�u���F	� ���	E1<m���[e~����*�嚂���w�D���^8L (�i[R�@�g�|����'�)-��p����z���$��>�轜���λ��P�D���bh��������ز	y�?��D}��W����t9uxR�w%�I�B^����%��γoaA��l ��=���Alt�����ȵ_�u#>u�yo�M̝e�]7��Ct��%p�9V��>F��T�Zz�/ʕ���X&�4:�gއ�^���I�P��'����?�|u��C�Σr��2�^1���_AN�f�Y���i^�	���1"�ps BSy�˺Mڰ�)k,��w��t2y�D�BD���h(fS�z;Zs3~cH�͝�v᪰��"`��P���zG�H�O��xC�/�6/�)���^�ƈЂ�e���t���Kך�<�xQ]0��gQܙ0�@�]��f!�����,(�uy�N�I�F�����l�P1U��s�$�4(:�S����3M���C��I�~|M��=���Q�:ف�o��s�,.���QBsF�+)��`���g̓��n:rg{����d8����[i{��dC���
}��$���y�rJ���]As�J������[����G�oH�=::�Q;�2���A&%�{W�6�S�s�;4Լ{�C!f�S���ȧ>� �7�>�]Ω?�v(;�]���M��oix-�h	s�g�v�������m΁6��^�������%�N��W�q��;0�q�KS]������^j�f��I�G J�OQO�צ�m��N3�@���{H�Y�B0*����r�U1��Z�g�Q��֪���(;HksM����	 Yo�P	�FT���gax2�,�`�D"J����C��2սO[��cO�7af!��	R|�k��-U�܁�UU&����S* +���V]�œ��+���0���y�7T,]��.=Q���@Kw��Q�-��+��T�$K�k�Fl{��h�ͣ��8�1��#��5�Ͷ	E��&�Q�eb�ApeTf9u�;wN/��xʎZi/D�!>�Ԃ��·7֊(��KUxŤ�J^���ץ7� �YKi�O��C!�ݤ�`Ն1.L��ݝ�.��h�v��$�q׌m�������n���f�i���r�B��y�eWh2)4e���h� �`�>v���6��a�t�{�
����W�;�z����݈��p�,f�S������oG�Y�����Q*r����:��9��g��\%9C7����HdC.8�@p�����>�F�~ ���fy��4��Aa֞`�����e�7k/�E�P0
��cs�:�IN��X84�&���:�N����#�y�X8;]��:@����N��"�_U��N<+�s�`3t�U����O��7�lM/r�*.�9� ��l3�_DDF:�����&h��8���5z� ՟����;���zD�i�X��*��>��������{���FJ��8?�(�1/[*�C�A�18���q