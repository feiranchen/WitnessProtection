��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^(Q�`QԤq(�"1d��_��M�oЧu�Dt�2�3z����.�`�9��8I����w�义=� ��%��3�<w�ce'�j�A3N ��>Q_�1*�ǜ���*��'�G�BL^�#(��xw���ʉ�T sV_UC���9RC-^Rǽ��;�E>�h/3E7�p��K���F/m��:|�FK�l:p��ZvH�YC��c�a �~���E�O�5nʭWv�,�����?oB��h2�UЩ�*�yr��8\�`K��l��p?�WK�t`��bis�� ��9��O̢~�x�W�s;��4�l�Ȱ�g)�"�2�^���v-�YYB�Uӣ�Ԉ%H���f�P���n|��Ł��#���	d.������o	z���P�׻{��ӟ��48���-.��S��d���#�Vm�_F� �7`����SODt>)_�ZT�&�S�g�I:YS��s�] �ýW`G�I��Ow0z�B�w 4k��B�@7�|4��5.�(o�MT2	؟/�O�9�y��h�\���v�+]8b�u��n�����C����f�2�����V�KG��2�xc�i����n��WvK&�;���-.(��|A1�%�ی)�nu�
�3NN;C�,��(?yR�b��~�wP���'����������5h�^o�aS/��I^7]�~�p)@w�5hZ�'�{��6?�  '�f�U�7=��[���1�'Z�"��h�Ԓ��\��}U�2��d��0b�~��k�}�m��&�^���X���Z�A+�]`ۄBV�l,�+_?��Z�G��>}Ga�(�m�LD=}&�yc���	S�P�����OxZ�y��cD6��e���Y�?��g.�'�2�C>�@��j��>�dH�H�/�N�(e�5΅��8���	�?v2�+�{-]�>��м�oe����������vɌVJ�A�Ԫ��C�r�.�E���>$D͵y�:�VOf�ȋK��z(�3E�9�1��FS�����ث#YSs���'4Mϑnm�Yhஆaf$��D��H�" �����)`��D�Ѧ��AK�y��5�1�N"T S��%iK���|��W@_�E(�"���eq��L����1`��z�/��Xq�`n�����mp�9�`Jm� ��b��AKBV&P��">�gp�q���x�߮β��"�E��-�JC��0�x˫�Ka+�N��֣S]�4���%c��~}�5G����e�Mt����39���8�oY�����6,Cq''y�=Zi�0�{VX����y��ABߡ����K��4һV�!�G�J.���.�����v�g�D�gy��"�_�`.�"YvXM�ռbs������_��4�"œ`t諁nd�A2��j�5Zʐ�j�K=��I+�e�t��A��h�7jnD P��#��7�#s����d����<��;o@�-g~��E�f��q�2(��"%�R^8�J�:��T:��@F������k��2+%M;�`����U�t&�MnnrW>bU�{l#aY��J��&Gh�J`����^���ݲ���~y-��sj��Mz�s�W��^AD�?��sԯ��Ŝ�9����@��} 5y�7ZJg�n��j`�0�PKK�Y\�)��NX�*����D���F&��p
�v]s��
��N'��1�{�0�J!��dYU�wJ�Ze���7gh��;p~�� F����Z(K>|wy]�?�.&}�M����w�}c��R*Lq��%NP�:q�;��X[M���Gր (5Ez̀�^�6��ī�?{a7���֧,}���K�)�u�KW��&؏&�i�p9���$]�amu�AQ�\��83�ӡ��mEh��4a$�w��Is\�:��C�$��#�9�X�5+zy.�J��&
mt=�/���R��S?Y��{��0:^ �q�p������]u�P����ۡ�Jxm���XeY�C r,�m1�'�H�Z��Ld1�.�tp{�FKQ���������vYKb5�����j��T
�����f)��bͷBw_%%<�A0;mV�چÃA�K�f�����@�g�����Z�=t�
f���j1���o��a���g`�V�r7NƷK�ʓa�c�W;��(`

�����y"w�RD6P��.��:���F0p-���mA��&�}q����t�Ydh��V�K�X<!5w"88����0�"�yD�D�Z�x$Q"G �D�\9�\��z&(J���qZ���<��L᫭֕��PB�e��an�Ϗ�YL�bto�͹��ǋW0�!���u���c�%�bhS�u ��"vM�bs�aN�
֥!��`.� �V��m@��3�v'�~C6�r�Y��F��I3{�߉޵b�'VO*�O8��;y��O�Z�r>�-��Gr�|�<�h18&����^�>�<>���]��Z)B��-��po�e�m4+����w�WȘCh�>$3i]v�g�����ޕbhFzT0�djͽ����/&T�0�!,��F�S���7׃�n�x���!�@֌�F�@�a�FS��(bH����p�i��:�6��P��w�Z*���eS�+Sj

�]A�s+�a>,���Ű��^pc��y@���V/���ӞqR> l�j3v|`���:���?���ɥ�]�Ǐ`�_��<;y�x��3<O����8��
)E�L��B*b�3���zܫo���~Je.�(M�X"WQ���w\�P�U�3�<�v�k�z�b>�-(!�*�s�(k�A��C��!%/p��hgDX��.��4��UW\{��Y�|���ť�v�/���]���ـM��ͨ5x��ϰدϋ+~1��� V�A�:��KA����Z�,Bc�1Mja8>\�
C�<���UF�O��
(�O.���x��0.`�a�X���=�%5�>��HxA��/�=	IZ�9��{����BW$!4��Q���GUH��Z&�ܙ1Q����;��U���yx�uE��7�,�
�j�Ƌ]B90���I�tH~ �3��h���T���U��.�ӟ���T�Oϻ{�D_h�>� �g湦[�o������q�0����h%��a~�~��j#%~�z�Hg�@@^�7��J�@3$@I����6���H��L'F܆��]f�'���J�����$5g/P���tH�.*��`�	ʆ��2�?'_TKI�@�f!��$��Q�_h៱���Ey6�$*�z_�u���3A/#[O�"4e����r���2iQ���%�Ƞ� �Ei�5ԍQ^����/��.�x�Dp�r�>�H����� 5�F4~�Hx��������s������x��F�!�&Ⱥ�}JOWSX�q�n��q�L�2�e�0��9$&�N�<!�E2����JLN+Ղ8a���+{� �w��ͥ����D�r-�o&�h��HQet��_ص��I��"\�	��|!�	m��N}�F�A|-�+�)��"�"��p*�<����I�u,qI^�՗��O��bօ�Z
�X�@�x���{r�h����^��L�_��
+��e�ɢ+��=�l=��sb��`��z���}ӧQ������11d�����x��dT���O#hN�iw@�s�j���/y�[��b�~I��(��x�<0�ه��x�G�z5ȢhG�hĐ4h���&���#�WBǝ����G�XE�*��e-<��%^����9���߶�Y�T�ym�}	ޡ��B�O��'����R�$���R���Ea�k�$���	������,g��V � oF��_ �O�A�Ԩ�KoX�_!;�%�N��9U&d�Ռ*`�c����U-I)8\}�y��s$��~���/�(ޅ�N��8�GᜳJ�3����Ƭ���l� �n���!;Cgkd��_r���5��.j�ɂy��ǲ����7ȶ�w��ɜ����%�a� �\�umTV���:��9%h�5��h�`��O��=n�#3*�rX��"��!��@��_-���E�>�Kq��l�x�����`��]z��"5�g������@���,*6�6��Q�eH��e���I/w�m�/\IO���I8J�!�����f�@/Y���S��F� ��h���<�s�-�y�>�)��	<�b�Ќx�^gj%/T�v����h���Px��L���'�GŠ�(3�%���+�������*�1�C�h�t�,6"�-��H6��6��.'�7a_�t.���p)v?��3�;lac�(�Q�8[%R��r��|�r�Q�4��/�4ζi�`����d"�3n�(b֮;{���d~)S�Y?�LE]�ǭ�=��z�!Wҥ�nm|�r�d=N�'͊�c~�S#��G6���6�w*R+�oX��g��!�R�|6òn�T��._(�=�iȖ�e��&j]��7��,Sz�r}=�靜v+�2X�u��R-7_�(�e�nZ+�B�@	L�o���]T
�3��T)�ܗ�h��Ķ�v����ۍY����V�����~��F�I{Q�&o`�07�W���#rI�8y��	 ������(E�h�"S�8P����$l��,�2PKݥ�>�i!隁�&r�c�#�Iw]��6��	X�Mr�PRȈ�*����3�F�.�i$C�$���(iǯ�%¡��pJs����k[��F��¡���F1<�N���vm8�����]Y#fШrܥ���Qı^d���#-r�vW���"ڱV��T����K��!���׵����~@s��AfP��h(L�U��_�WQP���:xí)N�<Wy�S�
%���mZ6u��7���M��W���քc��T�9�a��ڮ[�������áT�z:fGz�ǌy3�Z�[����E��>E[Gوh9f����<�U{_a�KӺZ�߷���tG���`g+�p\�9xP��Բ�����l�JH�N�;׿����$��1��Jv�x_��hD��Y���u���W]�??�!�q��̎��a�c|[���D�5���l1�'��n��(��õR�`���!j6��!uo��pV(�v��s�p��"4-�Ev[� 0��r�W�64��Ca�����$����H��c������#�dx�`A���4��,|��kj�{*�_3�E��	�VF�D�1�f5$_6 �-�P����MGt��G��3vC���[޼|���
n�7�P�p�Z45�z�ɪk�>^����*�J#�
(
�A�;�Zl�Ƅ�}dHAC쵪w�����e�u�;��ڷ;v�?��DB�ȅ٣����5�3W���gi����q�5.�������K��@!�y����S$!�r�U�!�?%�>�CE |��S�<���gd;���@dx�}�Nl�I�G�~ǜX`�"9M!��M����j�7;}[����Jl@�E�~z^r���/�$��+����^-�Fom�(7�d�W���v�>��dP֙��c�(�/ޒ��%��F8�9��0��N��q���r\(���J������� pnLk��7�����A��10��E��|�v�	_^�iՔ��C0�m�DB!��Jwe�✯��F�vh�˝���"J$��41f�>�#w<M���j���4?�v{��m���<*�V��	 ��j=�����j���1����v��������[��y����9��U`��a�[�.��[w��/ �%X��$5aE�_�#�J�@��Nb�Q�/��q?SJ7�}�LI�,i,��_r���Ԙf�)}X\�+7;Y�b�hnf0��5Y��13�&���$%�B������)�g� I�&�#2H�,�R?�T���
$����7j�l��~�W�No��wI�g��\ ��
�H~���U��%hI�Zx�#&�a�v]��eLo��)�B4D0�u�6��~�Ʋҭ���5Bs��'B�<�VS�'���}��^΍��}�&��}��o������ŪFn�#��N���M�r"\��w-�Tq(8�s�D���w��iUCmp������f��G��pQ��Z��/�k-���4�1���&r��1�^�:��6���aO����Cm�mͶ�`1����$�Z#�X���u�c/��S�&�1��{P�\?��{�� �6G\_��u�G轈�;�����&��m��D7�A9bC�J� ?^��Z��`p]HS�����eXr�ŀkV��#�,.��.��h�T������`��Yc��S�Į�O̐�zD���KLaVCnh�7�6e߂�+~qC�<�o�ȁTa��8C�(y0�r{�!�}�&<��1l����7� ��|��\�@jc�)� H�(�
������{�L{��8[�.�C���(5�D�̹*5��	�e��@�y:O̟35�Qo�Z�ߘ�\��aF7+m�$y��� 5"�t�b�]�bh	�d�/Z�ȭ+������p��&hmWG���c����f_�1�5#�y�*���iZ�\��l7\=6:=x}P)��42���o�d����6�-�5|�27�^Fhd�
�8�?5k��/0���%�!AyV��{�D&��[ta;a[�w��&����Q�K[�@S���A	�Z�~��#���r��:"���P�*$�;�E�_�j=��|�P��&�7�_�ψ���
Pw��4	'�EF�/���V��FFa'[������,W-�K�H�Q�L@��_������v~�f���1��.�>�r�c�+�kQ�y#{�O�/W��|U0N^��ߝ�Z����P�nڼ�����	�iq{M*r�bj�f��j��W�m~e�f����
Oڏ ����u��Q�#f:ټ8�G8���OH(�񈃓⽊�e秛������� �,�(��ɺ�Q�9M�����ә��1�(jрM�6��+�ȈL��E���Wc����p�!py�*O���ȕ���h�����|��`,�3Nf8\�4k�dߏJ=$�;y ����#EQ^�t=�"��E�� ��@0����o
�-���̫N��嫣��S�m�p�wF���T�Vc=���0��v�_��c4ރ��t�5��Y/)�w��q�H�bi�7;���5B��i�2�M��`W�+L�/eYD�V%Mbt���Uˬ�3�r.��m{��\�\IYIf�:G�4�m4��F��G�χ�~��OЋ<��`�4�	ݤ�/�+j�a��zK�s���q �g�F}��i��`R��;{:d%�$�O��6?��/x`�꛳�J(a�۲[q'|�ԣ��Uð\��@1fu%�>bh�@l+�^V��뚥���`��2ڶT���C�5׸�护(�ġ��!>��]�%L0a���T�15��T���v�_��2���I�A�|��ySĿh7	O4Iϴ��I<�bv$n���a��i�'�@tL�;���ࡧDN�����{>��d��&ꤔ=��_�F�A�f��*-�!��%1佷"�͜T�F3�^�탬���"�^5u�rc�aS���ok��(��C%��n��~�3pyl]�*\jr6�Mۯ�);+v� �wf	>e귃Q�d.@ڕΥ�Ah8���B0UI��Vyڸpk��7�sj��]Nq�Uy����ap�n�t� �U�HX"�ΐ�l�����ϒ\ �X=���[Rµ3����rQ��KT� �@��nb���1.L�0AF�� �șo�W�_��Eϑ�
X謢/�����c����(�ː����zGnv�ޡ�OL����8����w��~�<[�W��_��|�L����<ʉx�X�XF���9��L�S3R��=�%*�g��DyK��o"M5u�/Li�o��_B�����4I����b����37�F�EHF)�8a�a�;߿8*�ɨ(�_�?.-QK��G����" ��`���5uw�΂�0Ҳ���ڠ�0ͱ�ze&ѷ���6o�g*�w �VL�>f�Ƣ���+�rx^���G+y%�ޭ&�@0u���-|��R�H_ܪ/���@&�jw	i���58"
�~0 /La�饛���}��U�)�G/��T<�e����^����H��z�	���P���|v��!gQ�j���窰181��a[%~�s�
p9�s+�Z�?�+�
�9����g�^I͙�� �
=k0�ӗ��,ґ�J���E	�! �)���(�ſByx�/��r�b	�Y��$�vuW�[�!�8���G��I�>�����@e���`'�yh�q��|�O-ʬkH��f��.6�;�`̽�Z�\k�7-�?�b�6��K'n�9���_��`����6�V���x}�y`0"9�nx�W}�q5M9O��mFۿ6��҇�Q���0�T;F���Ϻ�cj�l�B�����IB�z�L�q�X�Y|�N�GN�9�.5Ɣ+��;�q�'N��݋/��w@��V�i[m�&A�"x�FN���ʑ%%��#�k�2��ؐ��	��������w����푇�cz��fN�_�@Ư�I�R���w�ՃG�K�o9���k	�8�йE�� ��~��bHAR�1~���U���c$\y�J4�mt 3Y�o/��6k=4�n°5u��)v��tl�۷U�����Q��GPq�������~샺2F�$�ǩY% U�WfD�
�K1E�=V�:����,��M[8-ۯ��M�A�[�g ���9-n��>&B�9�ܧ�ͮ�{,*��J���F3���w������o���Ti����&�9������=�e�2�,*��*��h_�@��(zz�����"'u �y�kh�|)���;�|�����7��|^ɒ�MDUO�ٌgQ*�)�qQ"�8?Y���o;l8�C���ޚ{R�w���N2��\��a`�Ђ�Y�*����/@`�`�F���33AS�-�w��\e�>;����[���G�C���N�'P�`��O�k�4�;y��&�����%�遟�@ ���Q���IҴU)��z˩��ѮkCtl�]
J��\�V�Hw~퇈1��@:z�N��K�T�Hݲp���28����q��(� N�ͭ��BlJO5r������,���s�<Tߚ�����ﻴː�s��D��aH��7#���;�%H ���f��w-b�O�J��hM=����o���/��3����m������=�h��Q,f��@�<u�xv:��b���k�\����
dD� ��cͼ�%f�����Znw]k�S�Vg��0�#l=>� K��
�2Oe �y���j��d���A�yd��j&<i���m�G.Hb��KW��/[Q����~�LUQD0�պ��O4DS��S� 4��m�tQ��:2[z��~و]��B���3��i��(Z�N��v����	�&5E�nC�4}�a��f�T�1�xh �ܸ�
�s��D�8�����9�v;�u9O�*�^�"?�;�r�p#F�O��$3=N�~;ݓ�^��q���h'<_ǃw�}P�� �p���@�C��¦>b�G3�1�N>�`^ge�[�t�ѕ�G.�x������B��Ak�G��pI�'D�ɭN�� ������$�� �!�_��;�&�,��ҩ��6 i�x��J\UvCǯ=��z���	?L�G���Y����#^
c�]�e��;˷PҮ�/ �ͮ���_�@�_�b�e-�3�V��M�D˝g�J&;������k�YQG���ݐ�F�xU'�Y�0�ZȵA�Kh��L߉�_��|:���0��u�.~I"���!'h|�!��V/�y�a�
DM�`AY�\�2dr��f)�B�5s��17��"�Ao�Z{>�=�S&'T��q]�K��3�'��k��ص1�F$,�פ�vbIN�*�Qz�J��~z�Q4$��DA4.�]GM��h��i���	2Q�6��� ���N�0�́m���bP�>y���
�W0r®�5K�:�b��
���7s���KE,�x�{����=�q�(�s63f\~�^��Ptb�W�塌�sk+vc1�y����Uc��?`�q�ȃd(o�BҞ1A���F-�-�j.f�=���w��!ռ5T{�2+�kn�0m�Ԥ}��	y���@UtO\�羽�#����/Pq2m���U��mÏ��p�x/`ƀ�D1�oD/��L�O�K��`d�'C]G��$w�mA��@ ��ɺ0��_N��<���LUZ�T�.l��%�.s�Fhe&z���f� �V��UI(��4J�o-Tnr���"s�ɿY�m��c��Jz�����H'>�0ۄ*3��Ih��o�����x]*&�?� ȷZ��/�ŧxӎ1�)������9r��I��}��T�0BaI��G�����V�вK����"3�Z![!��c�����~1K.ř�d���\�$u�������6}�¾�
q~�X����C�*sX�祎?v;mJ;� J��Q9ݐ�5��3�	���œ���e�tT͵h%��w�/-u�ޭ��`�1�$j|��M�Ny	ڏ�+�J�ir�9�Mr�D)�#%[��F�qB�JEH<N�N@|^]6?�C���'���EPKv�)���j:H��/���Āc�=��_�s-;5#�~Ǽ|����tY���|Y�;�� �f�0j�+9�ɻ���Ԯ
O��M�\RN��[fd8��A��ݺ��cr���J
SkI�e*�i�y��s̘J��[8��t�2���q�+K�H�)�" ���/#��҅�r��;Kqr$����I�~��G6�$v�|�!��К+N���^��A:� �["l�\e0�Us_`���xJ%����:�V�������~f@ˉ�<IKG� }����:uآ�SQ�J�w�v�0���m���&sk������.���̈́�9Q�L��XO��5��P�\�t�/=�����LhnK��x�^�I�����]rW�̟��)��hWt	��ca�Į�b5
8R�C���h�*�&�� |��;�t�8^Z�����$D�|w�t����ݫ(�����#j�F\U1u��u����E"�p�K��K�����rr����E�5�䃧� �����?�M<�m�����5U���sH48V�x�%�b^a&5_�M�Y\��f���c����?	�DZC_���� �I~��&(G�����7��n����;��+���a�a��.�u(�؏�J ��2+�x�qw,�!X��В�s��z?Ԁ�4q�*�I?����2H�nMhݗN�:�E&��w���mr���Z�z��P�J{E�y{Q�ҫ�LG�:J�bͿ�_���Wb���Y�Ob���4�T?�2�+L�g�(PE}|�|G4�t%�������^yzM��Piar�Ȫ��N�u|&��	��"=�����{��+��a��t��T:4	im�K+6i/����!*� ���(��L�^�vI	���v���򱾈��ZB���+"�o/OAUؒ7���VH$C$~z�0��U�ʋ�RBY�y��k�g����6����|��P0a8"�h�W�c��[��D$����Z]DR������4C�F<ƹ ��@���?e�֨&�ڽ���:F�#�k89T��V��l�� U+�;Eư�CJY�,�cP��j0U�VO&�ڂ��Xz�B�e���$G�u�}���I�,f���=JA��c'�N�����j#ï�D9��b�{�p�Xn���~��Q�Q��7ΐ  ;�iY�Q�W���\x7"�'8�k�j���*Æ�gꩋ4��8�<$���)�I��^�Y�ge�J�Z�{������ewQ|�M3�$��+�8��\���p#���X��D��>��˖O����#�7�R��[;��}����nE��e�2��Nl����>:��L	��%+����גm�j��V�u
��:S������^Q^q�L�F�6�E�)Hd��������v���o�QnVˬV�����	��JZ��0�78�?tH�����K���"g��Y�� X�x4���$��`l�0a$��+h���x�U���=1;��7�7.�~�F�V]�����°��ꌡ<ɮj"���s�/��S:��ڥD��D���Ò�#JHs���CG̼�uzK>�w�9��uV{�[\tr=hf����2H�Hcl�TL�R17��q����#�Hs;�KW�� ���K�����,��:�O!���D5䊑�r�$��5��LD�$<���O>A��c=ֆ���@�~s��Zϕ�F|.��J��L�Y �;4Ld�|U����IkU��@9���h�&FYQ�����c��1�jd��b��W�����?��v��$�5���m-ީ[p-u�
OS,�ɗ�@���/�h<�>�'���i�B�O���
"�[�ng����θ��E-�Nɠfð՝3v@	>���]E�b;@ɨ�����^��c%~{��FH�@�u�Tc�3!��(� N�^�t�zO"�z̚������uT 1?�ͱ�r-^T��E�$��gJ�l�%A3V(��q��pg����.w�͘�����v��[��0��&�W��P��[�t��qY�����h�QΘ]�5��<q�����������+41nj�]�o�357��A�KI�m+S1+���L7�;��տ���F;��w
��y�R�J�kw����,�^[�X���횼F� ��4�����$xH?�2'���(���k�8V�Y��-Ǹ��e�W����,��fD�s�M���ôғ����q�H ��Q��_K����ݟ����L�^�����z@b�zV�����G��J�NhbT�+i�����3l�@?� ��:@S�]q�lOQ�8�E;2;nǸs&���N��g鮥#��ܑ��1�P�0�~C.�oPV�V�A�zU$����="��`��&���'莺XU`!�!:ū�q�C��݋yoY�*��?+Q5��![����4�%.`6?#����a�	�<Qrm��E���j�vd�|��!��9�K�S69?/_��Je���ǻ���ڳF�A���^M����|m�s�!�;���=h��~��y��!�uKg���݌�13al�ӄe��x���D?�^x��p���.���U�_'�E�&�f�c�!�
7����Qބ�z扇��
T:�(�����{���}e���K�)?�HN��kѿ�	-\���ױH9h\��@Y���{�F �@�S���,�v0}S� ���z��-Y19���6�|���z+zܿ�٭�+��،M�����>��������|�U�����׽t����T�.�.O*����Vo��-�r�n�.r~?dJV�\���[�/�|���ʊP���)��J��g�Y0~6�(q��ƚ���W$I�=ʹQ�=2K�8&J#����u��H��Sì1�Ҭ���E]��k!�Up��Cz�KT���yo	[� /�M�V��fѠ��r(��VT�!���/�ŬL�jx):'5��P}T�y=��'l˷�m$�����{~�kkD���i+im%'�a�5+� �!f!��bu ������e}(�L�x�LsP���!�ρ}�|/v�Il�� ��h�����#�75�%�C\��@"Nc�x!�FM��U@Dw.��^��l!��6F�_ҩ8,���55fmT"J �Զ?X�lou_a�L�)�Wg�"QO+���i�=\���^��K��L�8
��,3k����aRHy��$Lf���'�ς@Y)�NH���m2i�!y1M-��9Sq��`�v���r��h�*�X�.;ٟ�����r�OL3�q��)4�Bƻ������R	�J�:�c�}�!�9SV#�ʖi��ŒH���o�?�k��)�ے�y��4}s +p�E ��
�� ��J��æ����)�aht��懥���O��]��t�\A�ˈ��;췮>\����ue���{�n[���tF���g2�pI��7MT�'��"����[���sE88tk�ST+�1�����5��+�6�5������Jz�<2�ݿۘK�\�����ќ�������b&8��Zi��;����5�ԊԴ|a�/��[��~���K��2~������ D|I,��p�3���l%��ݖM)�|��4qn�̑Y��������52wp��dx誷�}��%����쪟���-XϷ��{R�S��H�����7��{��ْ�Jr����!�i�W���l��YB�N�?m}�Di�D�"�9ķ�3�X�i��q�El�{ۉy�����5>��+b�
����[\�G�#�rV�v)�g+����	fB^Z�?����)XGVH�"("�|lI�A�V��)��f�t�~��*�l��4֓�P+)w��>Q���/*�Ψ��]4��;_�rr:�@�x �h�B���=�������K��V��R�`"4�����!�O1������M�q9������J�w�nF���JDM�'i��eο���(�8�	��J�^���Wfʄ��)&�`��ov�i�ݔ��ZO�]���3��eq�gT���{WNʼm��q��lI�A�g�4�K�s�΀ІD�֦��Y9*w�ݐ;�C]���Tъ
�,c9�����r��0��#Aב�I��'ĦG���'R�_�,����^�T�`Hj�0�:��Z<�fQ�~�E��K���V�-�R0�XJ�!�so^i$$��:K��H��n��_�&[�YI�Eԣ�Jtvk�
^(˄7���_ˀW��
���ҡ�
;��>_�O����FL)WSvu9��,c;��7&(��AM��Fd���w�ݾ?R9'�e��p�*&{�g
	�6�4MtǑ;9�d��5�\:WUm������WS~8��d���q�v��mW����n�'l�]� 1(����X<��0���[�����~�\jz$�>F�����h͉�k��}�I���!�lo�8r����9jYkw�#�U?�[T��vx{���jT�2Ű�)8�u��W�H��
�bW߿�,����l��ی�IG����;�хP���o��ڳ��w�ZJaW?db�8�p%�vW����9�G�~�PAڮ\����@�D�6Q�97�W�}�a"�k}~㐨Q"��$��9�=
W'ӧYR$oXζ��G��@���6M������\��H19Usqw�3#�y4�D+���hPF4��PT�	崄�IFR���on�޴�ݦ�$�^Jj��0�@�5t��(���᡽����}�ۂB�	�{�X����*�e=�c��3!)�pe���'��N�0���y;���_B[��I�[fC�8��ZɄm� �w�r,w�hYsJ(�ܘ��������\��ќޗ�Ŗ�,7y��%����{�g]�X����5�u�w]��6��ޜBz�Ҋ7ث�R@�m1�i SW���$(Z�'X_
vy��Q�ǡ!���+V�YB�����LoX�RA��j
��XE�p[S���Qm����۪\�-������oh�5����0xa������$����߲dz�!s%M�Nˁ���H��"�2V�YC1)��X�ɫ��s�#�gT�ed?�����>=M�@���(�7	���}_����Ca�gg��f����t2�!���;(żJ�o�S|+�I��@*�Oz�2��E&�w!P�d�:�~ʊ��pDmv]�>O�3i��`,ɉ�����h��c9O���o[yU'1Qw@�,@k����(���tڥ���ڶT*�-d�pT�B�(�k^?��t��+2��M��?ӗ����v��(�"s� �%�#�~jHv�>�,Dw��ID��r��A�?��ld��:��=$q��4e�}�o�`����'�Ԯf��~���< �J�=��ްtY)gy;�\��Q�I ���E�i���"�y�	��]�}$��O��e;Z>���L8
G������J\�P�'��YiQ��1��� ��T{�D|ɬ����Đ���c�LQ�*:@��k�MYY)˿��f��1�Z���jR�2��lC�"���n�w`aH�y'4�@q����t���5�	D��P���Aj��P��k\�C씌�Z�D����Ę+Hڥh��������{��#HcIP6�1I�]��<��ä��`���oKB>4	��D�K_��ӛa<��颤w~�G�Θ���6�*��d�du��,�5<kzҋ˭�;?=f�-��l�`��L��Aޫ�ȱR�JhqJ����r�9tjK���qQIAG! �{O�}T��S̬(q+W��(�?_t|�j��CXn?ิ�X<������i�ԡ�6M��|�|���}w�.�)b���5�_���U��^�˚�O4Y2M��;ߏ*3)�6���iòw�3�͉s� U]��M��޿�a�G%wd}<p�{�W1@�3O�HI����T�r}����l1DA���i�#p����X��ަk�a\n�P�\��U)���o ֟1�$��K�� �!�8�tԔZ�#��b���YȺy�&��1/�����l��e?��,[\�
U����aA��՗����,YcC���b����n	�pu\�z)ҧ��)e��\��Ld��Q˔�f��:�M������QYCu����)�� �1��h���4dkfN2�	���'�:�Rf��@�xĚ�=��w���%�ÖU"֍$��h?�ёWJ:�A�/�B��c3=H⁤vv�J�*
w|)�X#``��V�""�Ek~i�I�I�M|���IT��P���ǜ�U�*K����b:��Yz�W���x=�Vg�es����ɠݍ緲<Cwk8,U=ɤ?Rkx��K�wA�3��MG�΀��;lV�:�Z(��w\��r�_���廠}q��En���9-���j��r�WJ�������_���Gk��UG�Y���±�R��̎t%�i �u]s�^��m�4���\��O(���
�dLe�#qA�i�x�O�:��}g�<�Ov�ɡ��V�n�[�0NM��k�r~- �"S~���Ri0/��%�����s1M҈�L5�,�O�rAM���l>$�l���(��� 8�pš�4
I%+}(ոߏwZ��sO�f%�����ڼQM�_��I�b�[�����z����%�TǪ5�\�J�����z ���[�"�$�ӽ>�`��cx��y�����bu�,-���<5UL�:�d�e�x�$�����&W���DX���%6�b�-�wgw����|�3Nx��ZXìi+� $sos�w����`[�?<��W�2�\y����1�*���lP�Q�J"�K�!��O�t�#��W�6�\��˅���Z�L:�7�g�mg�5��,8��[� ΅���E�͗' O�	3�Pώ@aL�x�!g�,��z�gȇ�(�yb�`+��z��,�>MS��� H+��k͐�잾V��1T�Avm��#�ʭ#(d��T��Е�������n�j�1��,ǷEu8c�r�t�-�����L/�Ș���\W�������@�}��?�Vˉ�Pu���g9.����={5�=Y���&]�h�9:����w����k�)��	��q��ۺ{�:�DI��s��&8n�#x��aȥ�X��M8'�$l�h���C�(�t�Q�8	Byة,��Yj |��3�'-�&���;*��O
T��ٝ(B�.������¹�6'�1�rI(E"�wb3� �0a�J�M���7��d�k��Z79�Ú��"S��ZR#�g9��+ǌ�ދ%4�x�n��Y'_��_J�٭�L�����u$&����f�������&��DB6Ɔ|���7N3��0哹~�����J���_�s���&\�Mm���Լ�r=�e}���B��.���O ��=������xx'�TsJF��t�C^�O͔j����?#�x!�=�q;Pf^(ޱ1-:�
�Q�wi�8	T-w�q�%ǥ�'�Ә�/�zG����[TJ�I���hݨ�&[�����9z?�����ʬ��R��I���q�b>p0�B�C��d�H笎�e��G�8RtZr��gO�3��&����"�;1�y��?�����tI�:ZRG��$=`��L�
�K?x^8�F�N��}�f�Y�V�ߋ'B���z��u��	���Pv�����mG���aP�/e�w�������Hg��AyT���v{]='��u��R��H�{N����;�V��!�GzZ<�j�n�OnU?�^�waN��@F](��ȇ�U��hT��j�[��n�UHKm�BCG9�,*�6h��jpҙ�����"�r�7��y����W�J��+����L�	e4ze������q�\�:3���a~:��U3'Е�N�-
%��	��*�����HA�P���j���z/O�$�՚�儷�v�� v5'Js�w����}����B���U#�+N�M�W��{@Q���ҋ�_���
�;~�j�%k~���#�R� �)���3�*$(h�#`�~awZ!:Eb�h�@�N���NA��֫K���]'N�p{H�@9*�t�����n�a�{��?����a=
�J9`b�^�k�Ҽ-��چ5�e�u)n,Zdua>{������J�׋+W��M�hU���
��+ժgo���ƚH��{���&�e|�Za�E6���)�;���ȋ.�~L�_�g��>���N̘��%�Z����T�4 � �p�(Ñ��0.Q�&J��*o�(�6T��-�+#@�pj���0��n�쓔+t=�>-J�����T��B1VL���Qi��:�_���ǔ/]t�>jpX5-#�v;e�]R����.!�h�Ϛ߹|z�A9ɧ���\Ґ�?r����-.@��8��h8����\3u��65Hd�?3����<EL�0:�՘�_��m��!��O"I��l�V�wG�����$�wae�{�~j�d��eP�:���(����N�l�6;	���W�DR�m�e=L�jw�VT�f����eǀ�12�K8
g��]���1���YY�!�s���)���^ڐX�a��bs����j�?U��	ucS�97�aDH��u~��u����?�E\v,�?��y"Rg&�o4���^�k ��/K����X~�[6�f4��UØ:*�)Ws!�Ob��L)6�`i6��Y͹������Q�iE`�2.�?&���Lp1��c�J����ǵd�E�����Pz!��"&��ȷI�m޺7�@�R����m{����o%?�Si&�pZjKzR�g/���u0I?-W[P�L5&���fʷ�OK�7��a�B� �p�	U�M�a��p330�꣤��w�����4�}j�J4�	�U ����.�A�q �bu�ܘ���J>�o�߲�a�*�H�_!�;g0�k�N�~��|����ğ�T:'/	����}ʈ�zK�a���myc킱����V�%�œ�=Ɋ�М��x�~q��W]�,~�K�_��l-B�Ǐ:J�%ho��|��{�N� ����b�4��ɍ!�	�w�O�F��  �+4ׇ�e�°i^*�G���<�	���W������l��ݙ�2�2�	�6QyrP��r dKtc茁��w�w��V�r�B4�a�������^=Zޑ=F����SP�=U.)?ۻm�t��0���L�
�p�t:�kZtd1�"�>j��>��)'��
�K��F2���x�>�����C�<Y�HBp�G�R��58�҅�G��>�U�eu.`�S��w��$�ð�����`��jL�Y(�_ʫ4���ɲ�'	��Bjt����K����bX.3a�T#@_�y�P=�w���QSL�ҜS&%.�RR8�?��w| �S(t|CŸS��繗��y 5����9���=�_1��cc�Uf7u� �Jj��	��O)���'��.8���)t~k݀�?X�_p�h<�ҭ�M��n�`����淋��hu����ȗ�[2�\���1�&n��8�,(P(�9��̭d�nɪV�0�i�Y�J��b^�p`R��¬�����zL��.��X%B�T�5_�ϔ&��:����`��H G�>۝�o��?�^qC̫�h�5��	��/�Iv"'wR���,�����Zu��H�a�'�/a�a������/eہU[ɅD���:Qz����Ŋ\���¡�+ě��hS@@Ia�{��Վ֞GT�==���e�F�L�|���Lt�ę}@h���t>�N,kS2K��7V���B{�S�Y�MM`Z�T�x����p"2�?�I�;�r�|7�5����N��d��&6erE�&N����e�rx�Uv�`(Nᗓ�o�j�o���.֑t�T��2Ќ��Bƫ�'%���ag�(�����[b�*�d����ܪVwK�γ�R)�a�/x+�==�Gn-K��b���!ŷ���j��E���uH�~}T@b�>fp�^{Q��Y���Y�	�A�ఔ�{�P��d� �.A�T��W)��3<���eH��jhfSJd����C��\NaW���l>�����X�m�u޽4KȖT�=l`�C�R;IL�3o�tƣ~[tu�u��N�R��Ż>~L3Z�r>~j��d,p���C �G+���^j*Ks���/���7�б��F����f�������́�~m���$�(MU�Pޑj�/q���,��-�לW,k�ή�P�{�.�C\���I8�D9<�����<�ɒ�����9��9��y�ߌ��2������T�?�����k�)T,#�Q`���E!�d�Z�[沕0G�c��G�f���bnH��@k��uG����܉D~�8pY<ߛ���&���