��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��@\�r��5#�\G�6��j�@,�j�k*_n_C#���,��(��?G��f���:�����oR�{�c�X�dˆ��۰��\��췬-��0�A�0v�.�̍��B�́A5�A��J<De)k�+�o�,Ww�>�K�/B�"/�G��`��9������1|�>^z��%X��c �+/L���O*P*dB%䱖"�=a�I�>t��-Kzl�����Q��a�`gް+?�\�<�����q���p��wWH�q����\��c�ģ���*���#�T����ݑ:�ػԥ�m���]E�l�L�=ݶ��Nw�/$�J$wu-�#c���,�5�&9p��vrMx���`J;kf:�ƺC9�B��!C�Uk�p��B��d��Kds+
?�'g� _okA��5"�.53K+f�S�^z1��?ˏ@^'��Cя�#��J�Jc�~�*.�6G�H�%T-��OfJ�]Q��/}L���"-�'[DW�����y)�;��>Ȧ1t�bV
��}4�%y��*}�B�_�s�5��AQ��H��ν��ա��d�kL��5��ƀb(�YIf�O�I����e1^/|[�9h���!�r'9l���%���rSbeg���5T����F���=W�a+I��ZJ�.P��rO�朳�`f�������8Y�y�i��iF.D�)��8T���]����{u��cl��/Ly6�����U��aP�3�ܞFHØ\�� <n��o�8Hi���Y�	ć���e���(J8-����A�M�	 N����j�8k�:<�^��	�z�`���%z�"qǋ\rc\b�V�R �=�����
�v�B*g=��Ҽ�	\�����A22q��7H����s�8��3ؔk�T�͟�t�.p��81�S�Re�x`Y̶ۆ���j+m�ů���TEl��(�e[%i�h(�C���ꭀ�O�C��ѓԋF��=+v3�[�:������sBv�JaU$b6*t�m�%��Q߫'����e/D���e&6h�$��?>����G��]xZk��~9�48� �]���n���bu��(��x�/���R�R�/׊/����f�y,f��F�(�!Qi��2���p	�$\0�E�]�?~ه�r�A����R�7���Ex�ڶ�&��@hOO���ٴ'��y����>���܋��i�C5K��}8��/B 򤲚$�P�{�I$f������.����\����h.7H�{T���q�w�����,o>����� �Z�2G� �0a{3�va¶-pt>��/A�M���e���N�1I��:�`j�F\�!����n[�0�ks�W� ��7��:�W���^�R���c�eY��Hf��̕QH/�U�(�.���^���^)��@�{#,��a^��ԅg9<!�+�#I��#��h�P�1�#&���F�����e$Ǐ�:�0'-0��������*�]Dwl�1�c�ƑU{�#)E��;�6�Үgjө�[B̫c�A;����ygXC��:i��,0_̌Ci)�H��C���h��(a��{���(��D��&�H����+GSU(������]�]
oH�*>+c�Cf� |QL�5��Q�v�.gK�|O� ��}��mkW��KU*�%.�ga�	O�?83�EM�E�~�?KK�:��h�!Yp�'�W��6nS!~b�S�BK�b�se?(�N?���W��0�<�0IP��:�+_�w��P������찳����9�[�$[�Ř�X���#�� v'�/jFWщ/�i	�:7��O����usނ�љ�B�e�p뵺j;R�v���Ԛ����,����4�D��4Vq���G��t�{���?�Yí�}X�#5��f��Dm2�I�k�C;��f�ӄ���00t��(d��L� PŤW� �@�Ļ���+���u�?2��O�� OCZ�?�l�������غ�A����E1W���7Sv�lŒ�Z�!�Gt��0Yl���y���$�Z�m�	}�C�f�s����{~97�L�<�`r�Z�<�9�QU�j�{^�]�}K�|y�kdNġ�Kz��*a�>��C�ϲ�=B4(c���B�ǒ5�@����)���/q�٤2��7 �&K{3F��m��ZuV�j}=�\rH��G�r�L���ö�b�P&�K�SR����48�UH�K.� Mt���c�=y	^��?����b�<Uu���	a����Ћo?���$�o]`�E��vy��U`7�p���kDF�����%A솂e	][n�a��QKFV����;�!In���_X?_$��3�[���M��LU|����c�q@�_�J��yb�n�/4��>�
�@�Ƴf	v�"L ���m��B����,����Ou�Z��	�E<� ��R�{�y[��MH��L����d����b��V`rJ��<�k��'�� �/��QR�@�uǸ��C�D����f����tuA���Y,j�� f4�����!@�v�l1˴��rfq�vb�ƊD��Wԗ��n^��"�d��E�D�P6�'��n]�ݳ��|w~�PA�V#0_+����q�F*[�� �	�n�1���w:t$����	�/�L@��u����p�]8P<������C�E0k4�0Q5�������q����x]RBٳ�\�.A�>� W�)X�'T�2~�b��N�󽴖-���/��yn7�zl�Z$hA�T��L����Y�W�z}g��!]^�yy���x�"��Ps�.���ř|�b�2�?+H�=y�H_����Ŗ{[���񘌞'h��:F�A���ɾ"�2�Wl�4P}�q_0FY2�����Q�)w�8<�[��lMC��׭6 ���*�&r/��j�����{�d��46�A����KW"�q��0���,�g"s���֚��A?oA��(9q���|j��Q�JR�r:��Ф���av tf����ī�&/aE�	���K�����i����t�*2w�(�n&V:��a
d�J�e`���9����$�$0@5�=V�����9g�����gƐ�Řj� J�,�<ok�i�$s���a���Q������Uh�j�(��*&SA�>����[{T�WJ�SԊ���j"����3�r� ���Aa��U�x����b�2~�*�]*�¡W۸�Vy|�Ȅ#3���ْEu:G~>\ˆ���]�e�;��G̼x��yjP�*�:��NoF+{M�Zw��k�"�DEدV�+>�"��(�V\(X�� �͎t��|�Z�}�j��#kl�Y� ����]��xuL�~�_tz��(y�Z�:����R<%w�2�从&���,��m�%c&�I�(g�0lrRީG�K|��L�\xH����v-:��T���kg��2ȿs3t�Đ6<_��TN�1����&V�W��K���S��&�n�:C75b�T�8'�J��o l���g�t���dxk�Ѓ��Y��U�D�G���7�Ʌ�v3���^��<�psi.B1.�P^��8$��2 �B�����r~�3��G"ӊE�:�w�7��
b��To;�j���7��Nx�����L;;�&�Κ�:���R��}�]I�L�;uS�L��9����l*�A��)M:7F�
?}'�-^	��b��p��A]p�q���� {V�Y������ +���S��	hR	U�d�zz�Y����Q���B�5OK b�a��`�5Y"�����G�6�X��!��w��sG�N����|b�aN�w�9��Nc�ʠ�>=p��p*�ģ<�����M*��A࿕�`8S��K��S����W���%�x�-�K�����2~�p�f9��S�I�4�a�!�V8V>Y�ѹ���S����+A�����⠨������?��>�e9��Ce��C�.�7�s=���K�~�ZFQ�����+�b$��P�J�5���Y������v��5�>%��w��qt>�mM�8�gb�[z����>��Ϣ�,z&�����4�{�L8�ȶ؝k�=�|(�(�mͪ�e�̷Λi}�Z����V쏽������O�����$~���hG .��d'�TuYw4데�e*D�
�W:�]a`�֫\�W�i���V'k��{��O�Q��g�o叔Fl�hv�"_�!��Y]���N���T�������8����86�&&C�"(��\JV�ذc�oa��E��хX��$���_�>��c���H��^d{Gc�ô�#�*Ay��cO��d�'�c�Mϓp�h�~d��|��),�aB����s��z��e�&l��B<��� ���XD�Ho��eE��A�Hz�n�m��ˡD$'\Ա`��f�w����¢v؈x�w�V_�.�B�%zs\'��m<"����~��r�댺�'��?(�kQ�2gXڒ��9�^�P�:P#Ռ��z]ʋ�	�	ey�)���	L���UAzr���FR���Y�oC�G�'��ɚw�������h�{,���v,�}���|,D�m��4U�6�)�9f�e,iWY�MsI�}��YSS��1w�쌡���X>g��2s[Ɨ��z�l3�t�:ő�1�Ü���6^(T�p-�YU˝q���ĊC�3���������3�Dx�z'=7y��oV��n%��C��t|y'��w�s�8Xu�&T5��ָ��؁���C�D������l����'fr�x<x_�I ��8�� ��vO��y�i�n2��^oy0��i�)�z�cL���_1\��]-�xF��5D�Ҩ���u����C��l�oL�u������+�	�^*��ï�bJB�������� �A��q�f�b�K��7@T���
T9�㻏�!`����'rZ.:y l\1�
O{�$G<�FM���h�����[8���`4e�d�#�,����{5�.l��>��؎^�5���0!�!�Q�j8��x�8����2��s��j�Þ��i�_hB�oS�N�j�댠#�'.4�2�u8��NW��[� +�L?I7B�9r����yO��w;`&-V��$�I=�V���O?^�M'�J~�]������*�!v��~S9�=�����8,�g��dT�G����sv����ɩhos�:�jz�ز|\�t
3w�XV��ܓ��W�>����K��������xwkO��T*^�>����ZV����z:5�ʱ�*�ۚ:s�V[!�A$&j���J��
$=�ؐP� FF�]�*���A���G�$�۰�q��ֿ0��ۈ,.A�W���JȽ',kuC>]�_UF�8i����gjY�+�Zf�kE��ş!��� ��1�V�r|�@�!�QR��4������>쪮��p_ %�J�U�h���%D���Y�n���ð#����@Y}�3���f����B(��&�G��T�^� ���mtj�0�>^�iB�s���b�E�=�\�=r@�� k������/N}�ٶ=��P�^����K�G�(�;��D������
[�$�����Ҿ����D3�,<*���������W5���t��M���2��e�Z���)vy��p�hin~iq���aoȧ��p�����+`�.=1�QAӹ�4� S׽K��w:Ep�L���x�����]�����~�;�7@s�8# ��d�� �"�>4�۳�.�z�h��mn�u��N)����(�#yȤ�t�R>�2̇Q�4'6l�ֽT�{��#yܡ(fqQ��m*]�>��jRң���(V��U��3h��H݃,�bl�?�aC���ccg��1��Y1�^=�Z~�5��@:�s�X�4V���4�GD�66�#/��sZ$���`x;Z�
�l�\����Xݾߧ=5����y�;�tH(�k���anY��ئ��,����۫���lLԮ�����42y���?7�:$j���*35��u\�g��p0�R��a@g{-7�5Z�'�[m� G����eƍ�$�S©8��.�v�.�!E>\E���"Sp�8�� �D_CRQ�b��%>$*%�ˢ�|�e�mO�/�[J�W�{�1|p��a�G���*\�Οa9�^%��D
C��f�-��S���r��i���h̲�vA*��;���7T0���ζ��m�h����ޚ'����y͸��w����-�L�0;?:�	o6Ay��s�S��I�~������Z�_u���}���T (Kyي&u	�4���pp�/�L�M}��V�dl9�V�����J��*�63¡��b��
�v� r<��oe,��y�m�~�����*;��Uq]�v79�3�����y����b��6���J�FT�G,���v�۬n(B��*��y���'����s�h���cȋ�"���ZF���܅�C��=o�g��� �K�E����=�t��$�.�T��+��U���4�rH�����Q�6���ϭ�m��ےOvw�EƲ�
I>4)ʘf�l��Żvj�Ȫ�v�Q�5X��0P��q�P��W���*5P�v}�&`j�`�&iJe&��ܬ�czI\��5LXF���*?m��$�i�j
u�X�M�_��� ���K����T�0�>J�DW�S��-��ؕN�(K����G�#��<{��'d�"�r�Oތ�F缐4�O�HZ�S�YUk�/��ɪ�.��}꟢a�: ���@Ň�Ocާ�j��7�=%p�T
Q�*��	�y���ɟ��bLE������uTf���&{���Qkɝ�o�,�C-P"�	A�����D�+�&lS�>��tr�����k-�,���)y�Q�4���!���u��װ�%H��4���z(18°B�(�p*ڻNn�i�˒s5�!�)�0v�_'1r�T���@,��d�[��G0Jb^��-̔�#p�N�ޣ� ���O����ˊ��͹O�'>F��gG�Tks�,�r���<�x\�uc�<��Q_���E�/ڙ]9�go���^2�^e��C;�f�\��?�{2�!~�oS��_�f�}�Im�[��-_��W�y�4������T�I� �����Rg�L;脌9J_l*^:��*nL�i�U�&�R��6}y��a��˞q�"~ ��*xx�w��i�甏Tg�c�Y�7z`>RJ�~�_ �YXMb�A�Ub�%��� �0�\�m��]k�yL>�w���@���n�mbz���5�].F��x���g�a~"����B �Ϻ\*��벳�]卪���y��5��1�Fe�(�!�Cj�K���0=�����n�a��
f����a����<d�����Y�Ǐ_})M\�]9�y��ܖ��j��֟K��葊b���-�G���
��� KC����쀱�ZI_�@?fp��e�u�I&��U�<����m>��J�[��R�Y��I����nf}���Nyi2}�D���RV�6M6\
�r|KO�¨	-9]Iw�����9�qi���^���R��U�q1���0�_UB?��")_�!�w�$�(�����^������꘎�k4調�v����ZY�f�I�M@\vΛg%��\�c��6c���/��,^5*���_l��A�Te��+Ƅ�a�L��
`�O�0�ե���z0p�~��S�:B\4F�].L�������vv�yi�hr"MG��(�|!_�u�=d�v����3Y�x���&\��Ct���b�CRYA�~�?���c3$J����h3^!�E�œ!�s���P��'r�hV�}Cg��	�|�km����y��fO+Ү�6�:Q��,RA��^D���z'r�/����ؘA��>�3�V)�Gi��B��s+�4m�mJZ;',����?@�����P"��o�Wl&��(%n���O�-G�@�w����:���4 �@5���Z���О�+�	xR\���7�IL�MR_DzXuv����ic�+z�����M�(PPz�Ч�h
�o#�W��̳VI�]m*��*��o��Gzu��b�k��t*�?=���HS�V��m�GK_��^n�zXn�<��D��J8?��dӑ��	�ÚbC�
e���c�=F����*�*;^P?�ʆ	7��@�淊��p��|qⱴ\rp�0�n�Z�C�o ��wUr��:��"ZI&ѕ�l�I��z'J#����z#��0��Ԍ�~n��?_gq�d�'�Y��[R�=	Ӥ�����8��u��3�)�]<�u��X( ��X�Kx�x�qRx�q�i���A	�w+�z� b�Z��� ���OR�I ���!��$�z�41����"�1��T'���]�Q`�����k/��h"��A;����8���|���ň"6�ZD�3<̙Ӕ|����}�P�:�o>Z��%�7�*!X���HF��HW�L��Y�T�A���#���^%֎q��ʼ�����l��7B�!Ud�Y*�9T�v��8� �NH���6?@��G��IW(�+*��yZ��ud'kI;r� ��q�ߩS��}V�.w�8�d]����`��鉖xH�#n�ҡ���;Jښ0�s�ťh~C��|�>#[�Xg@RI��p����54>�Vjr9��Aף0\`Å���
 Ո�b,��tބ--�ا?�V���:F?���@�Vf�1�E ��
רV'M��%�a��-{��� �^@l ]���7���ˤeXV0�/y9)�I�����Ш��r)*��`�T�5N��XmW���Ňd9�D�ǯ�/i�ub%�6_"������<繳� ����̦��;�x~>�26�?9��u���o�ko]��f4����|��Ɍl�>L��̳Xʦa����}_$+a�S�	V(��n1kq*_�#^Vo!Y�iP�+0�"�,�'4j�pM2Y:0:��+�5q}�MY�()��7���P/<�_��̖�~�%%cc���k�&!���y���y��It=z���<�����b����qK`t!/D�U�牏��ON�M�dW%�3�I��[V�*�[C�,Ev�^���&��u��� I�/�x�n�����A��{U�)�w�� ���r�z��㠎kB=�t7����LT!��ҲV����F�s�"ٵ���<���E9.6^�*���ʰRCE�W�HuA����C'�@�;s�˅�
\cm��3~��3��`.7,�X�fD�_�`���F��t���1����w�cGV������!:�6g�&�*�z�LOh�i�}�F��4PE��F�.\��ڬ��WoHpĤ󑸛�VqCf�_�����:�Q�# ��l�n���C�"|,�N����+�`rQ|x&���iJ3�v�-��4��a5B����HZ�R���b����YP��n��oq9,k��@t�>Jo�7B4�~��BX��{�*���隹�^�;Vpɔ��Е��Z�g_���W��~�l�!scz���򹽔�4)e�k��]/vI����j��ɉX\�a�sO�	�f����X	<�P#ux(� �'J[�~-�0>#�¢:�H�_�Ս��B#=b���$�{=
�zh'��N�֐|&jw�K/֝�ɮ��dБhv�ɋ�2\�3�C�e�X������9��������j�N:Ƅ~G������.w=f�]���^�KQNNV�wy�����x�n�"��$���[��mC=�#�������E�R�6W���g���H��b.��_�S5*W8.uYY~%mv%M��6~<�����D i2��Y�Cp���o�"U�9��#�\��Ĉ&�L�}U"���CW�-���=~P��\@s4���2}B�,���'CQ��,�HX�6,����I�ԕ*���
҃���� U�IMf>o`b��u����k��Q8�}���{��� /�=W���xߣ�᧼>*�=�CP�d�~b
?�|tr����m��1"{b�p5<�UI�
�m�ʷZ����<(R8J�^�&��V�8bl̨��D0�Vn�M
l�mP�d. ~�_鬺"Z<�Z36���Y"�׾�͡AOm�C����,���,�|>�T�9�H�8Yz�xL��,�g#���W-����Y7���]�)�5�r�_=�^-Ld���,��!9`c�W�PQ��~!kD}��qV�>I�yh�l�؊gi�o2f�m�!H��8r6"�g�r��ǩ����j�i��I��`ߏDK
�#�$ǃ0���5}[���^_ ��Y�����S��L���5r�Cr�/Ǎpt �Ī�j9Ej_ M��EI��� SP�f���}yPfS�N`����s��-�W^Q�B24�HEcJ�s/5�*�͏hZ��#r\��@d5��S�1�KJ,0d�����7J�#��AU� R2���e�f�{(���{G8�N�>U��I� T~hn��E�Zsb~>of�ׅIن ���UPl�A��Aj�b�M�3��/R�nOFa ���T*�U����6a�H��"7�g F�^'��;|š���i�L�s�h���2U#�aVe0$����(�?+LB� ��qC��#%L�*� U9�7u�+&~=��m\B�"0��+�>�a��*��L�7�W\�NY��8��V&N �!���t�.#�ޣ��	Q�I���՗r�{�)��LGa2>4wT�͔8M��Ѯ���^�+:�����Õ�*��eF�5Yi�ാ��Շ��	�YD9��^�ӄ�E���u'#(e����G��O28F�@�{�zu� ���'������2~z�@VR�MĴG�y��!��sx*B*z>q�,=��3�T����f8^i���5���Ϥ��ͱ��\���/2��8q̱�z�� ��
���0\�G�A<r���q�@��ȓ�j[���\SeB*)͓WۀT����1F��z�*0���v��<�eDRl��%S��{�i�=�I���h8�>��\�s�l�"�S���Gb>uaW��6�G&�kё��D�[�B��<��K, �}�;�CZ5���펋2��F7��
��Ӣ�L��3Jm�X�<Z����ݴ)ȥ�~qh[���G���'#U��a��T�߰���v�EL�5��ՂQ�~Ն�^"my�[�XE�$�,O�٢�C�h/q�%F�e������N���q�A��g�ĤO=���m98ݙ��#z���D;$+�T���%�¦�ܛ��ī��Q}��E�A��k�g�� k��҄-��4'��$5UՃ��<�����O��p7�������y\�B�����6��	7;�u��f\�jP���\�O�]�@$>*�;%�t��u�b8�'�B����P���	ɒ� �.�e��/����JCx��4�px 0��_�Q�b	�8p��~*�Hc��E:S2Oq��`��b5���j�gg��U��u���0�ɪ��0`3��ys�c�DGf��]Qp�&�]9:�O�� �{��&���R���v龿 b][�vD�#�IN��t����>oRx����2tO6��=�5s��� ��ۋ���X�i�Ӵ�������zh�̿W�.঺ͷ�m-f "�P|Q��V�H�4Dʚ�I�0|�&�q��Q��|_�&��mɻ"12�Y���>�Yw����,9:#(�����
֝85�Ь=@~�j+�����CN�m���n5N�:�zU��}A�D�G��J��Ԋ��:y6�,-��˸�K�hPЇSI�U
�@�؅�$ŋ�11����g�}l��MZ��Nw^2�	�:1S���Y (�����C��Z���\U6ː �;?��L�d_�©�`1S�qD���#]KLE��R�Y���#�"xh$�Y@�^( ����
''��x��(�q׆Ӯ����BҴ�A�g�:��%ͣ�A��M$���e��-!D���$����:~�`���A�;.�Qߠ�쑯�ԛʽ��G�Bc����xd�ihu��\dL�����׀v��:�#��#Bȍ;��(q���r�r��گ��� H����Ӹs:׋� �]P�'2	���~'�{
����P�Ө��=0�+�����p���Ҍ�%�w����)�}����Ԕ@'��t�1I^SW�%:�'ZT83k��2�u�\��Z����<L���Bi�X3ս�'|
�Z���/�x�Λ0T?f��Ե�5�(���CX�;��h��"E8}o��^�`Z�����ȴ�P�.��I^��VV�o�/�(A����[Ά����D���B&6�=e��E��	�Z�4�kO��s
�$P�g���֝�`$>���2LuA�H��V-a&**��lö¾
8�MַZ"Y�۰�J+2D^����M�k�t͵L`%������ K�[��z�3��&N��^|[�fC�o��*�'~�<C���V�͇Y�&�A�aG ����s�U�P�T{^T��`z;��̱��I|��|"=��˴�LQ��h�)=�7��Q�ڎ���#����p�>nO��}�IW����e8RkF���	$���K��ՙ.c�;�!�� !����* (����b��E��>:y�
��qCn�=�7�<�)=Us�T�q�^j��G��Ew�#|�^�=�ۨLR�Xfz����xb�{55\#�p2�}�Zhu�Q��6߄F��YJ#�ޖ�0�x�m�����J|�8�����u�BV�~x��aK�йY��gɼKDð�rL��H�~VQ����.�oo�9���>~ss�ӷog�e-��n��.ۿ��5�e� �)+��PQ��t!�U��g{K�GE����
.Q7� ��ާ�rn�Іxz�M����E�n��4�j�*�s�(ZK���A��X�k�);�	�"�b,���\�1�wxr��.q� ��|�� ����?ņ��|B���j��m�^���݀i�){����������e,Fx��c�~��N���'���\?�\Ia`_�Hs��_B#��Iz�$^�c���Y�
k���X}]��q�����C8��.pv7S(S$'1�J�1����K���_ ��.ۨ;cNrq>h�|�JF0�`��+���l9��pV+)�OzT&��m���e*�\eg��v�CR���h�92���a�Khb]#����J���P9��Q���/{�	����=m�:��hk����"�V����R������	����� �
S5Z�xt�z�x7���e鈓���ے߂�ŕϾ>�@�8��Yʐ2������1w���+y���A.���mFFv��T>��
����V1w�G�]���U�!�a!�������;n��D�>a7Ez
ѝn��sN�������� $
�b�n"���Iy�&}mEPX��D���̍C ά��Tg�b>���yЋ�m� �6�_�c�� ���-3KӒ	5����t0���,)�U�DJp�}[�H�.
��~O�������<�D�B�͓O��c�#(����Ə����cӘ�� ��,�B����򚓻ðF�J�P�G���	��.��͓|��`[�D�]���&;��M >� ֍Z�k�;��*�������"��_ �0]�����
�c9E��x�o��߈�ˢ� G�N*q������Y3���.�R�7 3��ц�%���bV"z���$�ĹJ�Kw4�5�M��faY�6����������$y�H8���H�7T4և,4�*+C�Z3�L�c�8��{�En1	��jL
��_�MwE��j`��6g�e���K��6=T�}y��Ad�ޣlDy�e�*8 R���z8�'�R;��4x��(�O�d���
�0��o��pVV��hu�4�f�H���T����-d<2�J�Z�0�P��U��@h���*B7���{\�TE��j���y+�u���&[��+&d��Ty�:P��~���!�����',��x89GЫ��L�[6�M��78&��vs9eeNn�M�n�������ʟ��gԪ�6��3٠&���w �zR�'���w�L[e���7:
9��!���F���<,Q�r����)��p��3L�(/=�s�"�K�%^�c�k��&r�/]��,{CH����[�|R���5�s'��O���O�Px�DI��E`O�l�{��R8���"YIUM�xf@���Ǹ����X����q�{��൅�O&qM��}b䆠���=D62��oG)ш�b"U�ދXl �0�JRHk�'[Ҁ�G��YՉ��dƄP��r�ʢ�g�#m�3����jk��Wt�'�Ч�:u���d �7	2�u�,����)m9�ˆ�8�Y���bm��y�ڢ�Ch�³:��2�@�2/�Q�ȫ�0��.Q��]�U`@
W���YL�D˻h�B�l!��#��g�jF�bR�,a��P���@>�Pl�=(ۢ,�`?4��� �A"qy	��3�%)� S�Ũ˔ܺ��z�C�F��Dk��o�l��rHIos#�\څ��8Z�`������C���b#;���A``�� �P�0y�`v��Y� �	�Ddp�����H��w�-��t�d��a�UqC�3ں��3w��>�-/�;�(��L��t#��!ӷN���� �h�Fٜ��Azw
�"�߿��h��-%�<�g}ҧ���1�{a���۽�yA�Hl5�AZ>�T%��R�A�y2�S�b���	kOAqI���[&Hu�#���կer�A���\'������X����f'�)Vo���>~F-�]JY>�ov�$߀b�d7���.j��A���[�����䆻bu� �20�hȰ��b����g�����}]�ގ)�'����#}o����
x��/e?M�qM
7�ǻ��k���N؀�
�$�L�{2��Nih�b�*it�e�|�5unj��y�2�x��yǧzE�h��W|_����<5@�z�'�V�|�jOI?!ҫ$Xy��AL�t�y�б�xRcH#�z���p�u��[�=�i/�bcC�����D惇Gv���:�����D����9]! ����sQ�F^��*�}���������z�7:T�c>�^z����p�!�y��B1|�!��C����h�ˌkO�xr��G�? l��%�v��o��#Wc�
�v*�)�/	��4�����:���眈�4���ȡo�J�W6�v#�E��
�	>$xC!��Z� ���Q^.��w"x��|�#!R��x�!A�O���$�FcQ5�Gu6�����'O�� ����W���C\�r�����(/E���'�s%I,7f~���i��o�&ts&jr���k"�	H_xEn�YuǓi=��>4�1�y6T��Y�m�V�a��7��}ʀn�Ӣ�M�c�����}`S��Ͼt`SX��� ����C��k��vu�Ǵ�*�6���6�k�|+a�`�;�Gy��w��������'��a"����]����N[�_٠F ��<�k�ٟJ�V���ZNQ�A�?s��*j��e����3]K��vL��'��SD�T]��	̓߽�\������ӾċƝ��h�����hd����3����*h
���:�e®C��[x�g<��ō�$O�oŘ����!��_��+�Hp�M�W��PN�&�!Q��UMɸ$d�F�:n�����]�DK����Y�S�!��p�#�� ��"�-n��
$&a(V]T��������½A��v�
��Z�?~VFgT TC�>S�)3�&d�[�8���wwη��WR2�)�4��Q���FaS�o޶���P�I�ߕMbujE6�25v��I�3^p���h��`C~�/����O�l+j�������j�F�'N���/�cݫ��[
@Ǟc��Ņ���V�{�&Y�,g@�o86zaL��,Y"h�����*Bك��_�Qc��R������`�"��R��;�w�Q!_VH�Ba���~o*UL��L�(pޅ4������Ed��#�R��/��n�'hc�RWY�A�Pab7چ��Gl��4��}��-�͊k(АY�H�rC�|�� -LK�E��Y��b5�f�&�@�q��ėMFܕ\���*A{x[�Yߐǥ!�����ۉ%.')U p��MC��V��?���B3���o��O&W+<�wh�����Z�����!	،��+��` $�M��O����Ij/�4�.�������e�3	J���`��"��x�]���g���3��.����?:��}��oћzM�7!"G�6
�i�O�����2mTG�M*�_���	�,t�m�uaꚻ�4Ho�O�`H��Hɾ�˗���!.�U���&i�H�H��|(�W��%�����x&��x�@^�C�w�XW���$�g���j�i��������h[.P����p�eǶ &��+Ta�s���6���et9�²M��X�X����Ыh�V�A�I��GJd�q��fm��^'�����!� ���l=�dBP6D����7?Z�À��|�|�e༈�/��D>��Wi�2~`�ɫA�`������k�n�o��Igy�*��=`ޟ���-g8�7�P��{�	ɯec�TXW��9�@�Y�y�w-���o, ��j����cL��y��=��L���zF�J�wը��Gc�6��_��<���U����R^��o��e_}P���4���l���@F�gR���G��[�Z��a#���V`�lpKlm:������7e8�����$9]]I�	97��t�c�WQy1C�>>W٣�����ϕ�9@���E�;�:K��"]𳝤�!WT�y�Qn0h�p���D��AP����G)���&�7�艔�(�[X;�K��p�
v�\���Jf�X+;�8�r2�3��y����GB�������e�����vˈ�`g��Vx����l�r�y��F��=d�s5̏}�>>1������q:'�W��e���`���=�aZ�yP�Z5�A(شE�]�Ɔ�o��G������j�Tz��NF4~������򐎰��;3U�r��Z�:0LȐa����H�d���eHq��+kOvM���~_�`,\�A�I���G��`$�z��.m��Q�.�ڶ���};ՔF��D%�W��tVk�]=/�!�B��5��$���^�,���ϺTR�i��}��BA1�oQ]ޓ����A��A;ID�N c��x�y���U)�{>�n��<��:~{����N@�R�y?�G6C�e>"�b&�o����j|4�Kṡ�1������C+��y�A�\���$✳'_+���ݒ�.�K�Wa��)���T��OMu����4=]����������jg�I���X�>�1���С��%fX�l%/� ��[���5�g{���z���c,�����6#c�������==Dx�����SH�����@��R<lȧo󑘻���|쥇:�����t!}��iX�ZiUN�X�;Z���b���i�sF������1��=�]Mc{{Ý]L�q���tE�4X�w@�W�>R�t�t΋f��\�v���z|Z� �icZK�,LIMy���o%�C���S�on_�ۇ�� -���,���W�j�"?�����e��f���	U�����|�z#� ���zS[��􀾯Dm�_�MTH��v#�Pg�/VgP:S��Ԭ�Ԥ�P��qr��.�R�Qq�b�8�*�����yJ�x �ۛ����S��8��@ʡ��1�3ȯǗzg���U�ђ	+|C%������둁�)�/���v�w�!�&�f��,��o��4�K����*&T.��?�-��4`��|�S�W)�W� �U72@Q.Cbi(�5+K�5�����HX�|�t� �Z�­��Y�����,�$�@vqm�\��زC��l-��_�(.�{PO��1z���3��+��M�vF}�D�[���?��1�h���6��_��i�~�����Ln^�W!hs�K؉2w���],'���?&���?%��<�VjE�G�0>���0Iњ������X(?s�u�q�Sz����u���T��M3�AFCXJ�|�4V��c5(֍8rH������Fm�A[<��"҅Bƣ���\�i/�/v;�h0��&�mw�d��зt�vL>�6)�ّ��~1C���mʁ|i�M
001�d!64b��$��ͪ���~Qq`�����'�z�ʘX:Kd����#�7�Ŗ3�*��{$ I*1�d1"�ر���
(i�k_�N���i`��2�F+�7�xg9�]�ϵj���LlX�c�z�dvV���E{��Oeϴ��48VjH�wf"���=�vj3-wI��� �,�1p͊G]D��(�3��iq����(p2V��4�(�=HC�Ӹ��_�2:�ȝ��1��Ð��ڨby��4���[�m��=���2\��/���|&K&o�7�S�AD瞡Z�6���AP&�p=m����"���{�6;���!a�]*�\/~���7D4���Vm�%bH��al�׭��^��!���7������E�GW����ܼ��Fc��I�=$$t˙quks?_Bt��jO*R���.R�j�)���B:$� ��A�&=ԮRu���� D�ص�rKF�]4[شVC���{��o���A9�/��]���a�B�����R�'��$��~.0[W�갍�����K'��d)�0��+��o�P��j����*��:P�f��2�dKRޚ1�>�jO���Uc'D̃��+K����эy1�L!y�t��6=�O�@������{�I�-�B�qf��1w�Fj+����X8�8Xۻ���ݙөhb&!Q_���6O��Rh�A}��&q����"q�~xS��d>& ��Ul��)�V@�c�w�q�QI� }�n��H���&�b��
e�� t��تKM�S�な2�'s� Mm'�,�oJ^AüL��4����?oE�%�FOH���"��gniI�W�!̤�6���D��%Nu.l�F�RM��C�	�Br+Z�|�)t��'�@�i�������>��ZD�������� 4$���b2��^��X8t9�-ӣ�j�7Fn�/E����j��V��݋g`؋2�2[vKN}���S�cV8rCX�&Լ0QWB�TY�m��અ~!ѩ���O_��I6�?_�h�B]�F�&P]ҢU6cF)�T��)yX��.�`}}Al]��&��^����:��+5��4-�������M��I �*9��RM�|��Zⶐ��c��yr8����e�����o2(K)·��"�/�h�$�<��
L�ɂ%[�^�^ݭøw��ރ� C{������.Kkk(ge爀�ٵ_��@�a�����[���]�/�m/;Uw��?I��(ɝ�D����_5�A>�xˆ��pNMa���i�9}J�B�:Q
�cL���w��G;�U�m��x�qr�|���G���0�J�TM�ۣ�4�5x��$.��:��
:�����^y�n3�{5l_��p���z�2|�7p�4�=�W�L�Ub~�r���~���oQ
ƚ�O_9�C��v�Yʹa��9f!~�z�0��$��L(hR��q J4��r�K��}ޚ��R�I�P�H�ёra|6����q�f̫��؈F�ҏ�H�%�L.�+e���b�B}�~��<�pꌚ�톦έw��8Yi�Ǡ�')�E���7���kJ�������P�6oL�pm�X;�rձ|�y�z�|��'�X����)���N�\�ˊ��������y[���+�v���������Z��D�Y|��$��w�]���|:�����GO"M�"���`���`4I��6�듌�m'�&��FS�7 �l�"*�g�2�x��wp2�$uS$A����|��q��K����3��gi�+��x���%20���^�2��օ#��u�L���àY���{H�*ns����t��ro U1�#&�;0C�42�=��X9����6��(�AJlՆ+o�?�܋�q�՜p�Ĩ��<��XR)����e�>�x�C	��i�QZ��~8��q�p7*���{Qfsϐ�J�l_h�?�FV"���p�@ĬX��������ĺ�"f��ѩ}%��U'�$�Qk�,�d0��g�L���+�f��(�" Ni��`ƵT���z���10�_����%n��:׸���m��H�\S�չn_���_FJLK��]O�/+�tQVFy>g��+�B�6�c	3_6X{��j%j��>��2�����`C�{=�4a��b�<Ht3���o0'XX�G�OP�Wm&�$Z�\4ؕ�	���'5�����K�W���G^=�w6� ����k�%콘@�~�Q6�F��\��hQ(��F�@�ӷɤn��D�����J>:D�&��1�Q�S���Oj�;�����($)��������G'Z)��'�a)��8����>�/8�\�@3f���ȶҧ�b!���LnEU>�o�P$pږ�
��ԝd���[��2�(��,��/m؜C�(�Yڅ�ݶE�~`6��3�ܛw��°�攖s����l@�9O�q�QE'�}���bs���J�>�awOv��򩎬(�]��2�g���LT�2c��`�Q�w�x!�ֱzg������pa)�����0w����V9i�E@>y\�� �.�2� �m.p���m7��+�����/��2p���D9��vh$�J���D�od�f�]��9��������y��i\{�'� 6�m�0Q���}�O�V!��v��[���Zgn���= ?,�`�7�|զT2Ӄ%��b�c?d��m�����K�f�����͉��{O�$�	>�Ij���s�RA&�!�z�Р�`� �.�}�V	�o��UZ݇��{ݘ(�� %����������l�93��+����nn���[�q���=N�$*v��,RG���������*"��L�� M*�K�Q7\>NL���۪K��݀����l�i9���纃��(��zOұӎ���i�,����J>��)maک�r�?��0�����	q9�W�I��%��\��b�ou̝��r;�>��oC��Sx�]@�'A\a��q��.Q�:$��.2�<XV��D�D-�yz
K'�<M���HD���:ǩ���k݊4�鏴ڥ�kw��[�E�D	�髌�I>@���N�^���^� ��l$I�ߌĔ�A&��m����t�����m	c�HC✛�S��~��/l�3o���dl���UW�jOK�_���.2�0JZ)��	�#X��p*x��a�bH�g��K}������֨�k�B�	8!
��5�ħĐ<u?VVJLJ����^�N�%�U�����
ZVw�^V�`a/I'�_^��ר�O/tȦ�0: z�0�ô��;\���V.��;�T�l�x��S���ݕ��rz�oN^���e�G��w$�Mg� �,��4o^�e�&�Q��+D�H��{�P��� y^٫��[��2��@`��E�~��jͯ�|��܌yqѺ7�=����������WSAcݛu�V���K�q�@,EW�7�W'5!��R�^�(~��)�]3��t�B�R���9L��M'Z�I*�)�gP��Jd�2��
p��O�����Q��d�Ӵ=�*�69''��6{��/�Zӟ��f���ݡ����6�5q��_j�\jc�*�g���Nn����A>
D�"�bJ0�����L:Fv�2�A�������`��I�+�P�2I��G�����!��8�["��g��\�I���;rW����;c.ձaB����%�Y��m�!,�=�SMĔ5�S�?�g$+���,
�;�I��g���|;n�oa��q�)�HV�,��i��=������r
G���٘�r���Ղ(�֍��:DӪ䛬��3#(䅒����
�|�ǐ=�WVM���+�M�挠,�:�K�	����g������;ry��_K�|om;\|S�`��&���F$�=�'��9e��cbKo{���oé�o�g���I�wW��� �w"ea]�nx-�>��1����U#�����W�x����� pJ�%��@��Q��۪C����O%F��lZԶ�I1v:Pg���d�}W]�#j�t^x�M7%���*4�&�J �æ�LE�x���A@X�,z<��G��@����[g&dQz��D`�x���K.<ױ�G�G�J��\�%6�Y��W�^��f�E��K�pO�T"��_��3�v���[�UZ���3���+0,�k�
L�n֬�}����y�`'v�O#�����	���%Q/{�����%�-�Ь�c���|V�+
�c�P�kTW��lyx�vȾ r�FK�re(C��N��_B��,�?��ZD�0i;'0��hnO�̓B�]��R��(�!�H����t�r�.a�	���!�\�oQje��`'�E���G*.FԒ��O'R����v@�㡈.�&�W�.Z��z?�D_�w���
��d�2�ŵ��ݟ~��a�q�!:ޤ��q��`�U�E�Ε�j����2�����n�RD�.���:�8m�B��R�">�0�:;�X+(��'��!���1�|w�:��t x�Β��2Pȟv/��"\a���`|(�'����o�;Bb��a�^��H����"q�N�3��u�:�}m���w�jnɍ�6yٱ8G��a�9�o���"Y�}5�.'�Ri�*�E@nvI6�v�	��R������@�>R�aH�>(��Q��<�DyvvC1A�!ٖ�5�M�&i
�����~G���!`rP%i�9���T�l0,[�8;V{Z�?��p�F�[Q����.#��c_�31�͠��[ZZ5��fx-p���뷣ȣR������1��,)�$ntl�] �D��~���Oh��g�{�e�����'u#lͺ�_nv�ت&�Rچc5���6����i�<^��fL�S�����&G�L�h�پ�d��`I�3�� F=�A�]�jH,rJBD��O%� t��E^��?���5����4���2��"I�t��NB9��nҮ0m�B-�|'Ii�Y/~��zY��}d�l���)�&F��;���*�~�z֯�0��Y�i"0�06œ��黗��=�,L���`�6%÷�tNa���g�)^#�x�i�W���n���GS�V}��cP:Oi��T3 ���+��ǈ�L`QT}g�����/z���"?�?'�V��M(*�.���vx�{�����YP&�dk��4�?��Ҹ��wk�i��Nx��x�2w@� �3���?�D���D6���?J���f@�t!���;C�E��ηQ�a���N���t�s�Nm�W���޴�E�=���qfWa(�#�3�V
IƐM������rNt�;�����IF͍������k��V���ax�pյH��/�g�7���E�����tH[^3�y"�I�#���UAA8�06�+�F��tC� �Y�=��]<~�t�O[��q�L{��� ε_���u�<e����(j� �	���"�<� �=�:}�*��L�ꋴ��F����>��z����������4�eYx(�E{Q(]��z�9�Lm���`�D���u�N����67'�L�➟�HY����ݣ�����jP�4����m�tw�*�a�/,�sI�h�|��<�YMw`���D��n�� ��C���"��S�t��SB�~v㙷�Qe�}7)�����dܻ�p��/}*|��I��G�]>��~[��c{�Y;�N؞��ǡ`�6�����
������bq��V>�b)h�2ER�T���c�7�L>R���ABr0�
�\ݘ$�h��t����Hky%.M\���G�ME܏�[c�%m����06
J_�c�6h:�k���k��Ѫ�E�FK��lc�C+ua>ؙQ�Z�Ꮖʍ�<�d�$j묁�2�V��r�t �P����t���5
�%G&p�CG%w:u���r�U$!����U���	���-]�'B���1�d8j]ÑP���E�'^c)eW�l��/o�������rX�i8���>�Tn�`8$f�<�6��!^�i$J0n���&�y�zL5��J�Ks�+������~h�C�~6��I�B��'��my���ނ�f������@�ju�������8@�I�D2}�U�m�=+V���S;9�ȥ�?�[jc�gS�bq��^X;�JL4�tr�h�d�����4�	w��F���l)ͺ�> T,����\z6~�2y-�k�0tX�D/��瓲6������rƭ
�\v>A[­u��e;/ n�Od�I���c��rX�J�)P�~9s����j�'��|z�ZHJ�]��4�h1|���N�fb�X�ƻ=��f�?>��ɫ�w�3�o����o��j��ɖ��c3w8N'��%i{�}>� ��З؍%��2��6S��3`=��q�r�w��̥H�9'�'����Pɕ�&�jU䡻���\.o��V4(��b�����R!z�����b�<ց����1�O�HY��H�k�Z8}S��ӑ��P-%J|�ʳ`�P���H�G�����Ю�}�J��m����r��IM�e���n�j���?=��eS�0>�q�h9�-dh�2Mo�"�Z������yNwÑ�K �?tj���|�	��� V�0|�H^,��Ml��Z����pJ���~��BjI6|<��޼]�j�]y`�Օ�$�C�2�@����YW;�ȓ?��� ;��P�ȧ�������ˀ(�������8�\�k5����.5❬ֻ��<7�a�kQ�lc���=�w�,��tp�&�x v�	���>ڬ�{h�#��Y��5��zm�V�~�a��t>����q�G��H��^�,? Rb���C	[k��u��!����:Ρ�Y��]ױ��������-��KK5���Dw���W�q1p��'M;{��IiunmP���j/G���`{�e����2-��
$������>cp��
Iyf_�ɐ�Q��PlyeT�tj��$�I���kc� !�
���U!��1N��W�8�}.~��F�����kb�=��P>�����Ʀ�`��+E�?�c��3��Dy:�v�N�tnpݳ����V��]�ɓ�VZ��)�w�
t+G��Rd���t$-��)u�H8)+�D���o����ḍؗ:�s�q��o�f��R��x�n�	�ξ�ۊ�.�ϣa��EF�.��s�?z��{����IB��'v��E<^E����,��]`�3�X�^-��If7�XN�����ڑ�k̫�l��~?��P��0��ޛu 
��T�H�<����?���=0ќU7��A��	�?є����p��5�V��Uf^��H$%k��_�.@��.��mF�mt�k'������N=� ���.��X��~sa$�y�E[�*��^$/�>TᇾE�~ZR�ܓ��`�p^DONJ��pĬ����.�{�vi�Q�H/-����=&�(`��I0+����>m�����3��A�ܘS�U%U�"�74���Օ�]E�B)ݪ��V��/�{��TO�'�0�̸Zj ko_����'�����	����pN<8�����m�� �Q0(D��}=d�!�&�Ա���V�#�3�㷈�����װ������_������I=3���n��Ց�A�k�'~{��(�UԴC��ʆn��}�Y��c�
XKu�)�+�#(>V4�P�`�NV�/n����ȝ�:��C�2�ff�p_�� �����Y*�A��|�+�X�N5�0�z�����M��R�R�����t8f>���S�8��Y��{Á��Z��=&qJ�ؠ�.��h����v���@���Q��(^�L�F�~Ɣg�C)�W읋V�n�5L�*�a[�.��i^����f	5o�F�u�G��i"��eO��Y]�|�;�.o�~ͩ�[�Ҽ���Ǐ�J��\.;�Q�b��v5܄�
�q[���R�M�J+�(��d����2�4�D|L"�?�Z�����?$��$?cT�����q/�b��Ҿ@ֶ;x���m\������)%v�#�ҩiǧb�h�x�[]W!>=6(K!�R��0_�x�o]L�n�f�<��u�CT�k��[*j��y�:E��!���ZU�%�3��?�)�Q��#{���Ɂ��k�b�.U�+����.���N���^㗻�RBU�d(��K)��{����W�p4&��r�h��0��=�~�����v���C<xZ�i�	"fJ����@pHs���ߛ6��G��`sO��ȬZ��������_g�t
whj0������ �s�T�1�m�x�j"k��S�
�l��M�	�z��U&����W��u״�"��a��TyVO!U����]㷆�7�C�rȹ5��\��	)5,*�p�Zf�TR��k�~��s����c5vFU����f]����������ϙp�w�%�1�ȣ�QC<w\k<$`��W��Ұ�3(�h�՜u+ݪ�Ez���8���mنDs���}���[�ݹ�?<ǣ���:`Ԧ�,ZD:{���6�
��m1?����M0���4�55zGR1A��KJl�iDn�GSd�Gn�����5,�tѺ{J��{�-�<���������k,J&��/�ɗ
����+c&ˠSY�Gݢy�$�d�Is	=N���Xp.�Q�
[V$���Y<X~�4�I~�|��KP=7��A{M(�u�{΄f^C��T@t��-ń-wz�tp
��NC`����t+��ߓ~���(�h(���$���;��~�u�oC~���?����ě}��_��5��:��� ��~r���;�s<��_Tk���,�Ԩ��L"��J�_ ���l��A43�M~�9�0��%_RƆ:����[�JA�����C��6Io$x"���J�5swN02���/�µ�#Ez���0��.�v�e�ܨ��Au����i5�2N��b7\n�=�"���WZq�|3=_�c!�� �+�Ĕ�5lyr̎*b�!~w�?����"B��'�����x-N������C���ܗ �-��,e�]�IW!���4�P��Ƣu4g6nx�J�щ����:L�:I�E�^yK�#��o�g��L�G�ւݪIf@o��Z�Pb��ϼ��yYM��? R]����ͦu:��O���HL�$�u��ՈrJ�quhP����0�"�I��`��/%ZI�FDmǜ�Ǟ��u�Lt[u�JNݠ�K��Q�@����Ȕ�v^�W�����X��)6/̞_i`�aj}13դ�t��H�~�YIS���M��P+j��cc
����a�a��T�����j��K�hI�%��,���>����%�A,�7�����?��1P�!}Y!�;��o���I甛��箸ow�Ԋ\ٕ�Ӷ~��|��3J���%`9�7F�v�mK��ϖ��I�L;.{W)��������Xꨳ����qDO�3HoԽA��Ws�����,kY�k,�iW�%u��i�������Sc�S�7���J��A���c��؊��h�ٞ����i�W~y�-Fb8dj/l�`Vv����\��)��O��0��b\��.�bQ.(k��O��:��ȯ��c�'�ԛw�}}~�=��t�4��qAqF��$G�ZQ�\�*L	��b8>���Q���UU���@MқG���/F��ֳ�Ƈf�� ��j�eh�t�Z�Z	��_=�^�y��m�(�`}�w\3߱i4;�����J�xo�B����J��$��F�@NT�wQˢZ���w׉\���bCoW��i���X:V�Ɂ�u�Y����i�!��+VV�
C|{
`�fG؅��ڪ��As_��_��b�G�H�da'5'ݱ�#KK������ad�<��L��V�2,-�ysmVðx��FkF>2� �vP��E�%��,���L�R���,ɒ��M��~���m~��)=d�Ͱ�8��Y`�e#���R{���;z]a@Uí� �>L3�x��t?EGa&���+8�F��}%	�����@���Eؓ ܑ��K�rʋ�?��.��	b�1�G$wW�����j�e9�-g��M��h}⪊�ڦ2���:˜� ��8 rb�>�MS���O�7kR�9�r��U��<v45�����X��?�9��βJ���Ί1H��SUΐ�t��V~�d��SκV}g��T)��SA��6s1�_�[�L��yW�t�D �Y�[��H`��*���Tt<^�'�D�����fo8�ZD�K:���\�e"}1�Bż*_ �͒�u� w|��צ�q�!���"��J�Mq��h���0{Xx�ZغT�4�{����_▢"C��ٰTw��ɟ`���g�l�]N)��;�r#z�%�^@�0}"E7�
派}'b�dj�&0:?�.��I��>2E�ؾ�	�o�����B�k ;v�T�~M^�)}��)�<Ldk����-������
C�>tvdp�P�2��A��!�.����4�!�;ˢ������A�I�~�,.�ʭ|��<�ߵk��ĉ$�'���=-kVU2����{&z|�CK_cw���xf,ɛ̵+�aHTeƮA>�*C}�e���cL�f��u����C�Y�C6�蹒]!�ql�j���cO$�jL��JX��I֣FO������4�\S�~	8Y����vG4	������7O�~���y#f��0!,�m���b˷��Wx�'U��#}�pI�ڻ>I�oN����ne~`$��?񩺼��=ܠ"$��{�X,$�ԙ��R������"����_$��u5Nӑ�\Y��D�RAW�m}gר&A�Q���fO�v�Da_nq�Ǵ�\�@;H2)D�՛�XM;r���W��A㆚Z���Zo�P�Q�R�Ag�>��ϑ
Vr[t���$՘�/Q�kV	]��s�x=�U-@ʠp�v;L���X�OZ��b$P_�~����ꇅ�a5R����d��hO!�A_�K�����S-��5�$�{�%ѣ����X�-5�zȭD=��q�%"�����a��
�ЛL1�l�1}��'��[���`���"�1
P4v�!RD�Lv{c
]a��d��X�Y���Ϊa-�d�U�i�3�:��qB��|��W ф��UTVwt�I��\�p����8UVaX@No,[� �M��Q�m2E��:c�{��s���1��
���L�w^�{�*˄�=�M�F��"���5��L� $ŀ8�*N�E�v��}��So��l�� ��te��|;�T�z7� q�H�Խ��.���3I�aŐ*NW�Em�o����:h[z%�WA#;�Κ:���k'�������X�n~��y��v�U�A�j�t �2pv���9=s������r*&��4�_>{X���%�X��羦ݿ��s���l�3M"�
B�>v��K���#`roI��4j�3�����f�&�vs�(�=%�+!��lނ0���E�n��\�:�K��y���7D� БȰM����U"�F��]� f�\��Ν��2�9�>����Tq��f�gؕx�u�O֒3���c�����C,��|����Or��V�B�V:"���z� ����TC���q��Aث��%|C���ٕ�(\��1k�24��X�;�G���PY�|���� �O��,�7��n<�dQ#>����ju�Û�F-���UȔ�������$����LcI'���]�0�b����=VM z���&{�����n��|N�H�~I߭0��F��r(D�B��jSWB�L���3|�1���������H�V
�E`�矑�u��G"ʯf�� �:���;\�̈�y8��,E�'�������|�4�_��}Ź)�Ө����;a�����OQ��n���`)��v�r]�P�RhK*�*W�R��M���,~$�Ӑ(gZ�@��pw��%;��>���F�n��Z�d�蛕�PK'����E�d�~SҢb��z�"{���ܞ7ڴ�N۷�-�I�x>-�4H�W'W;G�J�j�۱n���n �o�u���]D�,�F�d��0ox8�
����l��}����h���b/����	t��U���}F&9(*m��)Ch?�H�ǣ�� 1d�6T�h6Bٗ�[�3{Ӏ(�\�
%}��aDC^,�]�$;(�p%������˝�r�Maw�nQ��'�����|+��wݥ�Z�v�Z�`�V�% 6h�t1��3p�}=��0�:��D���y��3�}4/�J��v�v�H;&�6��a׌��s-b(II�F����z��Y0��tuW�|ћ�?�,o3g�7Tɦw`�b����I�*7��
��9S�??�/��T�}E��_����o�|pĢ�̵���_�@V��{�J2*�.N̵^%�P�����1���6��s �k?�F�ܭ�4�銍�m��l��N/��r�Z��_E��*���SH� ��o��Q�؅�ϐ+(Jۓa��87���Yl9��l����y&$7�' ���q><����O�l�-	���8�49/�����N&�xXnEU�;z�(�P�����V`�,���s�VB�KU��.�l3��^5���i8��pd��>�;�d$����PnU�7��¯����b�5~/���d�\X��[H����o��w#i��H�~�a�"փ~�$��Lێ�۞��2"��%0G�a��G�"�n��P�m�`q�	��y�t���&�ev��Ж�8P7V��|X��H���ِH�[���T���^j��3Ф�C��,��A޲�2q�a�X��j*��w���T���=����~��\ecM��Vx�����4>l��-{@�}k��N�Z`�������5���������!�5��^¨hI��hD��}�wi����c�2S���]��k$qg��Hsh�v�@�Kj� Gy:\�����IR��'��Jhݒ�����!v�Ib�FVgœ�k�7�zSΡ��9���s!4�槹���ҥ�-9�>�֍D摇F�N�gdR�2rc�:0�ﾀJr�A^Kk(�hp�<D��`r�H�r��k�L��֥3��g�"�^�1���:J�Y�h�I�Kݓ�@kH�e��a�L
%��I��k�ſ�搖�~"F#����f9�1-/y��i���ț�WN�����^��*�P\� r��If�a4m�"S/�@3�-�"�7j[B���)�<��,i���8�2�ƿl_�?�F*5�����Q�P�Q\#���S����p�-��T��F.�	��Y)?��L�u̳�M�X�o�i��B�l ب�K)Rh���4���W���DdAr��T��̱�k�N� >38�CU���C�����7�u�'��y�	������±�u�[b0kB��H�9F;��b�k�ք9�8G:�,��Rfo�@���
��[q�ES�����lO��=̍�jf]�����o&�u�F����z�E�1y�e���%�v!iN�^��qڠ�h�g3�jY�8ߡ��bS!x��"��2<N��Y�$�\v��7#xa0Lvf|���r�CEŅ̯�gF�m�\�9G�jI�\!�҃Jl<>4�,�Ӟ�z�r��~�*Fq�v�@�ahMfj�?��v�4 ����^օ(p���nh�)�'�q:��:�<��RNB�M��W�77�\E�� q���>��u�ĺȲLӉ�@�E<ڕC�|5릓�k� ������G�'6O��+��q��U]����9�,�[�"�A9�z
}����� �#=�o\L�Ⱥ{u�^�	���$�f�.�s�[��'B,F{r
-��	��+�3>fp��~�N���L�G�u��a��^�b`��p��}�����N'f ϒP�������Z��wy�+�T�T4ɕ�w�)l��IQ�&"7��[9Z�ُ�V&�M��2-g�چ*k4f�n�W��O����壉A��&�%��;d*%��A3go��2�	��.��s�\Oe�9��${=���꣝k	�X�?���cJ�&f��y�c�F��
�!^P��hږt�J LI���T�DF�,N�6K]sp 9-L�'�z�e����7۷��x���X���{�o7�GC�oiC\�a�TaM�`j���(u?�P˨(�����.�N��I��y��P����C��m�Q���[�Ɣ���c��hl�u�ܱ�t�,G�y�Ƀ\����l]
��F�S	�1SN=���?��g(i����ņp�c�M��0�y������G�n��Q����g��!F�"��!����n���<���;���v����)����Qw���^�5Z��1G�v~��V�zI�K=̅���`�a���7��H,��1���k��)K
���!μ��)ㄛf>m��Z�V/�TC��f_FF%�IY�x&,��wm�n�C���)�'�5ݔ3����@,*P `#T+:���v���@��;�Kgq�A�N'�%�C}�R%z��q������˵啇V����hU�X�DG;  ��##RU��+��t��˄�CZN��h���3���V��9c�R�����z�0��ڨ��.IO��qW�/j\n�e�Ӳ:�㨧�z��p�'FX�M�����0�}���ǚ
0����Nej?:=����t0�SOު:!��Y�;��^I����*���)�,��?�Y� �\Y����r��yraP1ާ�P4O�ʽ�҂.�*v%בӶ��9�Z��}d��ЮQ9�J��ZX����%��L@׻���ˋ�o��?v��w�Q����w8�>bA5�:���⻵�5[��zP9�[�:�l����5�^y����]}�y#J���ΰ�G{�	EH$������@�E�$M%�7����W!4��P@��̄>������XĽ�	�qc�����TC���$��@x�w��;}e}�F� �*$=�	j�i�7�pjl-mO�Qy�3�۠�e�ߡl����ȑ���f����(�֖{t��R���M�6����* +��?W|�R��}�]��y��mxcm4�51�-��������}����z+�V���Ҙċ
J��'��<���P!Eذ{��#��W���Y����H-~�-����Z���#߬����2r�<����n���Y��n�|��R�ϯ�F减���'�86��t��U�䨘T����?,ݠ2	�u?,�/.�Hyu�����6<�U9��E�����Of�`6��OF�k&����~��_s1��'��v�wɢ����&��k#� 'K6��L9�j��g�7}���d��
��-6�a�Be<Z9-��[��A��ᥑ��'��UU
r��؉
��#]�F�ܱQ�b�	T�F��Y��fBW�v��*�F��o�Խ�]B��6H��;{�#J�s�V�/�>�L���l����:���}�����B�1Ͳ�a7��u%�i��f�^����em��%L+О,A�'���qa�ҵv�z�4����&�.�v��֝(�i���</t'�d��3E$�����|��������-����* S����n�'B���{�X�D�|�;���S3�^3;I	�	��}\�Lj<Y��sY���M4����n
ZYY�޹=��.�;b��Y؈�@G�����ԿR��b��@�]�;�L��b�ڳ��Z�O�[1�,sߑ�A�ҴS�#�k���=�A�8?���h��?���f����o�X����p�q��d�ꀞ=�I�3\�;fe}Dg��NڼO�����{�-�/.�~
j���[㉀S�}�<��>��A�$3�|�r�2]�vƩ#xS|M ���j�0=��߲g������0��b��D`��%��$j34rnW$�>7`OL���l�X�d��H��5d	��m0�����Om�ha��K����h�|�����CSY�*E���v��QF��t�f$�95���A$
}R�/�C�c���G��(�%ʁJ�]P�YV����!&u�=�ޗ�Avr�rkcpZġ.!/;л�A�uy,�f�/���!s���N�͔VU�ΖY{�k��F*`�Kƽ���:}����H �����=I�حa4���n�� ��%2*%��+h�M/���}�̇�c��?N�_c:`��1�L�26~�w�� �����ۜX{���mD-yx��N���`<��u׽���T����,�����g����	���s�3V�T��Jni����f�� ���p���D��*Ƌ���Fѷky�������}�[�ы�s��y �D�_w��ζz'`���guٍV���k>�-.�svU�����I�A�h�bf���}���"�3g�xj�=�)r
��ޅ�F�e3���$�0S���#N��<MQ?�Qu|j+�H�>�����41gS+2��ǟ檨�:�	�	��M�[��H[d:�T�~hl�hܖ���/Բ���*�!U��*�K���D�b��R�>�_>=}�0���-i%�!����A�ynj�iQ;Z�O�Jg	OQ+0�6�]S�C�g��m�z��?��1 y ;�"�R�G~�f4Q�	�Rl.x4��;�y�*<x��1�x�kpK^�����:Ц3�ib+1Om���r�D�������:A�K|ɐ�H��a}x+f�{d��y�l׶�.�^(��YZy�&��.*G?q7�f3�p����[0>�s�M��B/Z��Ű��k�-C�tH{���|��!�}@����SM;�m�d	\�U_�W�FFIZ�f���9B�'�^�A6�鏺.47�����,��AA��?a=���0j6���f�����K�^}���\!2���c%&ۆ9�"5�܂f��	�T���/��P�e:���-.�"���C=�6����3����޷ni<�[R ^��V�s[���p@�����PH2�C��t2����	,�H�WJ	OD �7�.�&A����o������������ Z��q7o͵�dO���n�M j;�Jn�ka�C%�ʥϖC+Z~���v�8R�/ݏcz�{�{�=��d�<�k��S����TI�������eMl����L����S�ݗI40m���Q�0jrEõR���Z
� ��jf�l�XQ���o+Wa�E�q���E�}L���
f��,�
��� �F�|L�S�j�d��H��B#ڈ����g�vG�{.*ɩ��Ϸ��nd�$1Y��o�7�d� 	d���ƚ����� ����L��-�Q�����UL�fC�zb.�0�>�vz �w#��B3e����|YJ�I'lA���'|W�~A�y�bBYI%J��ǐ�!;�p�9շ�Q[���am�w)_���A���
�cNf��S�b�O��B?��s�s��{i�,�K;�{�ב��M�K�B��;Ȳ��L��+ei#
�_؛����������ǆ�#�0�j�i��])q�[���/ʡ��4���jҦ�H+Z�^^N�H80��0j���
��dk"��v7��(�qB�4�-��g���[�����0s��}��"�=�S�75D��+Ƌ	�U`�Ao��	bC��zF6٫����r��Y�O�T!����O�d���)�x�f�MZQ�Z�!lܤe��u-k�F`��ur�?�nJ���;��A<��55C���Y�����^�L�$��PF�aX�e����(n���;s��䁬@�M�/�ʘ�60�{�%�M�"�`�y��I�dn5�W#���˸_��h�I�̓�yp+}�����,������Ⱒ��Cd��r�O1N]�*��c*3Q��@��-���o��$4�]ޚHV>`
�dM�X��@�k�%!9�nȭ
w���n�������hĠ/�m�Q�x�P�_GC��]���{$I���4�$��M����)�mZQ�ܽ���N��''FӦa�5&:{�`�`�4��M"J�6�@p)�6��$A�g��Ȋ��T~!����2$�cS��x	\�X��W�hpƗ���2�8� L�n|Lq��Ґ�t���6]|�5#r����W�D ��P5�<6��/UG�V�
�ɓ�&v ��v��c��B1}1�<�KP �(ϟE/�S��-��,�yp/�;�%�HMF�k��&���/� =�}�����B��MG$%E�cؠ�� ��(u�C^Q�"����z���������	P�^�G�fl�V��}qH�m2("h�o��(K�HnVI��$���&�5��'��x�۔:��5�չ���|��D�:ʧ�rh)>&<ʺ��.�]��?2i1��6���+�v���ӄ�t��9�_Yh���ۊ�NBr�A��EHX�xi�܁=��
�g��{��q�s��-��ͻO��<j�����@Z�/��$�|�Tp4�{NT�k�I-$��r*��Xz�z�/N'%�Q���_��	�4����-[��a�Lrج�.:���P���8��.99\X�F�Ȳe@�� ����UQ[n!��΢c@畡��v�|Y�I�<lL~�ڬ/{R.-,W�T(V��O:�L���)/�iH��p�E�R��[�srw��6��.K%0�hi�s�ބ��`8�"�xĩ�ʝ��(kʧ]������V斿����x��4i�Py�>ז	��� ���= #�fL(�a25MV���E�|h�L�U���=NL� X��p���[���hP5ʌ�h�xWj�� �yZ������on�ҋ�ng����mN�x}���#��{D�+�A�wd����aŘMjᮍ�/?1��n��c�1�`Mlp���(>�g�S>�W�Ew�P%�Q|�A�j2WY�`Ӑ��,����k���}�.��;_�D)��fpc�����0�|�
v8��[���)�akm)/	��7ፒ��A*� :��S��
�M)%XVV�ݘ@��Ѿ(8�b���=>_� �S���4f�-�S�Y�Ki?W�]�b}!�)̶��uZ՞= ��tfz)y�2�n�ƪ���*Q��a#���<�K,��ց}�4�O���-�j���U�wp��1p(�	��l��S�i�Ϟt��7_l�%��bȫ�Q�@��81kNC�"lP�����ԯ�J[BܱKΦ�BF{n:g�#�D������e��d!���Eg@�=���H��:3.M\�_���Wn\��A�tP?���u��	l}�KI�Z1�����eD>[�pʦn��Y�v!�����֦wR���\sUE�f~���;������jkl�U��!ҩt޴����l�a�F���%(����	�tb�ׇ+�����8��+��,ve���6��
����`dW�řƹ�i��H�J�0�Q������թ����J@��j> Q�=���7����;P�YGl}�V�0�Z���h���뢝 =L\�&&��j?*å��5��k��Y�C8%�~�65��k�r[�Cn�1-8��ˀ�o{�f�Q�ؑ�(t��Ƞ���Y(�g�Z���Y����mB��m~���*�'5�f�V�.���e�:�S4�JQ�\��S�H�W)ɭ�r)D���n�D���X>B�����]b�]�Ɯ���Z�&��zI����gG���)F0�����k"���@9~r��ܞ���f�7B��{�F�5�!O��$�68��:�h�X�����wBE!}��k�6{�S����;wX}?��L!�Ɏ����,MR��x1�g(��V�pP����7���n^�0e̞��k�����8��'G�2u���Y��宲�,e7�45�8M�|f�H)��X���)!4�4����M�J�b�I+_l��Y˻������R\LP6Gd[��s�����w��Zwݧ�j�+0.5m���*=��"��0�Jŕ�T� ��9ީ�}�%ɻ<CY��h�C�����l!
��{�(;z�M	r�k8���5�6
ҢM�-��4�E�?�1��Y��0��š��K<R���`6����qy����qA�Wr��GJ�i����#i�(_�;|����ȝjQ>W���ܩi	)��L*�%#��c�P���pYX�"k�\�H�Q�gٿ�J7_�Pz1��B�nJ���º�D(�N�����O8��Е���u���%<w@��a�/ʯ�G�q]�O�z].GkG�xI�U�HA��6��=ֱrp��5(?|zod�N����ߡ�x�u`��:�.,y u'V�p�6O��'������c߷�6}H�C�����m�P�(���I����^n���eK#4-����ؘ/��z�k��7��.���B�q��~T���Q��KC#o#��a^���%�p�~9?�SB��@�9/#�F����ʏ&ry��.�#Zz��.t�"����5z�)�	����	+�J�2��C��z�3��I���@���
z��U]ށ�`����,J�%�#�#��Y;��ڞm@az�#��|���lG�[����åI�w���@}����~����c�/l�r�oz~�}�o�Vu����|���@$����cW��(���I�'��+r�&�*�i�����S�.���X'b��X���J�f�h���E��&a���gvŒ�M(��	#�ZXa?-��0�7�W�?��K̻���֍~f�j�d�N��x^���d~;]ȗ����ms>����� �T?���L�7��W���漞#�M	��tg(�� �cxe���0�����NJ��Z9��WAKF�p���Po��b����ۜ���ėa�FI���_��JFwl��&e�������9B����77�{��v��c+���h�: ��0��C"u������D�����t�/����W��!�W`��r,�YZ����Le��>�kwS$��d���d�tm{d�p`aeU��K[T��~��h�O"/�U�x�I�),z�w�|Fo&����؝��e��9A��IO5{��@h���q*�U�rd�I�`��ī�v]������D����[�Iy��h�I�ٙ������_�\�ݫFH��@����-���Y��
�$U��O��!��L�<�FHgX�bތV<oT�kX�	E仈Q�����\�'|5h>`KRn�Xtɜ��q)e `Ց D|�dMz����D���*6B������b_+i����(�$��+��p� �� �ٶ�KJ�?r	�Oa��̮�$d(9�l�����_E�-C��+��DB�~0�bT���>�)s����gMZ�PQI��G�)#FW�E��k޷OϾ<qm����ms�Zt�ȩ���̝��z�Pab�����|�"A`�M޺��d�Q�O�9��|�CW�T>�5�<��9��B;Wx�+����@ٔ�^�Y��|X���� N=��Y�Iy��Xg3dΒq�/��V���{�>i����LY3@��T���><}�\@�;�W��FL��QXM�h7y�7<|g���*�V�)�r!�g�"�Ӽ�.�5_DU�c2J�u��j��{����^%N9b�^�棴,�)"���@�GX��I�1;M�H6� hۺ;T��6<��s�隆 w��h�"�s��%��Y�ab�^ޭ��o�3ߋ����J���^���)@A�+yU`"��u�߯�0_�57{�tS\n[�!��f�4�O��_B��2�#Öf����_k�A�6�}�T��7�zk��1�>l�g <�ie�Ϙs�j�r;�+D��n�o��K��IB�����T J���vdnp5!�$�Y�/��񽭥n��R�)�+����a�[����d����"j-�<0'0���y�[~�K�9�q�4�'w�y��O��a3���Sz;	q�O_�`�Z�&����޸��$�E��2���=y�Һ��@�mC�
����}/����wA��$P���T��¥�o�k�Z��twI��.�+�5����m]��l����kP���%s��M�S]r����KJwD�wg|�J���,Θ`�`p{/)�q��9��ׂ\~j�t��)��|7n�����8b�:<�kt7b�ȸ�%r*�������;��[�����+8�d��H�#�C��!.=�� ��=����ѧ\ڒy2x�q ��� �2Ⱦ[�}* 4�O]�:!>�Տ01��m:�<=7y2( R�}���:@�\��	�ᇀ=kf�ꉐ���IQ��|��Msy��Q��$��1_�@��-h�ѐ��]
̰#���/BK���5�o�E��֘ɵw���R��D��F�Ǔ�S�?��)��=6>{����8�J��B{iƊ�����Ϻ7��J��9?1gP_�k�"$S���L���/�� ��«�Q$��.i�������<W����4�HU��۝�N7�����������`O��]^c����6��2�|XS&�w�x����N�
�b����H�O�A;gɱ��ZN��F��ý��K�t����yn�}HU�?�]X�	��F����m/�����?�,_$��ƌ�1w�k|��aG�݆+�cޞq���z��ǰ�YFg�e�.j���g#���9��rz�-���_E�CsfSო-a��6�����Te����:y]`�Ơ�X�L�ɂū�:��)5�K��m�����[����S�E�;a��V��ن�ߏ�%i��B��@O˂�����s�<#�JgpK�ؓ�7�i���9��7}<K����0����#+��f���7l�ߛm�5�x�!���O_;�Q��Ne���� |;�έ;(f�J��C2n�[OЅ����斑[t�����/�5���l�r!��f��Gm����.9DWK��~Ysc�No�4E�ƮV`�$�J�g�Ohaf������~�$�9�ط.�Tn_UF�#lSe�c�H����q�{®�U�Y�0������ɏN�#"�j��K�*��l��ܐPܹ�t�5�*����?Q�\��=N�s�9v��.��O�OG�HjU9�Sp���L��l��ͣ�O���X��K��S`{�Г�DW`�v��{<�(�T"����M�1 �����_ {^���e�Ik�b��Y�	ϕ�l���R��aQ�Y=���u���J����<bbi��>|�ѯ/ ��2�����mU{��lƐ�y(��� r�g�1&�&q?���[eC�g�H�?ߕ��������-4|y����4�Q�'�b��X�Q��1�E��K����d�_/�
bd$�O�]�fp=�n�P�o�������`G�>2��=wI��ӡ�)��������W��i�� �f���Q�y������.�|��6����Ĩy�ǜ����a^!�:��ȱ�T}4�q�ҡ��	4�|���R=c_���
�,BS�Z�G����D9������|�c�Sna얣Hƣ)��\��(U[�
N���ˊ�/+��lG]��m V_T�D��9��_�[�z/L|Hp^�P{��M� ;�k~ږh4��߉�VB��֓yY\YIT���ڐ�P'�qС!ۋ粉+^��c�ޥ���YE�h�:ֿ�0�b��� Bw�f^Y���]�2���z�"'���z��C���T�:Cl&���s5��ϑxƌ�ΏӚwD�oZ�t�,�<R�k��a�GD���R�Ze�Dۣ824ʦ%��� �G��&�?�����o����X��g��N�������'�/��gm�U�����6s4L�:����:׬���q�p7������;��к0M���I��qs��H�-����hW���b,z�4�h�N/�|A��Q�.���_v�6��X�ˇ�!	]jD3-�'�����\TY0��3�`ML��A^���H2�)��[&#�ۊ<�:u����v���F�]�	�i��ƉF�]d1� ?M]&�(MN����VmU�UE"JΨ14@ ����sc�Bq�S���0Z���x�x�e�0��`�r�B�E!9 !*��#�y4��aA���-Y,�T�?e-1����B/���?�$l�=.xvd)�f�_��ERc�`��r�k���|����ZR��I~�x�+)���X�9��e�x�����hb�{�IW�ǁR#����� u��TA,����V��^Se���O��I�&��8 �3��ڜu!�L������38o�U6#ԭ�@��� ��I�e����'�aj�4�r�Y��T@�E�(H>8�,4�H��$�.t���E���ӄ��n��K�Uh�Eߓڸ�{>��o���E��á�!-aY��������[[��i�[�I׷8 +��j�q�S��B�w�����i�*�ۼR�}\hN�Ҋ�M���ve�Q{�^�R��Vu:��	-���	3ð�z�Y�����=���X�b7�j�������5��X�k��עͭ�Y�H0�pn�b�]�+�н$��4��\��K.2�0��D}��v�F���j�3vi�PsW��	���]-X+xj܊�����{�\GF7L���%"ܸ�1J`(�:Aу����|Ml?��s
Y
1[���s�ۓ36¨RS��ع|H��,e�3�5�����o��oW��݄�/"`��eUGxI9�CF��a^�������,��Ё���\p��Zu��	,�7@��%��g��O��c���_�E���=�_e�.�%<��hW�&���O��d��s�烴M~L��!M��0Ҭy�N�����]؜��:�0�ÁW��E?z��ٓy�	���g�R�j�so��1�2St 2�_P��G�dIXh�y���9���d<��6X��S��8�D��U��@]o�W��� gY�o�����E��}r$B��{ܵ�O��o���tNys2�Q)�ϥ	כm^Q��GSݬ������[�ժ\����Yp���&���!��m�"z)���
���� �q�1Cܶj�cܺO.�R�u��Pr�PP���.F���i�%a�w���W����?�O6r��c��Y�;G^$�
:0'�=\ �<�����,�$�N�4������"c���=�j�:�݈qgKi}����9 �#>�S�^�w��(A
]1��&d����mb�|@�J��'>�3�V6~�����;�w ��ɍ"j}��=F'����#���j0T�g7^����w�&�,i��}.�����>w�Q�P$=�C#J���X2�8#����9������q�L�+�9Y�`|N�5�.�X◵���n�'��'"���~B8�'���S����m+DyjfO�����p���D4`5 ���G[��]��4�������X���e��X,�`�c�<X�j�������i|�C쯈\�a�"Q����������I�xz��x�rL�U���+U |c��qpl�
n�������'���<��%�\���Y��I��2ئ��+�=F�S�.k~O�sʮl��S;��N�$N��S-"�N6���;���'7$��E��t����N�|`3���"d����@��c�����k&w_���cbQw�黯dC�m��M�g�p�`�:(�������x�Kx�/m��8�h��X�~�~@HS�����W�Rb2�پ�g,rt�.�������M�����i���K�(�Ok��gЕ����w'�V�q
���8�G�9�� y-SdF���	;��&m�b��'�M{�<�m3(�G�����P��~sw�s��BElȚ�S��.l'[U@P	_�$Q ~�s�3�pא�W�e~�0���p@>��6+۽����](���<���2�X i���{b|q�4϶- �l����ϯ�$��M~ߕx�N>�#��G�@&gع*�$O��ʆa���>�	x`������)��}�S|&�$�*�_�o�\TCP"�cB�b>�0M�� ���ܶ��D�~JZ���I%�y�~�`8""��k�sE�a��B(�%Ú}�y�^̎��66��p�F7�|��y�p��6�]��5�X>��{1�����W�9�j����J�t5������ۅ'�B���D��E��|Af#C-����mG���(��ϴ�%�1΅��F��2��?�qzj�oT�m�K�����At�<\8M��5p"�u\ S)Ϫ��\�[rk`p퓕�}�q���1
%vp����|�F�����!O*'	�n�@���u� ���n8�ch�/k�/���W볢#���ə��1��{�zD�@�qȍZ�rE��%T@EYC!�G�^�HB�}�	-��ENY���L�VP>�����֬d`]�~@ 0H�OIC(e�N� u�qg���F��I����ih��7��#<�
Ɲ=\x-;"JJ�����>25�M?��Z:'��y{صB��ܣ�܏�]�k4I��&� �~�Z]'��r�ަ?�U���aT��8�WM���?Q�_|�=)�_��d�̢a���$�]�\,D]:�ܙw=S���>�ꋰ��r?��hvs�2Ni֥��*D��7^���S�:��镻<��
G8[jEE$�Fr��`X�A}�r@��?a�"���_����z��m�h���}�1���Lވn�j7�,�]������	(���aA|D��y:z�x^�c���yJ'=A3�7O�soF<&d�%�A�e� Yn�_�0weI}{&1&�ϸ��u$7t:��j�MOx�ai����&��=��U#��h�L,�4����Ý��+gEbP �іm0��h������n���+ey!��6:�a�J�vR����WU�I�B���G˔�������A��M�}R�2��K�@�\k�*rN,k'��7���B��'Yc�s�j@�ʗ�{O�w��r��B*p7�:�3L��:PJ݂���(��� *���!W,٪�/߰yWBq�������yIh#:�Ѕ�4��.ǡ�.F��TB�L�������&e��@�O�t̕8�YU���/s=˱�څ��1�Kz��T:<��	�������1�|Ƙ�k\C�ґ"2�>�U���CJ���T�t��\E��n,]�r�̡Sf6uz��l�u��bU�S����R��!<���hAQ-�%�ׯ��#�zƱ�h�>��%���*��I�!He���AJ)H_a�&j���`H��=F�1�6c �l��/Gi\��b,��? W8�Vƾ'�M0�OO+&�ֶH�za���og�����D��K���И	�&��	㭙��x����w&X�̖c7�8�܋O!B��С祅)-?օ����~����Q��
���t�@opvR��;��B
�f�8x���O뉜��׉0�_B�6���(��z
�
W{�_5� ��/!��Ņ����O�������'���̯��[���R�C5z���MG)&��{]_�+YX�>'���B؉��8J^�E���,���� �*�'	�`�y�Rۥ5f�d���1�k)�&��VDl�s+'3�*�BQ�Y	c_ɝƻi�rc�j(h�R6���u�\0��|�R�@s �zTE�]������nk�K���C�Z�xB��M�':���@ :�W��+�����n{�Q|z�yAf��Z�~��������W��aG�N:�v��цe�9\�2����3����"�:�$��B�.�i����w�œ��V�M�a\���k�D���U���{���l �
��I�ouL,s�2f35�FϮzK� N���ǝ��h�xIs2�z>ܰ��ۤ�0�zM�A���	��%r;`�vմ�d*g
BV�֋cy(y]�ʞ�a�{� C�����'��G�_i�_���7�����{�eٳ���G���qi�Oœ��F��"��0�-H6�,M�	����l��<�`�3L�,�B'm��kȗ��u��%�J��^����d�~����Ό��|�P���f�C��s��T�0��Ѷ�z��-�Z)� ����n��`���􌑴�>�1��1)@��h��h�܎C�6!�g-h^��P�96E���2�AF��Wusu��OUs�Ձ���G �7!+S��hW�*+V$��"mPH�HA�|�5���W���Ύ9������\�n���Ӣ14�TǙg_�r�"�Iz]�����A����B/{���O��i���M�{�^����H��:��On��{�P��m���0��G���MHP3ܗ����Ǖr8�� �0��`"
�p����l���0�N��.�(*����T	�Y�\;1GM*��_˃�ȏ�"�Y����:�l��#�[��eG�k�74�R�o�AW����B&�_f;7%�$Qza��.�����e�p�I=���I���`8����E:�[�qÅu�nC}cf����j�P5�qj]PO�2Tf�m�����av���$��� `ͮ1Ė9���.݁�����p$2p���o=�LʽcF���l��n�Pj��&��F����p	�����R���቏C��xzN�H�RaO�x�PTW%<Jd�T�쁵Js��֒�3<�B�{�Y^V��Ae�	����E/���&�����j�����:��vE*־D�	��#���v�h�ٟ�k1X��.l�a���m�������:Ah��s��"~��f�ۡ���rIf_N�C���~ֵϕ�@���fr.���%�_�����	��+cp��\��;���$U��g�����h�ڻ��H��ԕ�m�ɍ3��[Z+% ����L������BF�����1B�2:3������� R���E�x�N�-t�^e������+հјq���RX��]1h�ܻ��_y�yGj�(��i���Ѓ$FW���8D�*�E� 48�z��:�En-�nԺ�8�p>���5z�]4�J!3��~+�ȏ���m��||c'J0p�/J����i�+��j"yY�p����F�o�,�cӮ�x ���ɾ��e��G�����7dR�#��r�����f[�,������d�_@��u[�S���leg*Ȏ�wZo�*Yש�?t�5.��I6��FxY����]
?Y<�l��l9t�`�L��\=��C5�����i��*�e��t��<�Z���
Wb?����� Y���6�s��=htI�mͩ@������O�B}��,+eQ��֩�n�k�t�_��B(����m��bf�L��{un� N:��]���JJhᲣ�W������k��P$8�\��%�S"�w�ܯ| 8Rh��P��>A�?
��Z��k�KMt-ݥRב4��o��B�k�zs���$��xhq{M�몷�6�tS������U?,�������'T�����.ZGR��\6D�oe�Ma��;��OseۃkԇQ9a˲4ŶQ�z��������z�H��y��H㭸�CE��,��i�S�Jǆ�.O\Ԓ˥+�F����#6�䉒j���KIN� ��n�^���. �ڌ���V�B�x��R�����4�<tHb˘S�ch�?n��=��k��^n ��&l�z�*%i`��F�y�fc�<r�a�s���b�؊>Y�!�*
Gc�'j�v�#��Y�+�&ᆺ[�g���yI��5<E}�M��B��J5���ԅ�X��7�����2�+,���P�3j���Y�.���$�=���|T�f��C�I�@��r�ch)�O������Ձ�xw�}����4U^���/<6�@C5��rbb����K �\����Y�;��q��ԮwB􄐇~&#�9g Und�f؃�4���0�+d%�CG��k�o�|t���\���/s��%�,:
�*�M���e���W�q�?�^��_=�Y}W�r=~zn�i���N	M���?4���+�u(���C�
C�t.��L�򼎕V�>����M4����_��I�1�;�Jv~t���#,L]ܳ̉0T�bKRR::PV�aJ���Z�5
���l>p�&�A�x�S���y�]b2���g���o��JV�[���:��L)������	�����%�?�nn���b�N��(�l)�U{��;�8=r���1��>��8��#2CGΙ���P͟Q�*���;f�щ#2���ݾ"o��FSIuI׊;g�og�%�DMk�]�+����	�+�;6���P[�:��Y�J��.��htK�j(��^�0��oƶ�"��{ή��Ú�
�\�z��0[��G�-zއ��_s��^�kt���-g��xv��&t��������a"�ń��A��䱐n̒�]	=N���0�~��B�����+H�[W��$�8evf�Z��5���6sB�����=�M�ˠ������dݝ�\���i<�5t���D[h:���N݄݉}�m%۸<P��"�Q�S���l�^3D�F���h�p+�%|��L*���Aėo�7�~(fct�0��▬�yi�
6C'��:=���J��u(N��X�b�D;�r�?�*":�1�7�cͬgG�g�G�E�<�k��T���ԍ:�o
Nt�Qy9B�B���u��R�>v��b�D�dd�X�����|I4 #�%08ns��m�g��{oEV���*U�>4X�\�i{�6H�5�U;)��ˣ[:p ����w�˺�����?�h7���q���V����K}�8�^�	�4�K�5���&�G[P�TK���XZ_鿉|�IS	J��7P���H�X_��V��W�d��8,nhK� h���-4#�j^��9X��}Г%J��}�k����mϢUV�W�tg�x��3�c�F���m����-L5��k�of5�%��賰|8��>��̌,A)a��+�Z	p�����{���-�,�8��W�Βߵ)��L&�(U��\�ۣ@��E���^zc̹��+A����$����ZC.���a���T�n,	��H�dc��CA��ǫ䱼DֆC���峪wi�Kx��ǩޭ��L%0���y��5
��a��[,�2'p41����I���1���Kw -����ѽ�m�e��������.x�Bpv�Za�N5��H�ws������ ۷Z�$Xe�;C�Qۻl$� ����,Pz`H�7��cET5������A;0�Cz��Y��)�y�=��#q�0!�G�T'>���pMc�;��� Q���UYy$~v	�g�S��Y��dU��3��f�.B>�o�K��k(�Á�_�7�A�[߈c��hO���cp��K2G���'����B���Ƿ��Z����ѭ��n�z�Ό�zc�����?ڥ��`���t�qZ�%E��Ʋ!��I�iW��S��%d�k'�����AW4��ƍ>1~�(@�X��%��92�1ve���+�v�	�ɪ�����sݴ�@�D��
+��:p`��]]�y"B1�ү�^	�U_�G�0~�
��U��;`RY��x!{57���*�܏]}�k���
t��-TP.Ry������;���:WZ-M4�G�o���g��J�y�x��]93�+&��ɦ]Û���i3u�q�xh�j	��#���	�z��IG��6�"�E)���Ƣ��!���MH�k��������(#'��fN�\��8=x�i"ݒ�?���W�[��/�6��\�3�l(8g���_L}�-(r]�$��XL�:�u�ݴ����}��ƹ�`?a�狖�Χ=%�����y�$`"�߆q��YeA������l�N��mN��~;hY�t�q�G�gm���tu�_�b�{[�U!��i�)��A�!N��䉵���d�jB��^�r:ظȁ�y�R`�F);��H�C������)0�U	����% ��r�=��[�}_Mw))(mc+Ǻ�w1/U���=l�3�uM�@qz5��d	�W��(�����y+�&�ND�4�n�z)T����GKvQ��Oă�k�"f$ć�!7��h0���	wȧ)��w�C9g�ѩ;�o{磳�#!�g�FQ�P�5�J�����9u7Y--�aK�ur�� P���\��jp���4� L3_��0�{<�j{h���x�Rx�y��Ĩ�(o4�K%ǣt^���=����4Øo�E6�v/s��^�9�gi�%�3�*��X@�u0 |��%v��'�iU:Es�@�Y� �	�Ev�4��+�֊�Q��^&G��1l{�]�a�����xqW�T�j���b���_�vՆGu4�@��'M y���K����pE8}]��uze��� #��68���-�)�k!d7"w| ��0Y���v5��͵���
�r���L��.�yA�%��28L�������<.Z���R M�������mp�BN�㚿E��W���#)>,~�Jj����+�w^
�䦍și��jȇJ$.�x
n�lA���H$���<d^�Vw��"�a8���zw��.-|O�����a͢D	4� �?ӱ,��4�1t�~�Spi(z22[U��/�-Ȕ���1�����|�1�JW]|f"�iq:�
;�`�s��=�I�B�X��rS���6'��k/uݴ���u��--�f�;��m熙���Nb�����L��FQo�H�f{k}뚽�ߖ	����l �ʄV�
����W��2�ǫ��`\x9U�wr��Vb�ը� Pkǫ}*�$��[��|6�ҕf��+#w�
�a���*4gz�uc]B�� kxsSwA����d�_����]�)"��d~܄���#ᱎ,W@�֞X�_�C�+ah���C�n����J!�^-k�x�d�A��lP�e��yʆ�
�[Y��$�c0������u@������w������|�lp��G
�|5���d7��Vd�<��ZPۿ���h�z7/���*����8Q��	��l"�L�P@Yh�6f�&��|��!t����MK��rC�p'�q�o�a�ߧ Kg����+��I���42 �|�É�����e�
��/�p��Z�hi]��/�I`��N���@�N�{��V�f�����¶�8�ޑ�l�}�5�$������A{L�j��t��2h��j�	�����p�#.��XR�h��w1a��| A��&�]#A��~����ڼ��o�@g�A
�0����~���<
�s�;PR�Խ�5�h���_}ko��ª�i�H�M�V�1�e���>��$�t��~�v��F���~�G�-��1a���Ք����/3E��m��v��;�O?cfc��]�B2�j��(rC�֋��Jg�5��G-r)�	��\�[�G�։��{:$�t���ޚE"۴�A��.�wT�9�����%%�D��>bn��I�ܵc@	ݡ�}��7u����	���<�2�3H_4Cd�*�ҽ .u:;��. �-��H���>'�>��/�J�"�#����Y�#E����iŽ��;���\r��{Q�Ly\�x�pNsO}F��)2��ez\נ������"������8O����Il�K�)�G��q�X]x)ʓp����������B�@周i�h�oA	DQ�#�zno��3A����	Y/�!PE�P���4�q;٣e�$��6�nɸ������\�76���=0 ͍3K͘����	���%�r_8�Wv��7�0vu�۾�����T���k�J(s��)�GX�Q�S@Kay���=�$�}m*�7�m~@ibcU��S[p��rn����.��Z��&�K5��{K���vGk�d�5��Px�L@aJ�u�������ؾ�DD��-�(�0����N)����-D	���z��ϭ'v���<�qIy��QW����M��7F�s3�{Pk?��7vf_�5͛��h�h�h>��<�ŉ�k��M�I����o9���=P�t>E�����јh�H�w�`�[`ŵϩ��\��v�f�.P�J��`�y�{����3�`ef�Ӣ��ZC�N����L���4%��^���e嗣�εsϰ��V��E�r�g�\meS<�'6�*�1ESU�0F/�l;T�F��j�M�v?"��UZ:����(�4+�=�׼������%%|ib��@֏�����������؃֑Ε2{�T5+�� ���FI���z�)�h��4�+.?b����>��r��8��۫u:�ό\��0C3S_-T�F��G��.>�!�O	�-˄�7�y�}Y�u��\죴����~>VZ�׵$�B��=��S9�S�p��O떩c梅�$3I�N�%�����8����kt2���-{3[���GE�2��ӇlS�����C���ˮ��s�+3��u���Mx"q`�N��ɗ���j���[��w��b�d�s���j$û�����Inڪ��}��d 1�����O���(�}?.�V7�`���̑K˼�����?wW�)����5��x�2	}�+eu_�R�+Z��X�~�T��/�|1Տc@��M��U�x^ȍpo�7�\kC+Jta������5�A��DN�7����f����X�xY9�(�eK�ѿ�fo���ovD��BF�����.!�Љ����(3G�Ù��f���'E���^��I��\��o	i�F0ڽ�*��-�+�
HeӴ���t������$����|���-�-����z1�z�\*��S��Ŏ�O[=��5����K2����ՠ���R ��z���V"�o����e�Z5��@E��&���)~�-���L��Qy�RRӹa��F��d5�B���`��i_�vl]"rPT�<��^�7�g/��{V�4K�FR��k/V���<h�^��Em/�*m��V�H�9�r*��$4�i�����xԇ����k@�QOzK��lؤ��JAǣ[nP�B��3ܓَ���zg9rgJ����(�B6�����&��J9g:`�/:�e��� T����������?��<����C���Lު��!r�s�������=��$���`�c�*�ٚuPP�vBvI8�x���!����C�����Gov��`�%�U�U����a��a���'�e�,-����{n|>sV�^��W�}ғ����W}b�ag���}��ԓ9%�;"\K|�H"�,,8On�$�^��;���8��f\�_BM3e�ҵ1�f�>�S��>.Px@�~x�}}?`�^�{������D�_�~5���\���bf,�:�,:�}����K�Y��?�毞��-ĩ�؊
$Q��)���x6\?�8W���z��Y��*���y��9�˅�u������e�`ҙ�ZX��6�����2�2��-{��^��5�o�lRH�y��Qnc�S�!�����ڛ��}¼h�	��a���!���W�=.c�a�I��������^o�/j)�gj�E,aEL�_W�V���sWhCɵ�R��2�O�`=$��c{������V����V��'.��J;�z������}�>9k����F3KS+�MZ�=���<邺��1\���ș��"B�a��Ǯ�C���)X��<�PG�D�<�`t`i̜ڻo��-Ȯ�G�_ݱR�rO3�>��؟6��9W�E����͎���wmͤ&�(a~T���}l^} 32�,Oݰ�����؅-7(X0܌�ۜ8�Վ��r��X�؊�(fç]xB��������C܍�\Є��Xw�7�yw�g�w��|Œ�e��^���X�&���@�� �/�����C�)ф�i������V��amo��]�S2�Y�=L���b�t���Tf>��U���(r=]!�����w�ѳ5,���;oG�YXjv�G�����ly���`58ٝ;�f|�Fh�@*�!u�Sz�lT��y(�=�,�<�GD5�r�&D,�����\9"����.�|�-ԃy���6~�S{��|jsg09�(��7�e�9���n�o7���i*T^����%C[�'[�"��"�+a�y��`�?���F�IU�ŀoDƼ���#-��9�����Δ�����d	���y'�.�BY�=��)rR���g�E8��<��SR�KQ/�Nu�YM�S�˝�h�#����C����z�P�~��!��jl�l���"/W�a�dq�wX�s���v1�$
"n@am�I��=.����Ƅfb0��j>�`��dL&��{,���e�=Ҹ"ەM�W��]�����A8=��(j	&�9����,����]8�Q���j:�)悬f ��L�m�����V����/�8	
ǜf`�ɱ>��W�*�4�B�9I��q�FCPP;���H�H���oSÅ �˰�Jc�j�=S���w˶�҈S��g}7O")T"�)W�h!�*�x�)�^K�W�}9��Ti��RԨG?*���]��)C������8�R3��;��u��z�Ó�@h/#��)/��'t�x�\�h�=(�-�j�R��j��C�z�]R���^��e]�1II$��~-yb�_���/��:A>����$X�Ć���Ψ.����&�(�C'ߞ�ue���>"Ux�$f��K��&Bt�`�<f��ȃ�����'���tIhu�f;����͌б���9v����/c^��$6��HV}�@ԗJW���}z!����MƠ�����؅��8;�ll1�r���M
!��⟌�6�s���r{�X^ăi���z�h֤Q��$V��>��� $j)�M��;p\/�}�92l��{���ݱ���R�Ĳlh�g�9a�(זL�дm��a���*\�k+��ʨ����2oX����
D'�݋ޛ"W��9\ې�P��tNͥ��s��ɰ��|�w/�?5��Ȱύ�-wwH5�e��0T�~�/��Hj}�!�l����$O��R�#������rv��Bf���Q�ӳ!���p�����S�	��Wo%c]�@�7+�B�S�BQ����Ds����Y��Q�<�Ǧ�%4k�V��@�1hć{W#��4��T������TD~d����a}s�j"Ԕ�Ԅ���Z����*�k���}�d&�����&O��W{le{�0��؏6��"j�0�%Ov��Px�T5~�)"��!�����x�E�8��||�v%ZI��% 1Hx�?����C�*���|�6
X�B��Hq���nU� %��̞5�2wڷ�bSۤ��w;��c�ǚ�|�j�u�ѧ	�?o�D3�m�{�TmJ
cZ4�"�x�\����v���,:�����O�rp6�?$c�|���3��7�A���
�X��K��N���HG6kP�O%rWp]ѿ��P�M�,뤢��řxɎUO��n/�	//q�]���at���8�+����JE�ǀ��ZS#��0޴jC����\��̿�͡�a�p�T���Ddg��{	(� �H 74Eh�6�����>�$��=N����a���W�-6CR\�g3��Xzp�?GxXML}��=*x)7��F��%ˮg��� ���k��Ӻ<t<�t���
�@uRg�|���Q����������=��T���7a�����{�Y~P��OLcQ�J�x���K��hL�λ�� >�`]M�_���2}a��ɗ�����s��A3"n!`_��o8���!���+"\s<����@�r�,�+Ә�t��*�z�E�rl�������ۍ���ש7SL	PP�)L�	b����ig0�������J ��Ƣ� Z���S���)���"�9���1R��q��<-��W��돲�j�$���o���Y9�/�L@�)�a���s�Cw�'>(�j�Э {o��� �%6H:E��n��	Iz��]D�;��Z���N���睰t�Қ���{��!���$K~s��O�l�����w��RN�{C��u_t��p\D�7�y�䟷�w�Î%��9���(6�{���w&�4��d�?Ѥ�/�V��Y��+D6��8¨�������v��n�ܵ����w6�����'�����[7�y������Z����j;���j9�]�%��+i)��a5�=vJ��q$��]E�_����g�,;~̥�iJ�K9ܰ�������Gb>�g6�W�#�`0��w���Ha��Js�X��+�i_�n��}���ڱ��)o��@C>uGVs��)yx{@6X��W!O�H������)Y9���v^F�Ґ�`�*�����jAO#��9�aS�oh��`q��O-�_*����,�b!��([��ڙ�D�5F����|��^w$��e��|�5VCz5ht.�����6������X[ggS�`�}����6&)4������21�����y펐Ϗ�X�G��6׬���=B�V4t��}F���z�B1ցyF�qZ�

:��y�f�նJ,L_@�O8����Ξ�.T`psW��.����Bn�p�lr� �%#��.�S��%�ר��므:�:��1�ąE#'c3����6%pX�� N�2�.Z��W$��51�� ˎF���́��?�5]c�0�O�[�U�
D����E�BU&䇮'�z�x����*q=�Ye�xgߵ�0%s��U{˖�n�e���?.�_&k��;Hk�s��/�o�50�d��Er{�{ W������� <h���<��H`ʕe��%}:|P8*pˑӑ��.��N
�e�v���ݸwK¯�N�ύy+&�����%h��ѐ�����E��R�]<nM{�[�P�<�0پ�}�1jͮ+�^���EL��Q�B�\����(�
h)/�+��wia�)l��cM��}��
�K䑬
[�֕�L0��1e�E�.��]Rj�A�,
Kgް�mv~-'�!�����to�VӰ3�7�V"�eC�	+>�c�9#�AB/��sF�ͪ%�L��V(	����v�;��e
�bxn*?DMɁ��C�8%{�P=�c���
��!�Y����l��7c5C�}2|�8k�������a��{P b,h����s�t"r�EU�(	�AӴ�2����ƥV����iV���V##	�Sm�XOC���V����t�m���.�N�%��C�������9�����njR�نD8��i_�2?x��[�&b[��◍�)o��E���]��E7-;(�r�O=BKvBC"[ɷ���݆��j���IXs�%�ĭ���jSF?���d�h�4�2P2�}ǈ��������R�rg�y��ZD1WK���#��OE��ZSC����G�)�Y���vq���Ǌ"�����x�� 7_���28�߈}��U���������.\j«?����_ҏ���߰scW4 K�`�+-�mf �~��yGq=�M��U�jhX #�6>�������J��0H�4#7h��r>(菳���PYg���8J}bX��L�筹IDs��f��˄z2)d@�������.�.�z ���2��E񤺔�A:)v��@{�M�&����e|ߎ��6���$�$"�)�]J�ox��͚�	B��/�w!�u�9@���	�Y�ό���q�(��%	j�}`�vxw�L�v]��S ($ukj�sd�+�(���﹆�e���z���������>[y�s�D���U)Yy`�	Ѝ���뭖�R�uoA˕@/�qk��Ba�a##��~]���}O�g��1���ݖ�$��sY�;U�E�R��ۏ� �"�i [�o��E �}����_T>���/�K�v�	�����������z��cQ_/$ZQ����\���8�!�y3Nn7_QfObBײe(^���m�/����&�L#�0�NM��z�M-T2� 8f�>�v��u�������8-}��������%��h���S�jZ
��@��x4H|����� ��t6���/*WX���
<�I
f�ܣ^9�Xf�8K!��|�euF�),���D�����7�M�t�d(%�H��$�޽dݧ�T���ۑ]|	���ah�"b�5�n��į����WW�J'�]#Oc�k7#v�w�i�lJ��Wp�L#��#��X����l���,صi�|�m@^��((��.�Nk֮8G~��n��#�KH�����m�<j$,'���
-�� ����6^�F����`�y_˸(�9��	K���@�1�d�hz�pd�>s��͜��KWX����'����>�����Ӭ=b�1�/~�SY�[@lur\_P��T���y���lg�
�K
C�q��{��f�hF a�G`��Z����C��g-��1o囼��������U�bԙ�'a��:�I �H�z����B��C�o*`~}"}g_e%��"� ��#�zʉ�+tƉ��<��o��)�Ɉ���3a���P�J�L��KJ����z���36�e`��{pK����9j�h�v���@!y�;�h7��8���-�[�%_'D��ŗ�'�W��5�m���'���!�@���5�9�C�Re]��*o�6+z����˖�3�n���U\�>�-i.댨�Ӻ�x
l�����L��|Ѥ1�ݞb�:2VHگ��P�Q���o�w�G�
$+_j���A���QP��B���0�=��;���]�ݍ���+9+	�������*��e���྿N�%ԃ���zY�kc9�e41/N�{�^7����.MlV�:��@es����W΢I���J��s�Z��vx�g��@��B����2s�!1��m���=����2�-W>�p
��ލ�n=�ԃ�aḌܴ{��|����:Nz�:����N;���Ţ�l5a������>����=��U|<Pw� 	X=�{=�β��r1�b�G�a���\p~���{f(������x�M�.�DW�?@VA�,�El�����e�/X��K��@U(w^շ>�C Qs&�'���(Hbب	 紓�
��5n�I�VJ@-*�6��{l���942Q��L�3�u���J/=S���G]�?�	F�}`�����Q �ֺ�
Ҋ��Yd��+�0&t��v��D�zT�˲�P�V|i�w���Ux^��}j[����
a���as���HfLlf��L��B�t�J�ߐ��5>��+_-,Z*SW���'�&Tj���wJDS�g�iDE���[�+z|����YLr��wzR�.�V����T�=�1�qo�V�U62[@�����5Za��q\��G����^�7����n��,Pe%Q��ݰ��ń>�r��I�-�{l���D�8��ֆ�MzJ�è�-LL��j`���mB����x�8r��u����L"a��)�#��^���������Gk�R}�}�W���[�[`i�pbCN0L)� #bw� 2���ޫ.�g]��"�ı
e�;仛�İ%W֬q��8�ł`�ef�׿�p���:$��w��d��<��6��t��H�O�ε��w�<]�`?��l�Ty����+y�,�o	Eq΃P��OD�p�1K�:����ݤ7E�p6B;ڻ�]�Y���l�'M}��b.x��-��Y���30��oL.W�B&m��?��/ٴ��z'e�0^<�z9���֓��n,ĥ�u�F�%Jc�`���;b,c
Fۧw�c����b�f �[�"���v>ⅈ��tz)��1]��-$��kD�ʛ|����,5��s���K�,�8;�_ت_@~�4�⺀4Do`x��Ԏ|R"�4"��� ��oP�/w�\�o���S����D|x��v���0�18A{/v�uv��[�su)�y�(]����Vއ�5��IԼ.c�f�Ҽ-~W�������V6��8q�d��&���a8�����O���:)�������K]��K䌘�0�s#v�G�7�8��%PQ FN���X���j>���Q��x��Z9
�̶�M�կY�*��D����8�4}���Ǻ��`����
�����b���Y��j���K��i��wK���%9�2n�P�-Fa��[ ��s�hwꃪa��<�S�C� ��W����1`����b���8��}�Jf���pM��HF����Ti��E�Z�n+������/m/��/�{3i}�k��2��\�|��]���#X�x��ً�$�xDƩ�f,��C�S�1^��{�T��ֽ� 0u!??�f���Τ����s�E^����=�]"fc
�5k�����1�(̈́�	�o���l#�ѸY�*�yjOu>i�x~�6|d��Z�}��R�qp�Oo�7-&��*����ڋ0�UG}k}J���)��z�������Gl�Ύ,a�u'�*�a�;��o��.�=W/��7H��Z�2����E �=�[�_ԙ�b�d嶟�����B/N��u��Z�<���58�d�哀�"��\ɖ�:��e�݆�r��5�F��_ ��׺<+��q��/���}sFY��@�����ldm���{�h�$RJ��X�y|�<����ڕ�z��d�hOKQ���{�����%��T~}���̠�'tT�T')�ض���>r��AQ�}�$��3�o@<�t)�47f����o7o�W�x�o�Ǧ�$�W¥�1��`�/��lM��v�����*B*�LUz��*e����<5M<���S܀&}��i�-���?�8V��mxkmf�8+R�����H�Z�ky�b�g2�kӛ���P���5�,b�}�F�( �_�k{�߿�y��RU�.IE���[R}ͷ���Q���~��|�کFֹ6a�+[|z<�[���L��Kiw�h�㼝��O��3���^{���B?y�~��y��e�5��v����=�;�9-�����B.��"y���;�����x�z�͵�f>D���>���5+pn,/�~�?����1�IH��||�M����x<N�<Q��($�]V;�h�񕑑��G��>�v����ͬ�b��>{f暠5��c�������%X5��K�e"ȥ��s�*�:7��~�k(̃x�فt�I�į�R
4�j{���,��(��,�����>Ǧ�\1���n�W�X��#�q��:����T�Jl�qH�4�}T�+���Q;O���tRcM�`�>�l��^��@�g!(k��|S�4��o8�v�T�B5�f6����l�"=�@���:�����`eQ�3t�\<�s�v@�2�faA�3'U������R5�Y����"[�0S�>ty4mV�~�Q��S#�M�,hZ�-ㅈ����o��G�)�>�=��ڀT�@�6��߃w��&'��!�5�J ��k<��4����(,C�	t��'X(Z�c�ʢV!���㿟ܨ�Ȉ���U��+����K������UΓ������)f���=���6�XC�<���'0T�T����F�V
Q.Ӌ�ȃ�I��%K�S�5v���P�����b6&�������):`���'!����0�k�d�,������c���&	��\A܀2�Ȧy�W��dը;$ɳ�e�����rx^�V�dݱb�?�!�Hg	�d��uCZ��qnUr�
l3��.����C<��-��"�#=khr�RZ�F��}��N����[�gfn��puksW(�E��~�O��v���ƥX��t�t���o�2�u��6�_�a���n	Hꄵ�kZ��zaο���݈��H�:n.]B��~p���xA)�aT!�(|��"d��۽N���������ĦkW`em�ϗ�(����$����۾�ء�ś�Xp���Z��9��d��&���>WU�����iF�1��u���lE�K�;�nf}h��m\� уM
��0����BGa�~ق�A�� x�=E���M��̎�Wa�%�z�܆�E+<@h��.9�>HU8@Q�|�i�ˀ�+�A8w�U^|��:��J��wD�ON�]�H�)Zlkh\�Y���� t�dg��`��������-+�˻����{�Љ�&ɵ��*�=�",�9��>��Ń��b�3wg4��Z�3C��pl^	)*'l�[^kX�[��CXS5���T@�i���o�˶l�h��CMs3�z�xjCǔ����EFR�%^*���5yV��^�n���ƚ�Vޗj�gsC,�F6�I4�;�v����ʝ/Ϻ�m�y�Y��(�+��\*JR��+U�	sP�Q������a���\�J� ��\�6H�.�����?��@-˶BؔA�l<7�^O��/�ON�ֻ�Y���\��� ���!��~��'#m�XŮC��bLn�k�A���6��p��eNO�(\}YkFj�k�lݙj+�C �ߙ����Y�w���Һ2�?h��oU���k������ET=�X7l�p��V �Ը������S��Wc�H����W��x����-4F����;��؇�_���zZ��h6i]���Ǟ��q�F�K[���{������l;7�)���UC�AÂ/�Xi�l1`A�9E�!݉>�W����}�˻(�4���k抲�T�!�m*W��	{�|��$����vR�O'%cu�����Hs�o`��U�eJ�P��yЃ���B
��Ǉ٧
���6�Jz����LN/E���������a���K� �#� m�d�����f��(x4�����ޕ�j=�k���i!s��,���y�_:���=����ђH�>��衤A�pI�����F �g��DΉ�..	I���(横�]j���SKLe@bL6�݂t|ŀ��� 1�K�(��e^J�,5�Xj�׆�W%�]��k�&����n��-�s7��O��˦��[�'�;��c�12��E-���s2ޭ
��3�_�p�X�t
�R+��0�kD#�cտ�3�jk�f�djB������^�u��a�nW�#��Lo/#�/���@������?|��uۉ5��4���b�n��ȸ���
W�@H(� �?�0�Z�+׽J��h����I����N��Ǚ��kŔˢ�,I����#�\���Ew�[�k���>�����Ad6`v�Vc�ˎ�u��N���#EG�^�U��GT8���~���ޘ��U�޿��0�X�j��0��֑|���/���`#�ĺ����v��9$�P�mH��v�*6�׶N�do���L��!)f�虓2"��wH����>fL�b2��s��&}�!�o�N�yW	��7$�V` '�Q0������"��m;K���`#n��tIs��9X$���
��jZ"}���գyx�����IF��a������� ��͙܇M^F�A:Mg��k3T��5�9h�߯?̉�W�V��7#O
h�|ߞVDb-��愭P8��Je��]���M�'�_���0]x��A�!|��Pvw�l���s� �µQ
8aP�猀�)lC�����2�gKU^��QjR�2w_�t"��0sx~�Y��C(O��ԖW�3��߬���y��@���*��W��X)�4l|[m�e�3��P`�]�!����"~�1�����7������\�(�$�7�j���Y�$�ln���{�VD������W«�q��N���:�'k�:Nx�:vǟ���<�)'9sj�d^b�2�	��X&C��D�ŭ�G>�g��!�����!&7`�cw�EjL}��|HT-�)l�dB���E]���%�N�L�}'>�iR&����O�%��/O�>֐hPw��ʆ [�G�ii��עֳ�7/��Sq���ʱ4)e���9�S�4�&��9����+�³i.%����ω���1���IWu;�����V�,8�psz�)��ă+}X���<��{42�M-6�,�j�<R܈a�j�d¥�����Y���նv�g�(�b<u�J[;��n+҃���,���11ب����J�T��YR?���I��jVE��&|Wߺ��<��l��Ua2�b݅��\u�SB�V����7��v^?^�:�e�H�M��A�N"�W�F7��:���Ʊ���{>�.��j������$-h�J���� J�D���Р�+u�0u ��4�&D�\�c��ٓ銷�G���;�.�ڀڒ�t�I�̷.�����cm?��\[��}�m�n4�n�7|[S�
L�;��˰ʝ�]��S@T,t���1��&K`���T�C�V���'\~�X+SF���p�5�d�/���%���s�|���B���^u`�3C\A���K,yACD/�.�҃�a[�Lh�=!����!��(�&��i�/��'WW�;��>���X���y�X���g
��3cl�s��3!�ژg
)�5{s�j�싯�D0�7��'�f�x����c&�B�{�.���c
�Ż9�����B��Dq�t?�����`�z�@�+,��@�����B�ȡ\!��u�=��u<��&&R �Q�+���ȷ��Gʊt{�/HT�e%�ߺ�	��}�=��ų�2�BxAE��Ϊ�ϺI%����z>q��f���`���(����`i��9[&�Y�̇��Ī�5�ps����&��r�Wձ�m�2�V]�Uo͕r�y�tC3�^�)$!ko��Zc�h�ɨ����-�§��69Z��1�f��a��M��3�NE��z�0��E��f��R��o�l����� ��r4 4��2*�9/��ل!	L(��teo�x�ZC��퀜�w�|����"��r#�ڊ=�+�T�]e:r둠��������9��X4)+J����̇�~v�k`���!8���q]��sδY҄X{Y�Mr��j5k���RĒ��),��r��(4M��H%�%(�qs��ܿ�~<���5��
2������M�и�D+���Z|dm%�2K���/?�Z-���6=#�]Y�i�]���s��)v�z��3��شYR��t��I��0L��k�W�1���8(��A��(��-�����F�sۿ[�
&�χ��j
	�9��&����`k�jujQ�U"D�����#�-�+�G��HA<zW2ItJ���tKd��xim��f��n�l@�bhr��j��|����<�A�&������m�y��'N`n'W�f���O�M��}�T�̑c�Ͼ�F��5��I��6ܔ���B�6���f`�_e�����m�4�7��܆�
}�{��"���� 0�T�=\Y���A��Ң5w�R�/!��p�#� �W�}y�϶4S�)�D/L"��A����=���b=ư	UH�$�{���{v�t��������l�p�kF�/+�Bbz�&6Aj�������"�%'̼\�����"����!�p�'%�~24,`R���Ȩշ��+;U�����ђ��ׇ��}`�>�P5�l���������"d#v��պ�:��68��
��o}�⊱���l<�_78�ъ*��������k��~S�a�(�?�eb�VeA��Ϫ.�5l-��o���]�q���z7�0n���:6�9��Q�濘{�K?	5�n�1�޸��KAe^�H��Gh�ӕU��b�0~����;f�^��v9�Ą<�+K�<P����и\h���X�GHk�ʆD1�g��iA��@���αѰ�Qi�2����K�������Q(N$���n���
���7��������rs������Tݚ�R�3Yw	� C#��@Vo�V ����%�u���;c(�ߞ������������V�X�� ����Uӱ#M����\�`����}(�~摕^%W��$5�
֋��� !P�'������`^�*4������s�f�:ڈx�B}�l��� '�4"���+H��n����DᑂX�Y��𦄩��^���gH���.�|�È2�)�<Y���9���0j�d����1��u�k`�{�x�_�F����E���R ~����L���k�9ݧ4ډZ����MS��9�m
��n����]�>��}�x;�*�iľl� L�񨠯�Kqݠ�yHF������H|����g+;���wK��F��j�) ��6׮�BVIu."e-٦@�O�S�0M�o�©+4�fچ������ {;Z�r1���Ҋ�V/03 +�z��H���7��j}��q�Q<�52lx& ��^g�Hܢ��+�̨��V!IeϡU���V���.�����a�Z�6
-��>��K^N�<�4����Ƚ���]��S��E�� ZpR�#��P$g���yGH���\l��w٢�����U	u��ٵ�%��p���u�����	��ƀsFv_�me
V�ӹ�~�~����̙�)B8v�y$pB�@]�J�P7��6u�SC�qh��ҳ��i�\�٥����A%����T���)E�7M� �!/��R�}�S9Z��AH[ϑ�g� P���@]�1O6u�KM��xza�8�o,�{#�gq{ݙ��g���� Y��wJ�%/?�GBFz�ynDG�8�ng�C&H_;wYyA�r4y��ڞN�7b'����/���g��b��/��&�I��)=���1��D���q�yp�^������& �l~�;ń
*w&!-�L=�_%KxsM��}�.�~Z�7�1x�C�2W� �I'�g4+!9F�b�B���FדtiE��u�i���}�� �Ţ��
�*�W������P���R��J`���h�0������9m]�Y잙���I}�:ף�	�
P��&��(��V��3�<oCB�H�B~J�.�]uz�4t��o�p����P���ȓE	*F��<��8L�����f�9�<�S@*�%LY��]Cn�}�����U��Rp@�yvtswéP��G]�@	�7�D��9U7V~�A|\(���@$f��%@�ݨ��@����QD�0�FB<�:�-�i�9����~��*����%�����jp�뜌ҙ�p��(gW/�pk}q��\��
S��B��d��݅eҍ@�kEL䪄g< �È��Q>��^�o��"�C�����͛��j���z�� 1�o:z4w�ϼ
#�N��
Zl���	�0wFe��̃B���Po�9�V|�[{_�]���;��&H=�ό�U�\ސ2<n�RK�ְ��y�@�O�ѬMn$#^Ϗ��_��קZ���1���Z=�u��!2j$���{���Z������lu�/��}��ǋ��C���%3�ݪ��j�FF:�;
�Os� �N�n�<m�n������,e��#S[�/נ_iX�,xiJO�M'Iִ�Rz���}��2�:'C�bi-HfX��R�ݫ��ŭ�&�| 