��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&�����6u��%�R�l���ɒ�[������ e��4t{O*&�z"iM���z�� _��)X;�g�(������<W�;1�g� ĄY�;�MI�u\�Ĥ�P�њ��P�8��ڙzd��<�<�\(�*w���H"Z;#Uldi��N�]�J/��d63��Җ�H4��%� 3����W�U�s��V��g����i�W�~���1�c��*M��	`���\~z����T�Ut5�&�rryo��R[���&��3�� Ɖ�C���^X��{�a��'�f�Y�.��_�Һ��lL^��6+��q}�V�B�?3��-54�0+���b*���%���u�L^C�(��nQGz�c��W%�:���!�����@�d��v?s`�^��k[����پ<��z��#%���g=���@y�bь*Ҷ��
q���D��[��N�K��,l�I�7-1<��%����M���Օj��>�uP��j&��:�҉��Ϩ��;�A��#�ӃY��p���'B4}񪳥u�Nꕵ�՝�5߻\���E��q�I-��D��?���y������;�U��4G�*��y*mp�2�R	�a̶)�_�J�d�9F�t�9����P ���Qwz��NQ�{��;iw��0����i; &	%��|�2����-\Z����'M��EDSO�����}�	��a���%���K�
�k4�޶��R�`�*Ga��=t��]�
�	�B���kUS�:W~;�8I���G��t��F�٫��?����2|��/̈i̐��4]�!�!��P�4o��^C�f梡m»Ua$ @	�F��͇Bʳ��<3hE����QS��D����N�L0=G�N�'��v�<=�tH����gk�R ��Q*���M������z�t��#H}�3�	V��a(�)G�����_ �N���p����Q���4�=�5�n���w9���ISܳ�e�D��ӧ��@�{�mw?%5���a]��D���$�9��3�jaJ�%�ųA�����^lK�*�{��e�����nК!AƇ���+T���Z c@E�1S�[��i@z���4�+D�0�s���>k�Jng4)F�f������W��v`1�O�:���&��ǼX#����Z��⛪�&�b�#TE����%&O	aT$�fS<�M�&;�Ks:C�ׇp,�6���޿����Ԕ�� ��!]�����<)-�!˜� i��Y3��S�Լ�~��	�;�۽����YO.0ɶB}��X'���b��h���J�q��o'C�Ҡ+J9I�4
N�ſ����x]�$��Nڶ1����[�KT8�#G�u$��MC���(v����܏���HY\*�;g�Ԛ�L��*��2�K�V)�"\��,6�\S�RYc=ؤ$���k��^q�4�t-��d���l8��֦݊+1��W#�3�D��� 
��<�ZH���f=���C>.Ks�#ۗ���jtH]�l�j��uY^(Z���2D"wMW"�|F"�c�n��<���Wa��¥D��aJ5o[x�R.�EL��' ���|N��h��v7���{��lzj-��cq�w+OL�k��i&���%I�N�/��� ,�2\CI��n6����_(9�m�U�Dh���oU�����,�5J���/�^��zrbj8�u�b�=ц� ������l��+���_oN`׎}���͗L#oFEX��� 
w�'��x8/���#��~FnY�:ޚ�z�v�s6mwЯ�u��Bhx���A�2h+)8;]7f����l���%?Yɫ��c���m���UѺ �b�_ڛ�}�A�
������ʞ�f=��	�e��w�W�젦���?"r����qΕ)��N��=�:�e'�ߟp޸?ṭ����2w�x�O�=YG?�^����
�D"�� \�������>���o��aK|�aET
�����]���p�k�0rέ�@m����>�~�&��${�"�z�WaǑ�\��犔3��I�D�"���=�w�KnA�8b�SCY*�DU[���et�{�績����>���m�<v��:�*��<>S8����g��Z�{�5�@�4�rxoM��T�����Es$B�3�,�)�2-�+3��#����s&���E�l<=#7X
�gf7Gִk\#��i�ZtG	���pm����󌥊!t*�`��QW��y5�C@��<��x�<��ﯡJ��=t&����3o�Ѻ�:�%�NW32%����r�9��w��!>A�?ⶠ��.��.�*�#������!̅�w)h���ޡɊp�<�;��IN$�uz�q��X�P5Ԓà�:,<��+L�$�{�1�#�0��w����D��P�i��R9t���jl������ip��m�$�G����\��Z�p�&'��Tdx��`�`��#�l���vZ�R6p�ݭ�����a�_�+Q�� C">ߑ2 �=(���ڈ9>���c���xۣ���~^ʖz�����D��oW65��C3�jb�<f����Pn�'�`���q�@tL։�
=���W�+������/:R�3�D�O����S�W� ��5���b� 9�O�UM��]��@�w�8,�3^�V�mzժ�4$[du���3�'%�9h? t)��������&�ۖ�l.H�U�lM�s�޿�e�V@��<���Z�B�e֔[+B������t�u�&A��Vf�3��h�$��:�Tפ%%< �d=��Si�ǰJ��h�\8شѪ�#�S�O�ؤ?	o#��m��kOM�Wmʶ�	�C�	oD�;.�vB�~*�?��1�ڃ1ۡ<0�q��j,Jq�x���e���{pUgq�{��P�&�h<W�㟯~u��'x����5�7.���|���~635����%���Kv.��Py%Z�i���&����j�V3=4�P;������5�~ۑB����$1��P��e;�O�^x��JV�pټ
��ά���|������1=�F����pԵk�@�s^�~	׹/�p�,�w���ξ�����y���!iY�73N 3�^���j:�(�_�$���`������4�B?�����~��0]��'��~�Xs���JIZY(���g�)�N��R!Y�~��Դ�CP����P�ǂ���e,��E[!s��ݝ���0i��1�l��m�6)R��Q����ʯ~�xI��s@���ǋIэ��L���<bEV��dBs�,5J�ļ��?i�Z�E��T��Z��������&�|���يSAٲ�pBb)��!������)ɼ��ѼK%�ײf�*Yh?��ۋ��m�j%d;��$��A�9
�ql(T��d�������,o�y�O�m�R�3g	����bE�;2B^���mex�?&��gv�O���}�h�֫�����ȓU���f{ҷYL~���|�Tt����Rd߫��Ό�7��ɢ��H�������h�����^߲SC>`�~n��)��@��KS�+���{�l-�@�x������rI�Z�]��զs\�����NH@�D��B~���\����\?�SNxK���\{�1���M��&�n�"ߘ=���E��J���!�k�I�f�eC��qL�+j�KZl��[4޷x4	��n�q�k�e(�����3H�O61]�A��1h<��T�^�y��z�2�Ow���n�k愆���Ӄ�Քܽ��1��I�R��̋���I� �}�C��EiY@7��bǷ�r!z�U�hw�Q�#��z����Bϒ�=;5�EmR�%��j'�:�ѽ�;����e;6����U!~���r��{ۊSL�H��zZ��L�t,��%�>(�Gi )4��>>7�Q��6�����ӜhZ1I�pz�v4y0�71�Aܢ�ӻF��^#�����k�2�"œ�����{֚���>z��W
o5ֵ�6�fro������I;������yj[����.��8~η<%b�%Bz?%�ŗD��c�2����������	&�E
��@���)$m�����hq�ȃ�����f!�m����2�l�tc�\�*�`�דZ�ISV(��9���f{�1h��]=���$�&����l���w�7����6��S��<�	�Վ�󽨎dt��d��[�q��_%�)��n�0�,���o޿��5?��'�:]��-e�|���T���]�/)s�,��$.U���&��F{]1��Z��yǣ�C�%إ�:�e�wJ���'�?�I��U�����p��z�>T�<&f)��il�>�'�¥N���G�P��6��X
O��M?���U�+�����_�|^��I�e��}��謫k�#�o�^�HUZ�{�p��O��PyҰII�W�J�ՇY���[�<t��h�g6����D��x����W�3�o%b��7�	y�bE�E� Q�Z:�ml��L�bV�s�v["���_�����?�J�3�ۭ*)��۰_;n��8������Io��?&�x������~��AVI�yЭa����% L;����fAG��������w������9�_2���d���!����c��j�j{�]�:���e���F�&�D(�O)Q�QJ��UA�h�	j�����ĺ�$M
�vx��� ~~�2{!#e��3�����L�E���,��&�xNln��ye��L5/�s�m{>�V`Q~�I�	��d�6�y����}�3ZKBQkp��q�g��D��R3���hj���Zz��qõ�$5kS���[�wۗ\�����`A��蛀����R�༩c� ;p��|%`$`6T��ä��t��/<����#3&����@��͟_ù�%�O��:����ot!�۝3u��ci���0���4�Dvэ�JJ�����c.:P_.�o��I�d�����>ZҰ��O9�x��I�j��M���>8W�1�����w5��x
lt���ʈVaЩ��<[�{��{<]�r5c��ل�6�_���d-�I�NQ�>�6�+D��F�h���fMkя�ƶ���]�>iY�d�`Ӓ
��ȗ�T{U�Q�e�k:�o#��T�U\���i	��kTȼa�*�8��>^�5���|+;UxW1Ϭ���}84�uW�Pɇ�2����3Sf��m�7���c�؉!'D'�9�22���W�iCM��/v���d���1u�Dn����s-_�L崛����T:R�BA"Ͳ�����"�:�O�9g}M|�M{Xwѓ��Sr�UnA�ԸW?�����;���J�<�=۫�,����$�?̱���3�U^��6��de8=&:��D��J3�����p�"S
.T�����e���nd��¯�Ǥ�v�&������ƅN�	�m��{�͙w
 sl�67_�>�t�&a8�����B�4:�NАw�7Jx�@D�-J=#y�9�V<w� ��
�<��HNј{�l��m��-<��� �f�����éL�̩M�f����v���=�J�.�W~��48�����O�dv�\8�%�{�ǃPWİ�G�:Gj�?
��"
���ˀ	o�z��ڗK'Kj�Ota�r���zT����	�C��S*K��!>�vG*hH��>,U�� (S|��w����[|�C��IJ�NaNmu���{��)cZk��� U�ˌsNH��k(�<��xaW�w��0��� Bp3�1�D#ig����DF&��w~5$ �Y����\�[
�KSf��JM����b������s��l\�8k�aT<�e2Jƀ�y4�/e���r[������I�5�`�ڏ����/��0����9��e_
�"��Q������/�é��ʑZ��.tz��r[1H�@gf���r�L�6v��	�~kv���![+K��OLd}��gv�T�;�Z�ـe�C�p;�ĽM�2��f�V���t�qG$�}~Z�����ny����.+f�����V"�tGxz�U��ܮ�>�B�����b�R�)�ӿ�<��o�&`��=7$��Q�$�T�y�QȺb)��W�`c����D�8�6F��+"�Isz�S��c
E��&2��T��d���TBo͆I� Hy�jaO�0}l���@P��Vw�iԐ���x�c�R-�Q��Qb�����i��ɻ���l72P� �,�.-Aq���6�����a�/�����R2�[Ÿ*a��9��@w\�i�pM8JZ�s�+w��<z!�e�.Hi�1B����Y��M<�%P�*a$:"M�lY�Q�n$��Q����me\�<|�b�ӦG��_��|^Yzg�AM�h�O��a��%��2����Gnv��kvr�=�.a|�?�I�
���ah�;��Ů�C]_@u�S�[�'��7~x�m0�/�~��ˏ��a:��m�\��G��oL�����-�p[��?�i�sUƌ�F�F���5��I�v/N�%@R�] 
�AK�U���C^��(����ۣe�xL�I ӌ��~���o�y�X���'u*�C
uf�^nA㭇�I���ʬ��f"Cѭ�r��C�N�;6�5.�p��N�'�����Md�|�s�G� L f3��rI��p����b�!xM�̂��!t�49�i!��(d����WU�,�$�I�᪀s:c��Σ�ڮ-B�74�p�dp����&�_rꔮ�o�6��Z��J�+?���5��I�@C���ξM3���_ȶl0 cg怟�\Z��/*ܣ��a�I��((&ʣeh_����D�-�:�h��=��o��ِЙ��N�۪D���9���Z"W30y�2�R�t�@��z��������>�c�/�Ɖ���ډsbr���_����.;D� :���mp�'�g�^XQ����-�v���_�z�?��4��(�n=xI/��rJ���	(O4�S~@7��/���b�z�_1i��K�е1I�W<_,�L�2?CO�JX�Y�$-͵��l��k ]�7<��J3�m��]ً�������nT] �
|k�b�rf��Xgm��Ǥ����W'��~`�Ha�mj��c'�?�q���A�*�n�o	KЅd��X�T[�yP��ʷr���֠5q�F�'���)^�=���k�W.��x�zKC���*TM�Z�%8�H�Y�mb��AotMF%���"�	��?����jt��fc��n�U�@�P�$���o�-V�����r��wDl.��-�w���V"[��	��u�ņD^)�}�2>5�����������nH�+x�!�O��9�V�w��U���� 9.9w���W��3Uƚ�+F�\�ׁiMҲp8��ՅO8���g 7�ֹ���v��|�5*#vIf�{d�����nI?��ߤ�����)lٯ�J��sǱ��E'���j��In�[{,2�h�����bY(͛R�d��ĸ����ߦw��u������ݻ@�l?G�XFj۝��!���+	�`�E�?��UJ�Xה�GSD+�h�Q����'9�KGgLh��/�JxƷ�����U�VZ,�0���M���!΋I�'��qgf��i��\!�`���U�_AQ
�����[��2�ιH}�
�6|$qM�l����6M�����!~����&^�4��1��J$"���d�v�f�\�?�'�����=��uRbY��$]���F����	�#�����t�cc��Y�X۝!ؐ�oh��iC��M��N2t�iҡD?^�_�ޭ�-����C�UmR�Y���ю��Ɠ#:��/r"���T�%Pbi�����dW�Q�l�����
��������-ץu�E��ׇtW�X4E���A����%��6_���s#�-���$�×��:�`&�d �$� ��O��_�ՠ�k�
R:�*B�J�5)�(@md�����[cL,��6ޑ�^�����H�Q�i��[�Fv��JE��� �$11z��?b��_/���O���{�.MQE�m���,��zO��]b�.�U^&3�c�	���#\��#�Z��F)���0�f���'�r�mҲ�I��߫�Lt��bWL�������ю��ʅV�U�����^�D�7�'��d���@���%�A]�%Tu�A�F�G}�K,5��%Yx(|��G4�I��*s�'�ī�_�fe����o�"�6���0�9��婘�i�vm�K{�������^0/�vv�M�r��S
X���oVB����K`%��[��`��B�f� ���"T�	�3&���e9��}��[����3h'¥�]鲆�h�D�d�NN��fmY?%�D�^T�����|E�⑓6�Y᳂�$�	�9N�_;�w��ꑚ;\l��h½q�vV����*ܧQ� �>3J����Br�-�Kf���^AEKo��\�h)�u���a�$Kw~f����(��sڢ0vU���Ƀ ؚ}�E�K?(g�_W��/�-��)��T�'>����
��Y|BUx���{1�\;B�uA(KO�V��<XC�z:�ǌ>�Q'_Z�B�3�yF�������<-I0q�9��0zw��YwL���o� 8��1�S��bJ �X��	�th�c��Rp<j��__R�0�ъђ���Z!�ڷȋM4�[��[��8jya9\`�R2X�ps�`�AM�6JW�:�����Fk���-��kJL��x����R[Na �L'�w��>�쮑Rr�E:+�3ٽ��j�oKd�R��/������nԝ�X�����3��El�����T,��t�%��/��(B��|�%�y[���&a)@X��X��f�Ǫn�!��|X��ђ�A��wLcҥ�~})�!�o %&޾�����*Z��Ž�=����<�G����W�!��Nd>���!�yi�=(��H"9����t�)��O)�x�0,��ԁ�<xD{$U�u1Yyl\w��~y^]�e�����܇FZ�6/'4��@�e�|�j!���$j�8��w���T��f��w������7��v�ttn. $�&U��VF�P5x )��5��:�>��HP��<�a��,�����qM��������&�с��k;������3�rP�(zf,9#E�1��8���%���Ū����0�:���q�{vL��y^a�������x�B���q�y.��VǿX�`�r�4A�a�^{H6lH}j������I�S�Ĵ�x]엢�T�4�࣮E��"����x�t���g�hަ��ɇ��h�J�p��Q1*�DX�TV��s#5�Ī�t�u��R���?h�k(0��YhoZ����N'vQ�O��K׿j�-m������3E�uAᥜL{�Ћ �@@�j����9�{k�t�P�/p�v�D��$�����1|�;�]x(K�N��J�Q��"�/��/���XW�r~:?��[�������Fq�o��yxz^M�OzX�y���-z��~���!6���P��*�/�O�&�-�	`�d����h�/�X6����d�M���WDTƖ�>t<�&�w��h1���U����Z�Yg��f��B,���`� ���e�B�i�5M�Ƚ~��?��X�&��^�`�I҉Y\�X}��b����ʄ�"��k�����-�'["i	kZ(�� ��,q�8���z����6�k���-���{���M�U!���V"�cc��̢6�< �����c�%菹�UFw�DJ�=?���N5	��r��N�\8��=,��$Bd�Ɠ,m�'O��/RX�COCW�/ �C���Z�RB�*��ۍk6��m/r��AW�rr��8���
q�aL�Q�Ǥ�Ұ%��Bt���#� �Lhz��պh�+V�_ Bh�Ĥ�GSz�~��t-�[^m2b��7լ�A0�:p��%�Kz��h�0�I7����)0g��җ����xk����B��`�j����������~Odݙ���2��w��=�у�.�8B�=R�d�O��8�����žx,�=�������"ɀ�7��*���Z���u�ڵ������)�u�LQ�\�r��.qE�s@��O�ZH
W3{�p _��²2ȟ��"���rN{�t�		�rC���;\W��ɰ����p66�f�+�w�CR<�i�q��<�Y��A_r�o�2˨��.���į���9�q�AF�M联�D[H� �?�o�:�����D|&޷�	��cy�����H�����I�U9҄�)����4��4�����r`ˍz%�go��#�a��vڰT��'�l�*M��S $b��g�Nd��� |��yW��^J+��K����9i&�󎵒tx`��NXX�,ω�(�W�α~)��l�P�M�S�LqQf6on_ު�ƺ}�[�&y��C���U+s�$�K�?g&I.�����N���3�U	�3������2D�9
t��z��u��_�+�+"+@]bA��[���R������J����#j���^:����B]$�=�:�s�0��-=h[��R~�7v/���J�;Dˋ[�;˽C��Lzw%��>\�
���h�P���y�s�b)\T�����ma,���a�q
Dz�_m���W���CG�M�r�{o���`=�@Q�0Ө*y Ǻ$��.��l�c�p`�Ӏ0;�����e3�A�SR��o6�!^W�#��RE;��U<'�_�&P����p��!v֌u����I�=���N|L�D����e�i��4����j>�2|N��A�ɅW3bࡣ�8���kֽ�R7��'k�m���;��z�9	u@�}~z��^?�6˔3�ļF(�, �W(~�����G���{�m��F���	;<�.eo�=��̒V�G�L�������̸l��]�������<�;9�ë/���8�yA�`��Ϟ��;�}}��hxhi��:0JW?  ��&�%�l/y	gʹ�i��f��}���o6�3�c��Y�;5��I��l&���<��~�h��u���l4pŸ�V ��`�I�5�{�<"!D��q\7���}:y*�C�m|���p	�W��]̦�F���Wa\hWU.~����γ߮�pPQ�~�C_��$qI�^w�jHo(2'�E0�-N�*���8�|����w$�>��~��W�eDA���VXH���={�2u��f��ąiY�W�䠓cJ�L.j�d��"#��������( �����u�N��w?�.�&ZR���@@��@�c�9O&���T &"���p;��ox����;k�8�mV=��l:�
���^'JGž*qt�Rh��>ݵ�w栒WcW����}�VX�&��ٸz�m�}�ʵHm$����āx4�c_�iNd�R�Z��;��}��h�m<� �"��K�K�����]��"�0��V!��!�c��!�� ��_ЀbcN/�)�#�ng��\��q��/��1�E^"-�V���_q�T�2K�F�*���5M����^.8]nݢ�YڤG��i�Y7��i�}��f~;����]4���p"C,[cg��=��.�����`��v�ʪWӇ�a5��J�H�J��-QϺ��}�ē.���,�DȢb�g1�"@���0�&��c�.�"�������%�u�����l��[Z>�9�uBQb��;I"Z`�o��ZX>�a�q%�m2>����j]w Ӗs��A���#/<�
68��r�PB��Z6վ�,4gJ/�8�E����b6 �����5�2&�Ԗ�]�,|�`vi��F���u����_)�R�T֯Kw+�%f�n]T�:���Q��m���1�'�t�Q$�V�!0�K.h���-��@_������cO��{���T�55���=�{ku�o,��J2�9�v�#�9�J�Y����|P�U�	���'�B�S���bu�K�S���>2�I��ݸ�g.�J�q�+{�nV���������}Tľ @;���ߺ�0&��[!M�D�_�V�6c���/4���?MN>���f���6��TѺRG�B\
"�B�u���E�j\�8�$�wO+��;���<����@��[v��Ͽ!+!q�ŮD���V|s�7��ܥ �u�@�l��h�G��ǫ
.�4΃�g�"����w�q|Gع�z���j��b���B���ո�:�(�Ǐ["�)���By�V+��T��3A���I��;�3PJ�,��#�VV�������$�
��2n�T�Kd�m�$(������@+zb$Q����.��b�} ��՞���oh>χ3~�B�ec.|H�б�
Qmz���,�yLH�9��3�֘���$k�fM�%����o��h;��w���(�Zs��؇����̂���f��$��͎���:8IP;�K�?��C��#�f n�,�ת&W��O��'�ͼ����$��1\��=�'e�U�;O�9����Ak��м��.v5m��mў�3��l@�!�����4�)�фD��Tח�l�
|�J����N�{SY�����'�}"3�8��[8�b��?�%;��u����s\3��u������o�٭�P 0U�"�,���G<0aq2�{w$����!��d�Z̤�fW��h:��)5r�n5��X�Ӳ3Ƨ�:Y$h� Pͽ���W�kj0D�({2� �s�-.�P����ނ�|,�+�L�{�񟈉�8�c��Ƚ}�S~W���=�F�4���4_ۭ���,r7����_�3*���M��L��Ơl{8D�-O74-�
�j��
ӿ��iۛR��Sa�Ju�H�=7x��W��K-�B~��SZ�����T����r�{+��\ё�mv�X�QHE� �Oi���@�Ў�0����y`�  l���<�w��,q$�E8I��t,�����1�Wݳ�8YqN����Э�m��e�O��9g:�,�	�����I�l���5P�SO����wz�����?۷�n~�on5�_\�N�~/�\<��q��U w_i�@�����"V�h�>,�.��Z(��Fm_g���
Bx���X'���F��NŴQs�|�Nm�[$��7�uG/����wp9��f��L����	�u�n�}t�C��N*kyJJL���9"a�'��A��e��'�ȳ��jԠ��6j	�����>g[�{�7Z=><3���1�UҼυ�te�k`_7x���:.~ᔆ���)"yd� Y	۷A�Ͻ����/�3���6ʯ$���X�eOs<>�m��gn��^�	�*a��7��P��u�1��uZ�	ZҾʵ��,ɜ��i8��rN{�� 'f\������@�wܤ�`�8`z�M|3v�����Te4�!�h�1�]��Ŋ�B>��V�A2\r��̱��K\a��'m�����:��f��;#�%^Qj8ù���|�?P���j
ծ`��@�\M��D�
�)����CR�mK& �E��-�U�*�TJi�i�`�(�rt���|�tU��*����������bGXE�hv�3[D��z��YE��?,��ލ�h5�d;�T� ���I��s������%B�4Fg{�BçZ$��z߇��
v�0blË�7R��r,��"*sc}��ʮ�]E��\�ӳ�c�翥;H0�U���s񙙼���]
�Bj���:�}4���1�6�U�~�t'�
�8���ɓ�KͶF{��lt�؏��i��;����;�W�yD=�,i�}��5?QRʡ�(r��O���{\;VƝ�	
)�m�m���D�(�E��1[��B%PnU!�ͻAW2\�R�=v�7�=0������e~5}�;g�W��&���X����!X*=�̠NdT�"^L�ųr�ѤC��&ق�ffTX���6�KG�ë�q�ߛ���^���!"x��DD�o���6q&�V/��W��lcAGo�Q%媯 J�W��ܑqt^�y������%���t���.�G�{V]�Ed1O�ѳ3�z���@��d}�q�E3}F!uJ��+�jj��H����6����M�QZi<@�y���Az�t�?ԀL�ʈĊ}Fv�؂�Jٞ��$��a��X�E�Ī��/��Rv�D6�Z�b~U(1����i����JZEK�A�$V~o5sn�ǘ}"m�}l��i�9�&��7�5�\�x�\�g͎Đ�g�⛎3�;����1�<\��;n���Jr�?�d���Ck}�55�б�o��Mi�RV08�G�#�>l(�����3�/����)O+�W�.smB�:8�:�e����_$�����Z=_Q��3=碩\7�U�����8�^+��	�R'�6������pT���N��Ƹ�CN��`l1�"��.��C��ۆ"�_�_�<ғ,��e�Hy�P�w:-�"��'`�k��$��P,Fρz!��R`�j��x�P`!Տ�޳}D����RX ��'��>3�$~��j���|�k@��,|;��'3ܯ�A�yZr6=�V��Qr�Z��j>��(Yt�")~�9���#<˽�,v���`<����f�:���j����H��?�^�2H�SH,}p53r�>n���j\��)��Fa�'I`��Y�ᘹ\�It��2h$��FqT!x����Fc�� y���)v-����gV*x������ ;儏�tC�K���$0��O}51���Z�y����ڼ$�Uo?���Z��WK�/z��L��I�V���� h[�#� �����Ů6�@f��h�u��4|%��=�3�'z�rE�g�"��XBuR��!Et��M~S��$v�w��o���M��z�7&F��:ʕӄ
k&2�:��qx�t���d*=���D>QR��N}����k�GOT@W��q�{��6��KH��G�/�H�E�e�k����o�u��f;2��[O��m$J\At"�/T��H�ds���ɐF{$)��N/N#�z_ì�]X