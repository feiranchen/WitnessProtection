��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�w3O���d����>]5΍͚�S�K]�38v6�x��5V�Pe5O��>��{d&�õ̤S��%Xs�1RѰ��^���!�/�5��𨇈�BGw=�3f��u(��M�I���@v;��6�Ye !$�q7���ECB�� ��������PLg9<��+7�	�Fm�鵷�yPb�݅*5�R�U��ʸ�w&�F��E�s��{��� �^~�]c�~4����2��GĘ7����j�PP�$#�����xx��߷�D�0�b"I��[�e�>�x��<`ţ/�~�U�l$���gi:��F�̀���g >�r��ohrv���nZ����)ńFk@
3�T�e#?=�e���4�.)����V�l&����Fע#3?�o*ӯCIaV��*#��R��H�v�w�w�����6������yYۈShZ>� m�7�4���S��k��_h�,�;� rT��4'ݒ��[)�^��(�za� �qI�K��a�K=��`��M��/Pm�=`lc��$�o#R,HЉ�Z��Θ<�j!���?Ȭ���u����M����j�s'S��+�ҫ���ա".����Rb8�UU��C->��|Z�pͳ,�=N�@�8[���\�]�C㧣cN#��N��Z���1D��mi�s�{��OF��I�Fj��A�w��t�.9n��N���cϑ�*ď&�U>R��>�U5�U>��M���m�^G�-uaǟ�h[!�%�;��up��P#���U�	d��d��@�/-+�z+�$�RX�|<�M�&��?	�7g!�4*��:� (M���0��lc����`��`�kіqI�5%���4��5���9 ?[P ~��,\��$;��t���ڌ��?A��3-V1��{���f�y)V�pX���Q�чF���:���H%B��h�"֐��`�My�o@D�Q]�PK[K�$�kJ;�\���J�^�97Kޙ:�M-#��r�Rq�SҐ�̚����a�UO�һ=t�y,�@q��*[̞5�ƪ�,��JCŅ�¤��V�UQ����c2N���jʨ���xB��87�(�4��}	��d\���`���vF�76E`0�k��~Y��r�󆪤37��M��NV-U�X����"_\��M����?�O�6�3&*o��HM�iB`Z����"�,�z�-y��m"'�3�~���������ۨ8i�@�f�C�@Q�F/󬾉���ZS�L�F���@ZZ.n�^5�+B��Y��Of&����S�I-�ԍn��~����,�h�{��`�k\ }L�<��{�(r�#r@#Ƥ��2��hedJ��j�*��S� Jv��:�I/j������ <ɳZeă6���\'��7����ٻ�߽�xn�����%���_���!��S����S����*OqP��2�¼(��.A���(@頵�]����(�H`�M��Ay��c�֎�E���WB�H��3�S¸��Q��ج�5W�R�E#��Q7�eه�S����x[�`�j S�$���^��kC��5�A-r\�<֨�τ�� ���}7e�<;����X'D�;g]M�����T&���j���#a�x+w1�t#����bu�$�i�W[�7����Q��yҖ����z��F���v�k�9�9��Ft"B�{��UK,��{]��_��O�F?!��=f��@	�K�F�7Ŵ~$��.�j{R
J[a8��Jz7�� ����hI�J�A_���8)Xb[,G���v��5BY��Y�4d\k�$�x��~ 9LQS��x>^�~R��T`t{}�kDk�_��0f����pvV(�D�hk�����)0�Y�F�U�D�o����f�����#g�M��A����� AG�,\�i�><��1|]�����љ����[w�{M��1���W45��B�)�|�՛���\�����5Ϻ*Ɓʎ&��}e�L����I��0�L헧����x��w���8�Vťu3	�{q�AP��Yq�$ghZ�'XÚOzUI��5SA��o郎�_����[?��n�ؠ�e���6����+0�cA׌�� tj#���(������7���R�e�p5�%�n�[�#�=y�ӮKm�7�W����{Rj�=",�t� `/a��i�R��8A�E}($W�ނp�a.4sk�[S��!B}��SZjs�"�K�6����u�ы���lc�t���>����M�U��� &v���	@ީWv�feuԗ��JM���)A�w�-n2Ġ�}F�1�yg���ު���@��:ś\񋞪�*�X'�T�!�֏b"~e���߶ͥ�_��=���,����U5�r���^�uKр�H0r���`��TcӬ���y~\leI���)y)��Xq����:���O���\t��B�G�%�t��V͢��J!�'�B�ޝ��	+0�y}%_���z�D܁�$��f���!vB��8��<*�&���E���Ყ�lʬǩ�`���L4*�$��U�pbSf���U�l����ؕ�ո�h���a
-ec���c�{��#��`���ٿ$��C墛PQ p��d!���}��p���������Zt,ۧ��
��-�T��2Uϩ��4ح��[q#^��2�D������T�IZ��Fl!�%�I۽��<�;R@�d�˿��!��/���C�1�E�
�����%r�	7������'�6����	�y�g�(
�	s�Yҵ�G�t��n�3�ܲ�������H�-)ڻ�Y0�tOռ^�8���ȷG���&(�&���gj[Q�ψ���iC����k�fF�)&x���u0g��c�S��q���������X�>���sm���� Ji��"Ǧ�U������fw�@�f��9�/�IC	>I%*2�&^�:�j?y�H<;+��]Pma�n��U����a���<U��[s���T��8A��>�K�S���8�5�t'tn�҉S1�!SS\j�|������$�F���oa�_�hv�B�~QsU���Y�2P7�6�䄒���ZT�y����7]?�
��;��ˆ��0Cy倴e �DvR�ϳ�o�H|�}��pQ>  M@�"ONr�j���OK&����k�qʣ&L�d910,��
��W��P����멌���Q��o7҉�������Z� �=��'��`���q%T��U��5O�V~��;�+�R6)�IR�e�nk��>�n��{�^+��uA�@ɛo�� ��J $I� �!��U�K����GZ�	� ���q�_�I0��'������L��]w&W|䘪E?�r��~�Cm���D��J�6҉l��E������<	��%�_I��#H��!�	z��̆�����s�-�0}[�$�a-��T�>�oRqp��$[�@1\ߟ�A,2x��OT�\A�I�dU��G	z�ީTL�C8wAMJ�պJ���w�׬і�%�APԅ�kU� P�d���k˫�j��q��t�V9��"���YUߍ�*겴���Ɉ#r�n+�r"I���S}��Լ�1<_z^H�?��(ng��/��2_yv�.���g�m�J��WYUztՠ��s����H[Z70m���+����{%���Xv���u��A�(�VR�o����<���+���@����}w\��x��{����6뙄}sÃ��b	�1�K��g1Cd�5�>g[��Ի�p�g@]qaM4>�S�l 8��l��.�S$���r�z��d�F
�4K�0r'b��h�`��"�؍�u`*%��4lu��'9	5140�j�
�RVvp$S
K���)��<M��{�%���7��N����/	$�H��fEG�g-�2�T���r.VCX��#���-�9jo�NŠEdW��sG]"J�M/��*�'6��u�Ąl�
;/������X��=�Em�S� n�����g�+���(�$�/S���#?�J,�u5�H�(�j�_^>o�׀)����\_��Ef�p\�O&:
5?h�%��/�m���.��f���."x�u���: �QO���0��' ��)�IP���5��3Bڍ�ɾ{�?*V���P5����l8��d�Ow��)^��Re�V��?�I%⤐�	���&:^�O�M�/Oovl
��<ϵ�!�ԁxa�F�$��P��F�Y8T�،��~������\�^���S�mC��p���#:����\�&����R��S�HN�A�|@]�}D>@@3��G�	�H���'w�N����O��1�v���+ld��W�D���Ȕ�lyp/[gj�}\Z��/�������a:�pmn�A�SXZA��[ɠ�yo}PH�4���>��rz23*_��+>E�8«@S<�d����̜��=W�V��]��֡����rw�-E��*���Z�Y>)1�ml��4��I@��k�[%ha(�]D�������Nݔ���j���n�2�@�$s�?$<�
�E�J����ʰU�Y���h6BoO=M��<GT&kߑ���>ŅAr�N9����x�h�̫��E}��E�Rl��n֎�7;`���!Z�:fXk�r�p� 6Gb��bxC���n��g����r1
U�q>�8��{خ��G�UF �,ÏV׋��8�r;�FP�I�K'aڙ�|w�C���4�`V���`��� ���mp���  fx�-�N�Z�z7�����6@�+6�`�BO�y�q��$��������M�D+â�Q�.+@^�t��U��	��g��Qg��'�	-�qfI�{������!
Iu�*�r4y v;�%��&]�gD�2����~�z�?��`��$@d��?��+���p���cm�G���ͦ���os28�ݪB���UL�RN2�JGb��)���!�D�ڒv��}f�Q�f$����;$�M[��y �Y��y9�?��9Gx}��']o�9!6��G(X�I��lSA�|��6����тf4$Ř���`X{���F�WDI$Ƹ[ ����,Ѽ��ފ��14�{���L?��ؖ�z�嫊�U�<��ID�3��X�3x�h^�i�����<�O�s�j���?#1{-��.��N�[���%���w����)_�}z ӶyO�n���u�����4+<S�X��z�P`||��b��;�koȘ���������ZSl�#����B��kOܣ��HG.*��u�-gJM��� �0�Ϥ�K��?g�#��3z�վ��U���|Dx�1҇zT��i�:�2��~VM�h��\;���ܥ�q����*G��ߞ���u�Fl�jh�
W?��fFp�Uה'���<�N����w�F	�"�{��08���$3�M}�}'�ha����� ְ�9~Gb�0{��_�ݓ�U��G_c��n����X��Gmv�����=q�o���D�(-ۛgn���Xn�x2�@B�լ�{����	��hQ~�Y��� &��5�����挂�8���IM�&%�FZ?8B0�45�*$V�V6�ĲSy�� 8.��230�I	�����1��F����y�H�q#�� �F�2L�v���8��㲫�S�f_^!Պ��/\���k�j�A�����(�Q��o�7˦�f��"����\+�O!�i7(I�	!�C�����U����J��)� \��EḐ�v.�����d�w�Le$2ҥn��c,#�S�b�L.�E���p+Ynk�o�ɳh���ں�A�G��VS(Bf���Q8�n|?�������+�y��U��O�Që7��`�i��p`�;�HdI���f����Ƒ�K�ف��w��Jwl��A�fj�MaP�Y)�k�/�}nO����Kc�>�N
�|M3��j��[ʲQ��:,<~�x<��~]��+���q��ބ��%���1�$n���$9#<�-;�ɗ��[��h�����b��?= $/Ck�77����h/Jk)l~�'�B��ӣ��8�z��ݳ�F7�u�n5?�Od��V������F�/p�xr�q98��e��3����h�W�D�s�<Z�	1�T�L�v�-����S]�r타1�(�cH�\�Z���P�ŕ�
��8�m�����ji��$J��Pv�RKQV�jpak��,٣Ln
c���Sgɤfo�#�T/$�GBs�'�Rm)#�X$UB�͹�����x(�����uZ�K�$��:���u�]���V�ּry�3��)M��h�TPYbj+�� �����>ꙫ�H�!><���"|8և�O�7j�Mg��j2G�(����S����ȐM%/�^�KnQ���؊�4e��KK�8�����7z�RZ��]�~J���Az���xpc�eҼ&�!�pB�K)��H0f�ѪtH��i��?.\`5���̧�E_�� �;S��q�� X37��=�	��DwD�P�nҎ'�\����ұr2��Z7{��r��BT�J&�l�~�K�:�1i�ߛd����
���Ȣ�\�������"t� f"����)j�oGaw1�NC�����+F(�2�ۉVV�u�<�gÒ���YP�8�&k�^�J:~�$�-���ǣ��KǺD1���-�r�v�}A�k]��_L����*�+ѳ�u��tQW�������^4K�U�ʜ�I�"��T!g�G\�~��S�e�ދֵ`��p��U�3���� �~s.5φc��E���A7B�8�F���-�MZ�!�U*.�� ��B+G=�� S��Z��&�=�P�y�yk��_t~	P��c��J��^�������ҡ���i|��1�O�h3i@S��u���V����
%^E /���H�2+rp���zJ��'Ri���p�Ϲ
y*h���D�<���g�"|�GKgs㍳|ŧ;�O��s1wru�`G�$��z��l���n�H��Y?�5��U71��H�~q5š��ӗ����.������~�8M����mlz���m��+B��a���]�}v���WAd��5����`|dB^E�)S�Y�A	c���^��&)Pw�I��_��~
�!������l8�r��){�q�h��.���޴ Ű7�ӵJ�Ϧ�gw#�&�p���챿&Vd9�Ak�Z��{���?�T�s�P��ؐ~��E��)�rʊ�R�����b��$T���V�
^��$A|�A��4q��g�4�уb�G�2�߮1`J���[��XX�_��]��Y�a�S&#T5��Nϧdt��g����y5��������ۀ��%d9]In"����� P�9V����a�^���!23����\��ktU`;�EC�(ϽG����\�x,���&�!�I�I�M�o�A=h�1n���m���4N��۱�@��&�Oa����sj�t�s,0w�H����^m<M^�4M��@��?b����3��c����	�9����+��7�o�u��s���SFݍ�����S4�2��(9���1Ud�8�� T���NA$��I�]3�T��Ƒȷ�g��08��쁴/[׾c�Ì��Τ���R�- �:
Z�_/ ������c���,�޹��f*t�d@m�����w�6/�~��9�G#��߱%�����UU�a�P&r�|֔ /�w���=/��ȁ��W߬�i���©u����0�a��U	��!����7)�8x�(9������\VD��pY:��9�f�dr�$�BL0^�An��'59FU%Ѧ��xvf'�g!�8`��Om9�4���>����M��ӹ�H��VQC��I_��L���;����<r���I����
���h�/�ZD'����Xk�����h�Q� '`�������<O���㪶��8#�yr�8�14��A %��a�����]X��r1�(�-7�.�"0/���a��������'��8C撙
�w6n��'��NQC%��c�<��4)��\�>�I��
�c��8�,�J�֒�P ��EyJz:dsB�IY�����G���7`gB���l�+J3�`�q�Wڑ��"��aW�9��o���� �2G��iaϵ���eڝn�u�q��3�
j~��TF;(yDQ�b�0n;[�D"��)��D.-}�uנ.��̺u��8�-�N�}��t��s� ��ݓ�
���^g�t��c���k�$oN����'h���l&�/w�V�|@U�-�`����'��t6dk����<A`%�"�I\��Mce��t�:5'��<��H̯i�iC�^-,�*�#4"��$��.	F�9�:�f��m8=���Q{A�xG��s�+e�c�wB.�)�`�K�	.�m6�A��vh���㺇ÕZ�ͼ��?���H�0#�Yh~����i26P�X��1�f��+Z��K�B��I�>]�tT�~��j��ŀը��LN``cZ�e�skB���Q�.����:�p��#��m�6�d=�E��o�}0{�7�V�����m9��zM>En_��>e<��5wLG&�Y�h��ȳ~�!X�@vAp�r���a��}W�E�����쌹���S`	�
?0wc�L����`81T#a-�ۍ��=���8�-������9���NN���a5I�K���s,�Q���v������S��p26]h��Ҽ�v�����Ht��R��_2���ZH��⒬��?�.آi�H��M8�]>�Ѩ�ˉA޷,Ό4�?ǽ?F=h�"��������U�g1�Xd��Q�ʙ/�3�V��hU������O�ѳ�ҙ�ӳ���19�^��͟4(`֦���5�b�_�� #�/Ǫ�Uv(�ew�G��,*��A��!��È�����."/#��{x�nz��8�sZ�Y�Xg���6Bn��c�P���؁ځ�\�.OOpK�AQ�(�x	~^oS�ħG�a��0��M�����
CB�+�|�P���a�ŵ��ǽ�ECu4�[\q��N���r0��n��qn�@��Wvw�,��Bf�5+�+�"�}LW��k@��;����~�d�8���h�v�Y��n�j1���*�k�c�Zg6��
7&rF���|%��Af�EJ2鯀F��?#х�V6�D�q����\׻V
]��{Bg��O����Ϋ�֓'.��O��_j�����nU��'\��5��A�h���:��}��6x���_��}ۑ���� �������ձ�&O���#�h��ٍ{�iB9�0��CRͫF?��]�"۾��X$�ǁ��2e�Zf�8_dr'k�@(B,�`��1L�4����N���?���	�Jj�ц��pHzl}����"�VY7u��	�t�"�^C�� msA
3��
��=O��(�Ð�$0-�9:d���^�E_ch1�xk�����Q,(�;���I�k=�R��,M,[`^
�c�ѧB��&G7$ˣ�m�����y�0�&=j�y�4�*}���T�o���m� /�3�-��g�t]ZA�t�.M1�x�NGcK����"*������d-�n3��*#�g_��,���S�����I	�k�K��K�P�lWty��iJK�H"��8�����{��^'4ƨ	�z�dm��,4QY(%��^W	auI�դ�5n�#YWp��|�x}a1�
p�,��2�3/���T�i����b��Ø����M�A���#��Y�M�T�(+Xr�콌`����;�
�b�?t���Y�t!�JoJ�˰�+��lp	.9G�>�U�I�;^l_j�.�x4��� Vn�6�n12���`�ܹ)5�k�������}�<��vD��J�n��0���``d����3����m���W�I��4�Czλk�e�jCxγ#<S�W&~��3�A_��an�t��P>v2�t�"�����jH���FJ���1��ҷ�[w2��ϻs�'R։�L�^<>D4�W �p(�����M�#l_��a�B�K���G�6i�Ҫ]S7cJb^O�a�l̒�A�_q6�<��V��	N0g����I����*Y�����P� S.���).	cdNU�dp�1�MGiL����4�{�#�� ��j3g�p���"L�n���^w����*��Q3��U��	�_fA�s���I��TQP�P;����x }����U���A6����l�(M���W��(u��]�i�T�ƪꌀ�C�@t����T���bo��S`��6�u��C���u����V"��2��8-�^��|��q�������	�K�uF����W/v48-�}�z�T(3N�ข��}Z��K�M���6�י{6���F�Dt���q�y񽿲b�
nl�{/��p�^�?�{Uť�
���V��㕪�Z��p>7p2�@�����F,��ٓ�	|WH5��ū�浖����|f��2�Y���o�qv߷���ƌa�rw��3H/ހu�A���H��?��29U�8������nQ��+׏���gB�6�+r��u/�B��k�:ȂѬPE6߻)���a���К�۞1��A�:�)�闘B���QF��<]>U/�����X'�鵱�q	��v\]b�]8	V�A]�|Y�W`�45��ܥ�	���#}I�غ��H9��S��ߥG��Hj�X��9�@��8��1��@�6��(\EW7j��N�G�H?�p����@�)�u~|��o���_�r|�;��?����	R2�%)Ba�z���q���ˬB�Fޒ^>a�{pF'�����n'����$p���Z:v���:�Q��=�Ŧ/׷Ng�X��ݭ��N�����!��Pp�2eY7=G_p������ (���ٕ�qbF#�T
����T�� /�S)A{H�_D�9{�Q,<���p��!��5�`���Qs��M���d�"\�Ft�iR�N-g;�	m�m�e)E=��~b�j��®<?��'ȶ�n������45�F+H����ͷ8��#�G���W\���7��5nM��e&�����B�4m���������z�������D��q�/ll�a��;�-1�æ�������,C&�Wʫ͑�ܿn�z~<�
dM. (C	��Z�O���M�h�+��t���*���CIMbC��S�œ�oG��74��xU�hS5z�Z���O�<���f�|��]!!;)]����-f�{�����b�����mi�w.���'@��'�]U���y��S8;�_���o�ko�c31B;�-�H�"�|�s�J����>�$���q��s4 ��fx�I	�f4����rؤ�MEd�6����M���������o��c�2npBA�a�K��'NmL��o;\|�t(�R�_CI��9�t�9�'Ŀ�ګ��o/�j�f_S+	��/;��S���Њ�Ly�uʅ���D6 QR�������A*��˗��B���$��X��s�T�L�坃g�cŗ#�y�q�8��At���A��h�Wꈈ��e�7�O�C�����<���x���˟&U���=�#�4�t(���{2���
��9�H������0��:�C�Ƥ$���=r[z�٧Ju�|?�k[D������d��I��
jML#��P�8��9����r�0��/s-��X]��:��Z"
�2p�o/��,}�д|VI����?������+���G��3c�+����Y4�#���7e�X�77�X|L0�Ġ�8�R/rE�B���� ���u*jp:&D�g�oJ�4j<�1����wg��U�{U�(���Շ$�D�<:(!�"��)��p��M����1�Y+�C7Ռ[�wIr��"�:*/�L=�C�����n mj���F*�)�j��Ŝ�k�䞆+e*)�jiw#Uz��_�V!���M����Ns��"�&ƻ�n�#/�Ё�lZv#�4��P�U�+��H�����|�����y=O|d��q�(����l�K��6Co���O�E?構?����T���v	<f#�jvuRL�8��/х��˻�촵MJ�9�B���Л������RR^�Z }�Ư}��j�Šl	���u�4�M%>I!�9��hT�Rw�,�ȓ�&ڎ�v+n!pǔ �|����/5�&��l�Cj3˼���~B�͗������_��e� E"�OѮ)�`�_���7y�3!�,;6�0܊8�B2���5�kȂ�Z�r���z1|��n�'/�P�r����'��j�п����/�%����Hc~��6U^�ڇD=|c8S�x{hT�L "餼���*�F2"[��ٜ���'�Iә��(3|��e{�|����`��(�yc7�k[>j�j�^�ċ�ְFU���];e"�c�#jYnj�]���//��D���j���>HI�.rf@��i�|P��ݪ�NT�T�D�$iʍ�������sM��Kj���0�R8cl��V�px�����N����E�!>>}n��?��Zx��?Pq��������O7@������
��B�Z�!3)��՛���E�X�n�u��!D�s����y;�=���~���`h+���ㅍ!�4)���Ү8t�T�m��
�u�}S �d͜��ڑ9���g�D���vκ��D����2r����7خ9�Ş�H���$��֢�GQiz�S�U�W�c�V���b�L�VU��KzIW/��]��(vu���e>z�tZ4:���3t�G>{d�$���5.h�Fݥ����Fcq���=(�߸W�)n�X^���沕]i`3L<f�B^3�*����V���U�1)�6;�e�a���)�W�{��vb��ʢku��l�#9y/�u��*{�  ^k�9R��h3�%'�������z���HGjo�2�
�����>aE�А�EbчC���{��y�b��9]`(�O����d0vSʘ�!f�'���NeڊC
N��'�h\c�_���a��g�=��~����J�~�� ��ھ^�˚C�Ϛ�5�V�������3��Ae��Fr���c~��2��W�k���8��B����u?�(6�����S�maI�e"Ǹ+'�Ҋ��	s�]���D�%���c�n��0LT�,f�)������*��Ha:�����>5��rt@K���18�es�>�	T N�B�A`��/���t�Kd	��L�0��;�ag��<��F��
��Y+�ƍ��%é[��ݛ.ȼ�2��8�,&+$�&0��������r�Sr����%�D%�V��z�[��OkD�h�s����n���VE�}����B�z"�E�J<!vϿ{��%��b	xz�8��E��4�z:�$�7Q�д�S|4;����|�c{�%��J�缒�R�%"�.��N�cN���zv���B�l��^�W:�c�sq�Ј>F�.���:��`��}��,I�S�E�`��e���I���QIl̎��ӥ*�߽Zl����>�g��}�T� ��
��&�yL��eK�U�8��5����sAOt�I����^�e?����>m�n[����7���R�Ш�\����]Bi�7o����T2�w�&A�a8�����i!ˌ��$�3=�Rx�9Y:�"w_�V.�f�0HYdK��rMi���dC�
��LX�rb�z#����J�4w7V%����^��Q3v]� $����CUM@���8���,ѩl�s%�c����G�o�C�M%�H��j}L��D�Ҙ���$	1��Q� ��r��H��B����x=+<�\��)���@YȤ-��� ҷb-���?L�.�lB� oF��?����@/��,��zb��xTCQ'.8�g�uơ2:/%EJ�^���*f��xC�s8��j`���d�Zpb��Q�5T@=��w��J��Co���i�e���sڰ �uz�XrY�ٮ���������pm{��{3g���A9��i��>Ò�r<=�29�O|Z��(R�$9�3�㿵����f�e��2T����eb���"��e�Ӕ�@^X��Vl��UZi���Of�owm>�5�$���q�V�9I�N�oY (b$nx�'C`v�*_�&-�#�+�:�� \+��3��sf�^7m�A������^V�q�j�+f���j���$ �ɾ=C)�@[91���{M�����,~!��B�$nA�O* 2,��vq��-M9�u�GP��,e�ƾ���`?�Z.9�,�Ց��ēf�æ.|��_.��A�Y@�pk��sk�q��}���}�٬��]�WGz�u�aR��s)�& �c��l�
s��U��lFF��	a���;PT%��s����5Xj���)�l��ٽ����R���_ת���0d�G�4k��"���"yM����(�
w�*A�X
��3��Н����{X��iqm_陏+��]��xbI0!I�]jF��}�:�/�`����ǳ��a�3SI�R�gAc,�mgp9����	�ҏƞ")I�Ѥ�z���!mE:�+�RJ����s��ɞ#�Af�8��ӷ���7J��B�NL��[�7
P(A]�Bq<<f�]>��HY�qq��O�e��PD�~�*�n�OxǠ=a��	�y
�_����Ȱ��B_��*����tG���%0���<�������|��-������s���S���c�wA���U����"���еК��f]Pp��K9��iC]k��?�q������Lт����WF����8=�!����@#�p}�2Z�}Pp�	�\�o����{�m��jڲ�[���?��vnY�����n� _�i9Ok9-VI��v�&���nS�\e�v��0�&�Y�V-(h�����ӎ�$�Ox7�jE𩲇E�Q��Ȁ�x��~�z��;��7b����{3\R��L���/�pu)�B�Z��`}��������}YNH�Si���p�XS��}�����m_���Ei�b%��f�ˑ�=#D�8�|~���Z9�簾!�����P6���Rl�g8Y�Θ��ꧧ�g�O0���s��_	T��sD���/�b,�����J�!�~[�<wm�R�IP�t�O�Uȥ��<P��x��?���T��A+�>� '��B�]�'ƺg����R�U��H*��)�nV(�s�9��1������Gd��_L"�-�^
bu4��D^�7؎��9�4�a�t�Xi���~Y�}�wu@hv:&9k����b�,�RҮ��^��>�z^�/*c
&bZ�-��*R��*��σږ�+���"4L��j�g(9'��D�ί֨Qm��$/����4���ŧ�=�Sd�;���a�<�
}�Z�Y����/�+��ѐ!އqu$�rV0�l\{��PV"������l��67Hh(dVi�A8q�QϾ�� l�;|b��HM�`��{͂�#,�<3���X�y��S�.��ٿD��ѓ�cYO1�ݐ6�A;�j;��Qb�N]���8U�\����j�mC�$��vɃ����%�0f'��o-.ރD��c���j���e��/B,�W��H���+�߭�W�SI�O��ق�k)�"mV�c��D��������q:|i�=OX�<n�?��,����ĠyJ��^��1ޚmݿBx7_V+��?7�Y	U�i7t��h��2Lkq�2S��A,z�sN����X^�(�5�n���)��`�9`�J�"$�ߦ�:�CWe~i�T$H��ґ��Mלqo	+��T�%w;�d�l�K�ϓJEx'��I�}��r9_�e�{��c����}zf��p�7�]BΑJ���nl")��%G�-�	�I����f������N�p��X����V��)*A���������Q��M�ʖЦ
��m�r��[(i��;Q*E�@�~|��ǰ������*�3��d������-X��:�U45�^F-�6�1�#o��W�K�+$�‧s1+���W�w�P�~��:���?KqS�Tc�����^�tj �h���X���¨����=�Χ&X�K���w��2�����6;xܬ����4;�@�U����^ ���.ͧPb�1��=:�hC�W�5��_v��n��e�~uqȫT���ڒ6����Կ@���2g��W�,�\L�����Ĥ��4�'w�JS�؆)��e[�ۙfv��x�(�aݔ�>��&���1=r�s��k�I��m�;Ʌ�π���;�n�x����������6ףgd�86�n>���Y��]�}�,������v�"��~%!Iz@
:o��lm�8�u�\�i�W��O=3�'�F�;A��k3/���],�?����&�W0��:�qg�:K�V�$4(m�a�F<��m�j1ڛ���+��������f2���zP�2K5�p��H`�<�� )*��z���R���M(�?X��e������=~O����/z�����U�(�H}Q�5��[���g��gX��Wأ��AW��ܪ�}���a�̽�(O��:k'������~����B\G��_�]C��^��0�=��h(��� p�섵g,'�Ya>m��M Fm����>0���-�a�&��yHg����OB/@���K��`���{�=Z��ו�mv�X�x^�j��z_��v�d7)�е]d�GZ݆%1�'�M��2�_z�����0�1{�0��o�)��~���rUA��Z�,!�odz��%B�d��.�����hA~�_c;��"4@L~+W;�L�$w����ݠ��1[|R̞8��>��ԇ���X0O�ݾ�k�~V�Xt�Sk}�R��<�����їQM5�m�X�)�@e文w�p�����gc&�2��飅�;�t�=Nw���`F�4$kDu��H��(�������Ke����ؽj�8���da뤻���M�-Ym��z2�4���TE�1��A\���)O�Κ��ր[F�u�<�w���>��>@;O�"�3w$Y�}�.�g��ܷ���\4a�yZ��@j�)�k�/����|�w=�D"�����o��2*')� F�:��W�1%�p��!r�y3�
�)g�Kϳѳ\C�5�m��r|�-�"a]�fy<��Y�;�*���{fi @g���'��jd[���<#�4}50ObO�2WV��{��ra+E��$���9qm�s��BAbd�#��4���cAe��q��;�2�w��)�&\|Ӯ��UT��	j�E�<e�dX#ݽ1N�vPߦ֙��[��e��3�o��{Tr��Ϗ�&��|ۃ�l?\ΎN�+?����A���C����1�^C3���+d��Wl��W�ث�Q|r��䪂
ѣ�p�1��Z�K�єdcaLEd<-�62'�K��^�TBԀ�ɪu&e0Q�T���.%���]R�A�{�^D����׫���G�XK3j��:�,�ݾ�AXbA�y�	th5��MQ],��8�ͭio?^=[<jy�:s���c�u䙒�����ʖg�x�Ş�Oj��+_d�s�a}��d�N�'%��a���qO�6 �� �#7�6bڪ*e��
���%O�jY/��,�'Xc2�K�w.��X1�1��{��!�X��NEsv'��dh��u��}��z�HD�A��Vyg��(�V�6�屺��W�bW���Z�-��9����˃�W��V?kR�A�,b@�KX�� }W�� ��Ս���\WJ������)t��v�*�P���>*ѳ��ۢ�����sA��T�ԛ�3�$�F%�ݍ���ޜ�{f����;A��Gm�Eb��X�U��ρ�GKU'�ٰSS��ئt�אp��V�}��-<��<�����q��pY�{�o����	���˔�����v��⛲���z9��G��J�@BwD���GĚv�_�=�M�+\Ҟ�Η/nk@�yz��c���\�(H���U�E�#��u��Q9EĀ(��4�Js8�N�Y�q�6� �e\��t�{��+e��9�{t��������Ӣ�Ǖ_�f��t��� z��qQ7-_�o�^=	h?���d��R�K��U��@q9nT��h�<�����>��$�1���(�-��1�/������l��gs�Q��B�Y_�ִ:�δ! s�{V7?{�n��x̅�G�A�|�£H�-_d�MJ?~�"P��l7�b��d���0�3�><��q��#}Hw��a=�#�F� a|�Uv֑��U��DfR�ۂ+����M(D���}��5������i�\�օ˥=N��~Y}���c�.�>/>8�`�p����Jㅪ?*��7{*�˒��%iҤJ�i�טk\h=�ҧ4��f�֡��(;�Ev\ �`l����CLN:t�Q�L�5Q@��O�0��r$�}Q��s#��hY�<krj���{̂��E;�]��BΚ�袕�,�[0b��M��RA������O�%��G^`Ӳ�z�*奌X�L!3��0�N�W��fJ�l ���;hZ]�ʵ�*��&�\���m�K�y�
֙�Z�Ȗ��*dG�RdY'q��d�ż��<�p�'t�} ��˓��S��������S���/�p��ϻ��2�~:B���5ڹȯ�q�YiQ��6���V��}rT�nV��(�\ ��
L��,�܋:�U�az)w�2��5ˤ�&�,>��~e���n,�r�-�����6RH��4�h�ݖlzpw�>,�@F(m2b�D�'�$�h�bc�M���I#!nI��F��#B���ĶfҢ;��F����Y5�T���~On�,�&�2L�� �p��F���?�4;t��q8#8T[�sE�H(�$"l�DYH6�G-wh8�&[��B�a�4Ì_| *�.'����(/�6p�f]V�y�6;�� }�OW��&=�$c°+��ҩ���H��pn��[�V�V�UY���B;����*�-�&. ��O+���jN��
��'���-��''#/\I��Xg#[�3Z�/�1%��5;���~��Z׫�U��{t�(O}x�2�,�hE��,+K �0�QW�R"���=wcA��U	)Mt�z??]FN1f�a�%P��h;�`��7�8)�ੇK��oUY���O:6r�l�m�$�ݐf�z��ߩ@��F��6���K��s��k�uE�iF�/PV|�h<��͂O@�nV�Q*Ύ(W����������_��}��{H�i�ʸ�]���T18� ���#���e9k���	.���+�/�q��7��!�@ .C�����x,���g�Fzl���F� \���"�7N,��7@L����׺7�-k�`O� گ.d�R�|2y۪@
7dI�Y@�&e�ߕ�g�1��25�{���:�q��a���l|�׼��1#�z�#V���iE��*��FQʐ��_d�{[9�P�����b��4>��O�u_��@�v@D!�����i���v@=iB�����G�p�3S��eш�w��$�U�=�^�_��� ��h��xH��#`�8�3ֹJ��k���%J��Q����̋ �+��ws�@�Ik[j����C�@
��L�����գ��x�V�Wݟ�)���:`���b��_=F����M; ��\ 	� ��!����z�]B=C�������&`p#w�5;u���C����Ij�&�����:��k�Z���0�O��������SQ���˫isA@�V�s����░ul�k2���3Ca�E�Ʃ��ԭҡ�a�ކ�Y��t��>gI�QFhN���mӉpT���f�sR��{!�}GCb�km�D}�̾G�r��0��HȖک`��Ԁ0+�|
�^�����f��fm�IFH0���S�B$GGlF��w.�
m6���p���m��C�j6m�Lhy	���[x�=F�ul��<���W�pGx!�֚�o���wj`ȫ#��2u?-&����ث�k*Is�����"�v�'նO��̄���c���u��R�������Ӭ(¹��җ��NXo���(�Wv������[�5�7�4�I�|�S�<eO���}�)#��r��W��}�'�Q&-�t-=�e���bҭ*��x�$&#�0!�W'Tm鋊����$��#�g��u��#�B����M�"O�&}�QG$�Q��n8�L?�&�u<7(�=iXţ=��n����ϭC)զO[�haY��GtT�������kL�O�=WQ�[�Q%�y���#�0�w�ʽ+%5l-�Z*�#]cA�$+Q�e�wI����EaBL~;���ޭ����R��*����ݢ���'J�2�]�+;sm�<����O�[��p�����J)!�d�^���R���}/$4rd/Z�W}�"{_�c"�˖[�"��	\���Uu_9�	�x�ja��"m�T�D2�� rn�����֓%�[�6Ɨ԰]�5��)Ȱ�׋�S�ܫa�$u/ �ߜ�Jb_va\9��&r�m�Y�O/�����T3������T\������wu��h���$�9�8��K�n��j��q��4<���$U��k�u���/	�.��������=U��{�+�#��4�&g|��HZ�:^zQ�(�;D|�?�-�j��u��u6�6��}�yC����8�'ې7)��֐�	���	IUb����0�Ӿ���L՛T�y���g�^<N�0e����%�kI��(7RtT	`D�\06p����c�;< P.�N[>M��ك�+���>66�Ǥ�M�D�������K�?Y��/ļ��C�re�� �Q tF�-ƀpesQ7����&��?P-�3Ѧ6�<���94���*����=5>�w���8Ft�/=%4FyRѼ��$��Y[����O�`q���@��w� C�F��'��=�Jf��{|���Ğs�����r~�A��H��#�[�q���Td��{H�^�5,�7�l�| JXu�/�Ȓ�1~.�E�������R��$$Ok�U[���S�KʅlƟ����g\�;�&9rO	��v"$��j�g���v䫑�������8��^��Z霝5�o�� ���KҎbh������{k���T�$`��z�@]���5��Ѡ`R�z��t��B�o/�
�}�9��d�F�.G�^����Y��Y���r�~m�J���2*.\0�G�p�	j�T�cb�ŭ��L��w*_�P8�]G+;��M^[�`=M!�J��haR�D��9���!U B-�i�`�m+_y� ��3^����eC�q��,ٲ����	1kY/���25�#M�~W��� -2��kz"���e.�(%&B�"��A�L�=�Q��U�(0�E��Z�Mv�H�kߏwtP�����jI��₮�*܊�j܄gD�:�g!.A��pAW�:r�����M�N�=����CS�2��g7z�༕�0�%��J�[�H�G.I=�wv���ȥ��Ǥ��Q�N�Xip���w�xϊ��bE��ր����΁��vBT�0�cTE��p���J��@Aq�
����~�k9x������>���fk���]I�U+�.�T?��0�Pٚf
�;"{�v� �{Te �a<�?���X�����cm���l�����Ǚd2��\��R7z/A]��ul@/���z_���+@2zx���~��z�&�ʍ�C����IR.u��ۊȷ�7Gw��LI�%F���WI=S��G�RUt��W>�܅W�q�D*�[^:�8��0Љ��7��V����HT5�X�p�þ��L�&>T��>���b>���Nq'�! |L���y*f�f����Q�`:��g��'P���8��g�4D���X��C*��E���O"gV4������*��E���s�ضT���������v��o7ưH����k�8}m#�9��ZRս����$F�a+A��«2���)���P)�ʢA_4`|��v�^��W=7,�e�oD>ȥ~��6�D�Q�~FRT�+�t�.������t�4�$'�^b�-��|�|?������%��X 5
+��
 ��tSx�&�[}�q�^~�6yb���0^K�`�@��{���y~�}��u��X�6����q�_Y��u����ȥ�Ȗ��6X~�� Im�nk����W�ϖ���J �DV��pT�5Ǵ�]�!���"�)>He�O����ᢓ��7Y;'#��~�V ��t��jH|W���|����M��:D����癩]�Q��y�{`Oj��6gL^���u���q�
�fo���92���À2Z"�^p��)	<+p~�
����{�q���_��F���Mj�u�W�����}ň�%�l�m�VU��0��m֗x⽭�<��	����&���:Į6��A��K�#Ӑ�3��6�ȥ�ہ ڻ7���im��Vn�=N�O�g�uh���lx_0������~'�X�P���T�������E�u��<o�����nߗ'.��nz��3*��qO.�vi�6T�40�=4kӓJ���O.�a-=��������@ʞ�W��J������n�=� ��Y�in�r
d���>u����d�~׈�E��x�
�oH�t�rj�h��|�v�sBsF]���
9�,����F� J�׮����L�[r	:Չ�n4�������$�^>,��T&�+���ktaH!�ئ9�3�+�S�O�Ox���y�@C�	�Z�U���/P����p���|�j!�CJ���x:�JJ�d똠���u�F�t]B����$4l�"ǻl��V��',%�[�n�0��M�lZ��C��kn�Ṗ�Yj\�韪e���Ȣ�Q[[�B��=Ex�dF��ظ�g�b�-j�R��L�~�ZY0C�}�T�6�t{��v���	���j7D�8�Ke����q�Q
A��S�g5�gI0�������I�5e���o��+��K8�G���t���U hd���i��ٴ���#�r��%�Ȏ{f$��D��jhI������n���%oɠ]�F��hg��%0���w|���B[�B�X��\�#�GE����	2�^[3[���uE������(�u��`���$[ |��{��w&7w�!}�c����c�>��ozX5�c
�� �jQ߃G��J5��C̟e�u�~�v�Bx{_��i@�N��Ն��d�h��$��3I��Սa����X��Ƀ�(]7�cM�Nz���i�<��L�-Ps���4��NxeE����;h��kf����+.4���|Q�x\U���+��-|�k�H_���|�A�=�ǘ�H�悲�
�Ր�9R��(5��V:�DG���z���>�%sr��I���a�����ฟ	  �G.%|���A�}�YĐ�W�����n�v*���p�M����j��ŞI' 3����`�!����U������#I$2�hR�F�C
�	�����~y0f�a�0﮳���#�r7���۰!o�0(��dP�A$4��{/�u�0~|�B���aE�E���D�!�6[շr���f ��K�l��.6�qc�������s����g�r_����.����Ր���ʷi����Tf����
��֛%���3�,.�.����%h��HW��;�.��֨F���7��ҳh�l[.���F4�hjϤ��@�5��ͼ�5���dS?HRn()��N� �j��/i���EGodY҅��q�+3�NJѼ0"or�q���,b}���?:��n�n%�xG�"��T��wd,<`'�{2L��sf/X�E>����mن�y�x1�-k60e���rBs�L2���\A�/{���I��BEFa�jw�<2vP/�ëXCj|���(��ޑ�ϯ��ۗS�����>j�Z��W7";��������/�{u���%�'`�3�6֮��&����Lz���#�����躭~��=9ȸ��r��_�s]}0����?"! X���L2X��(�<ͻe�{,a\�S'��#�Ly\�|v�ǰ=��\����2�=�� `���p����-gu�yf��ϡ鵂������H���f1ܱa$�d0�Zw3�QD�=@v�:�Ť�~��$�
�m|r=e+q�[�Um�[� G�>^�w�f@�!;�����>'<[�c�+V�q���VX�]>m�$~m\�X*G׉?��V����/����L0hq�S7���p��L�J)���j7���ߴ�H�Z��I���MaX^"�%�c4qn~]�%���8Ɋ$r��ŉ��e�5s�.~�R�z�����p�+�0�z�]]���DS._D)���Ig�!��0�%us�q�ү ٙiH�'��/,`:ny�㽌�m�wy�W�m�KbRF�������O����|�/�v�Ωsgۼ��%�
7�p�9|�I�l{3��f�`ύ���=-b�vE6-�P�*�a��=&=\����+�ۀ��m�n��H<�ro�Q�@fv2N�Փ��$(M�Z�|.7o)��Q��a(]�Е+p�c	�f���J�3�q���_�i5����}�T��:4!ud�j;+S4��`+��]�����ZB;E�iY-!̂]��#���Dpe-�Rh��Ǐ`��o4���{#X�o�l��FI�s�$/S����Ec�	4(O�5�Q[�G [v�s9���+W§"����?���'�=~"��Ϗ-A3��TiE�mof>]���>%?l<ZVX�F%�Ԯ��ȥ�X5j� �f��ו��Q�b29��S|�M����=Y���Ff��-�8�b��#=����̘�\#s�7Ω�j̱�n��k����鑺�{v �[ʞي�c�uBy�rG��l��eNLl]�ŰK��K��~���X�Lt���*"��kEq��c�V�ц��@�)f��\1��M�8S�c6
@��H��
@hT/:4u70�B[��2Z4�db*��0�F��V�­��T�c�F�[��?��˧'���v�!&�q_(�G��p�ǿ����?S��U"'�?��aI*`��NV��U����[w��x������J�<��ݣ��Xрr�0����;��F�9͎����/]gU��^�d����{������'ܾ�e�]�K�f<n&���m�H�S���q������؏s�K�f掽�L_q�ṏ[F,�z�o�����K���W��~<#���B��������FIʊ�%E� ���(�R�,1dC���D�bS�_�m��Н34_���J�#���~ �9tU�E=X�q�xŁo�*��^l�uf�<��r���l�RI$j�i瘧����0� C�>Tb�+~���>9� �H�aX I��`��⌉��/�@�S]��H�(�agf��1./��B�]�A�:'��1�bq�`=xSO9Cf|�OМ���2���?9��40tB��4��/�a��.Z6�5zTP�8�y�VH
.M�ɯ0�֥��Z��VQ��m�8�,�C�����eM��d�2�6��B?�q�%D�����e*�EA���ݕH�����clz�M����ʦ�_ѧy��s3�W��s�¿9!M�&6&� 2��ķ��ni�o��|�p��C�����Q����9����&VZx]T�k$/K����U5�8�Z�*z��3	����j����Zgd �o��J���)��vB��'��O+�����P�iPH�4�h�v�T��Z��w�I�@,�Uɪ��fe�X�%	95���M�@0Q�X+�Ԃ�ߤ".�,W_~$���|n� S��OF�E�1_37y���j���3H�X/�\jU\�~�hγ����=	�f��uA\\ӓ��1�v;��wūq���P�j@m��-�܅HZ�eP��3��0�QoOGæ�f�����6�WG�p��(�*�+ ��/~���a�j�<YE���^��K�m/2�	��:���9׃tl�(2v��y�������pq&0Aϸ{y՛���E���N��)i��3��Zg�~D-��� �!ֿ�xZ���6�4�
af`1��|��;��5mV�X�g���T����Cq��V��ʿBB��ʏ`\�㬙���U�o�z���ɞ|| �.<���ľM��㧼�ʄ�g�7pMjj��M� o�E_
|�2��m#��v���w��w��q��+.N�;�Na�AN͔ɴx;�9���u!v[��Mk&t�'�Z��m�,�ʁy@�wJ��O��3�g������̓Y�a&}kz�,?��Q�s	��Y���o�߯�9ǫ_��"�4ظ�#!�t�w�I2i+Q���櫋~����;�����k��s�x/��Z=�P�N�
1` ]pK��a�O޳��⿙IM$�r��$�?�چ!@0��	����֍C��>���.B��7�_+�����1e:O3�Nx�<�F�WC����r�w�����r�V�j�f�����,�&Kh�NF�bJ��^S)�#ŦX��o�%*sD
�� C�q%Q��|��G3�M���r�R��j�%��2�UB�����)��/u�`6��]_�^�ߣ<��!��"<垆�v|�y��������&|�C��<�A��X�ː����Fh�"�U��f�ֽOk�^��w�?|�.G���i��}���]��5.af�.Jb��0�g��)K�0AFũo\@�LN�R���C�.�Z���6�������@'��/Ѹm���no3=Rl����uM�ͳ�� �Qrc��� "���[#՘)����؋���ML�2~e�+��1��qFJ��>�[�Gq��иG.a�".�|��`���ϥ�T紭�����?rGx�\=Y:�΁��{ �yS��b��W�UIRhQetcwnҭ?���YA�zl���o�^,qV�����mq��� ���@�������S/���k��)��kr��Y{԰#�Ò<jfg��4���t�Tל}r8�����������*��Vg����^�m]�~����9�N�%t;��uZiH�$�I�	�-O�էmi���� ��(����1�Ɣ$g!�rj&|>���_A�� �(b�� [^[�4"CB�]�B�G�#��s�ln����Q'\ؚF���{u�Yd���������h�{O���U���>M�ފ+���y.��1��}���Pz��$?�C\@wP�O���޶ �!Gz�|�ZQ1�O�ܣ�:lA���}���f�ԊZf�*N����������Mu�Wޚ\0��P� G83�&�m��x_�n1��g�D����J\�Sc7���֛)(2��u�R��J��}_�Rg�hx�A�ͤp��2f�����O�ܜ��F�'�q��P-,9.��H��Y-]e���H� y���Ԩ����Z ��8���M�r���jfN��&W��W
J��#���K]F6N��$Ǹ�� ɐ��N��y'�9ט��U�6;hmج�x�(4����3�K�k��D�y��`�ڢB��O�K�SP5(�wv��˽Y�Y;�10��Y�����
>��l���l���,��K-S�ým� J�YY*���f��h�i5~7j#�d�J��Ѝq0?�06��������t5F��y"�C���~�cW���y�ӗύ˚w��@��:��A�W��aW@�2�&'���wg���[���
���]�&��yؾ��gL��	2�Y��5��شn���$74���#���^[ ޯN��A���G����}(V:מ:1d�u��/%b[���S����Ɠ2+���*y�G��/��;-�mW���"(MR�j|����9Vk�x��I3����ϸi�ґhZnd-�T�����f�˵t�7���H�~���W�b섂��z6μm"�^�������"�.$�e�E!np@gm^͑��x�m�&v�9�F�֮e��9�6�v����K�o�(�I�l�z@#������ݙ w>Q��]^V�D^�\m�\w3J�s�R��R�j�fN�Rn��g�R%�(��7���[ݥpJ��!� �N� H�o�9�Q�Ή�����ҩ#@Ю/��	�l�/w_�� ��Y�p}(�u�?/�q�5���|� x��ͤc���Th��Y_k`Fj<���Y��o��õ�:�;�Uj�aJ�A��Ƽ�<U����)*��{ݧ���L].�cD7ui������\0�+I96�s+�����M`��g���^�����6=Q<��ICwf�,�.O��	�h��d��B%*o�k��ٚ.�>����ju���h��YJ@��{13~o����'+vW�l��эC�rЇ���Lݬl�!!�?���y�J�xk����C�O>!�Gi��Y��d��G���&2�H��k�����w�3���hT:e�nA��#�;k�?�-;-���&���D�r�G�o"�s�ߒ9ǥr-`�t�AE۟�~��M�m��ύ=$�
O�r�V�BC����;uV+�o�8C�i'$ҕ«���L4N����yz�$���&*F����� �Qe�!:Ʈf�Z���ح�����N���M ��;hɈz��}?]]O��=i|:t!	��^Cmom��<D"X��G��y��?���b��.t5%���l$�7v�0.4u���c'S���U�2Z^;�'e�hH�WL���A��.����Êt��?���FU�5�~W�C�!�е��3	��LL�A8؟��Bq�Q�z�-���"w��L�g�j��ϟ�2��{�:/�#>B�	�@ *86�:J���6�����i�����7���ꔸ��i�U
�sU��i��0��ܡrc��(HL�+����cZ倕h��
�n��%A3p�ʃ����B���J4��ζ2�81���q��)�f�o#Y�Yӡ�`�H0v����O��4jc� �\b�zв�O�*��;�1���R����23�9n��aF�ڱU��Uߝ�~ݜ	��הy&��4y��gNȠ]��w�yP4˖�$���9͏��B���
��.T����Da���}��$fe��nHڗ�\}��¹H����ؾO� e��$�j�k���᪞hK���I����$�b�*��S�U	�
��Z�c�u�����Ѻ�;�.��Y�wLPe6�{ݳ��(��Q٥f�����J�hŋ�����|�'p��>	t�4U�y2���~b�9u�w38`&�m�1Zq5"�����N�Ԟ�5�F�����aK�v��������v	��~h�@��07�j��#�b��a��?�a��.'J�y+����~J�.��
��Dx���8�vV��~s����7�)�C�c����G�DS�����@7�U�#�"����؈*T}�]T�xUc���t
�R�v6�=~Ҵx�zy[�v4�d?$/�$��q�B�I-O��cY���H�/�JE%�N���� -N�(���ɲ�y�L�A-�}4c&� A a8�� ���T�i9{�r�h�o֕*�� -���C�����8$��ҁDFP]�p�|+�I�0̆a7��tO�hȐC�30�|��U�=�b8���Q�΍i$�CGɍ
i<��ꔲLx���,����B)L�HmÊm1֑�ٺ�L � A���m�����d�m�}(�}�vqR]�0�@���u�g��:�nG;�2,�^A��*�U�#ɀ4���	�h�к󊹾mGW�q�	r홎�1x�8�vd:fkUl-9�� ���J�4�C�jGJ�`�����|DwaI�u�W,�}�urr�X_X���~V���tN�T��Vη^db�'���\Ij�F}����c��BrD�;���i��K2v՞!8����m`c���12�;"'�f8�E�P\����L�B揌5Ʒ�Xoe� �p�Y*��'߈aD��6��҄�3��f��'���M��� �HA����������2��ȇȜ"_t~�����[�k!���Sm �
��.o"�J�X���f���xo���Q�dT�;N~?�|�ی���:�ɩTCM�r�!}�T3��EH���/�c(}�������@f�++Wk�����xЋg١VT	�v��e({�o�1�Aadۧm@W�����Ęޱ�����m�d��m�A��m���g�������ƒ�a
���$ ��9`a���S�[0006fO�Ƽ��j�k���ޤ,����%��� ���w����sw��~6[\�;�cY?��YZ~g�ꑚ�y��t��m���M@FĮ���r�9s��/���9��m��� T��},�p��=�-1��#����d�@;�h �L@ڊXȖ�iϖ帬����=���CϘҭ}�E.��p�nKלw�|�Ǻ7�� J���:*�6�ԭȅ���%팇�Q��k�Y/�I�P����n�w�0����_���NSx�>	�J�kR0z3ކ���l�2���N��i���?;�)�ν�W�J��'�����L�u ��N�f�e7�Y( ��o��e�{1�lq��5�`��\�	��3[�v �c�;�.֎�4;){Z�E�5���wCy;��b�����a2�f���d~:��=�ӿ���c�jܮ_�l��0��ܱ�V4=�F�9����;�(�4V ����8�{YqDV��_4'h�`�f#B�$U���N���x�/��进����2��T��ij�'V��2�Ҏ�ϩ-7��t���ptK禆�^��K4	�N?�W.���8l�D�dW���aP��b�"'Hh�)O��!I ;0���ZEb���bzf&�b)���}�Ja���U�>������ڌyͶo|h�=�҉Yq����?��6���b�XsN��@�.lȡ������ߍ���`����`�'������Ѿ�#`Ԩ����djY�Cq~�oI��4��َ�{��&.����u���P
�ό1�N�AV{��N!��C����s��G�6�*�I���QDs����u����c��N�3T�T���%�zrɌ;vXs��i5�9�y�˥�`�5ܙ���c����߆Nni��?z����7�6�g�h�7�L�����Gv{��k4��r���0��&����0D��6�R1�� �Ic�	x���Ҹ�Ep+�K�w��k���ōn�hJ�F#m����e�Qŀ���)�
�;���a�N�t#�H��C�רك&�yn�{������`&_
~�2L��Bq�6JJp�R��hX�J7��q+'���@<_$��xti��MΕ�������˪�ks�!X����Vl� &���fv�
�غ�J=��=�)����oƭ����YlvN�fI]��&:{E������1���w/(��Eq5U�m\bZN�:6ٮHnL̟��X����y�K��[)�&H��y|��Q�5H�# �s~\@>���?�N�Zr�Q���J��gRH$^�K�p��H�����7�e��JEF*�oʭI"I���1#S\^k��b�������H<����n��H?�/Rw�K,�*(��Zߓ�2���1�nJ��64��-zzv%+�t���p��4�B6l^�4�j�	�v���ȁ4�MY�Z~���2�hA�H2넀�0�o��9�~I�v)a��KV�2`���l���= 'L�e����*�M�cd�Y$Hֺ��H��o���#���� +�3�X"�u�n�Rc�Xi�s"��Z\*�嘸$D7��Т�G�ֳ�{���
�y���"Y�"^��q^��|��N0�rǴ����s\���z͊"��Ͽ� �,J��>մ)nyD�z/#Ot�O��hO�v�aM���-������^&����BVE���~��Gd����`��Nl�K�3r^y�@�{��D��B)'����g�	���F�� ����n��E�/���#?ꙟ�CYc`1�T/��N�{X�bK���e6X��!�"N��W�}� ��~܍�Mqb��S��$�r�����������5d�Zsy�Ͱ�.~8
� F��TJ�%�lU,]u���?�^أk`}H&�3<oP��ta^hS%q!�d}U��A��������&���α}��AD�|i����K��M����Ez*���_�$	���K�v������@nYї5.�YY9HP�8����� ��X�j�X�N
�se�g�j�՚�L[��O1i���4��	�{�GQ���
)]M�K���$)������R�����S��ܘ����'$�q��0�i��b����;�͵*i��j6�v@�����n��5ˊ�4!IQ��'o�-��p�E*�:poW�t�	�x���=��H0����d�}Ք�� &�s�W��j�ZÕ�~�S&k#�eF	"����Ĳޒߙ�7UF�r~P�i��봠����H6�4�/:3�_�;�?���B�{��87�id��* k��D�*�B�#��>�HV�����m��哌��>\���+h��K�$`�Z�f��:ǜ~��蜮ќr���c��/k~ͨ�����'��쉖8;��ޥ�<��f��D�~�;VO�
O �v�]{���m�^nB���
rW>֛��M�z�F� 3>�k����o���A^�8K�7�^2�J�ͣ�H�0��P�"C��3-w-��!f�9��m�km�\u��Q|ʝr�|<�Q��͊b���C9���+���\�8�zPi[��M���:���]��B�3ұ���ͳ�� ��I��ʓ�� 7-��12{ѕhX�+d�s���o�M9Ձ.˪�=_���2�F�؛��2��;��'��A~#;%��&4Y��v��Q[��MDnQ�$��`{�/<ƤS����W��+�E �B �����f�/aDm�p�v�ӎfl�,k�-�u�s[�ο�~�y� ň�Z�6�OJ��x�iE�*��<F�
$Ia)@_y�|�.V�m��V~��y+�"bq�db8Zտ&S�%�n�d�5�o>
�2*��E�,v��*y��1B��k������
���
yHk����x�Ը3�ʵQ����d�@6��2��Dh
dv�I�%�2�]��%��O���O:-Z� b�z-��fB��;��$+�|lҵ=���Y ��@�2���o}�­?�b�5y#ф]���`i�k����zq���r���R��6����K<$��Z���Ub�[_E��$��7��g�v5�9�1Y4Uk��P��I5���$xS=�4#� ��ܛ�`}`��n\�@wc�������6��U�a`��1���5�O탬�m�62�G����YK ?8�a4NP.hi:!'ZŖ�.�׫�����~S2Pfk��"9�g*���/�[�8b��@1k����Ha�@�7ڢ(��Rk�)P�g�i�c�j4&[0/F>��,2_i;h��C�����O���|�H��;{z|�@x��e&Jp��V�c��1j�_Y�h�T0n�={չO��闰FW���:I����0�\�k�m�%�"�מ'��
F���i:��Sia��$*�k'�+��S�����cpJU�&�S\y/�����H�dE��p��LN�蔘�eY�4a!yIz,hm��k~��$�[��P0�w�Aj�_d�Ō_y�z�7�S{��Ǥ|6�*+���Ov:���.��f��9�Sܕ�%ȿ��\�d5�AzȖ�sz��40�
�xc �++9B�6t�"�V����6u�]M~���S*�Y�c˘RU��EO��]�^��;p�!U�C���g�M�xW��<�C��8���ߍ�I���;'�ñ��J`��*��?e˪��+�#�ЄS��|nD�V�?v������c�c:���%��ш���z=?O�!#���/d#������2�ŷ�݃ݮ��FfګH�������l�f/�bT�q0h�L��m����'���(������}1�2�n�cټ*<���oթtP�?PJ(��7!�Fc�
�� ާ:�M�X���7f���ґ��6P,˴>X�y�w�T��V��漟/O�s�X�I=#�����aX�cc�����)G��
3m\�%������O��A�:DW�6Zu��{F����e�Jj�lp�el.6�C�k*/��	��<W}�Y�F#6a���U�	3�EBu���R�h�Γa>�dz]	Ҧ_��L�V��#��*x
7��J��_�Kc���J�k"*��������UK�� ]��^�4��}2hb�N����� ���ꎫ�t���b�?4Gw�3[�����]���P����ʒ�t�gk�\4�����`A��%�%��ے"Y�'�a�VV��&�N�x>F]��u��iߋ��̓]q�r��K��i|�����Sg��������:U�ɨ��ajω@#^����=>�p�	��#b�|d*�y�
[�i��@�=�{	k��uH�Y�\�I��gH�QlƆn����VM��4O���Q��I�º����v���H�&M�x��P�HGR�	��Znܓ7f4I�b�s��#d�L�]ܙ��Y�ء�Hd��!����@#��w��|�^OK3ǞB]�#�ł&�$7�O���M5�����4����[��^k�L �k�����T�����lzڼ�?x�UIS�<l^'6���-&�\6�f�t��KFm�Դ�� �M �UN��Xbd'��B�3�`��9~/�b������c���:/^��߶�	�x`��u�q��3��ί��1�Z5.��{!c�����x��̃�
��:�X��C�]�'�C��{��1��1�I~�L+�7I�ưd�'�������hUIuu�G	鲑�jt��k����S�X���%ʡ�Y��ȝ8����R��_��=�|7����@nRnjhj-w���H<�؂�n#`A`y��XtL��J��<~�ʳ� H�Z�u�s_pl�.�.���[�y�.��W�l?��p�#{�
���,��G��g��dﻙ$�PRבI��}���'��,�XiH��%��iz>P��˹D��,��'��Q�&{b��=!�M3=��"��~����ä�af��y���zSA}b��Bc��:Sw#��}���9sl&�Ѣ�n��w"�#�Ĺ��s^+�P[<Y����h���P,��#��렕�M�����k�J&��܄ MT�m?�i�\I�i�? �4ǖ�X�B������.�X���%�[[|���4��"�#~����� �{[Q���oC7�3��S~FǸ���E[�?��>8+a1�֢���@ݙ�4�n̆>4[���>�����L\ڐT��lGw�c[�3�q�Z��X���� 2s7�A�_������-����{A����ٞV����d�8�i��<E��}�j���A�:בk~�˰�w�����z�<�ͫ��Q \�!������}��-)��^����z~����c�w��˫U�d�R�Y��oX���\���}ee�&��S�[��W�O]�O~|ۼ���j^P��aNՊ�]�b����3�~��W�Ӕd{�浔�xa��[�EDì&D���yߞ���M4�r�ϼF�
E��9؁�'��G�7�cyo0͂g�*Ɂןa�S�G!��[�s��͇;�W�o�����:'�{$'�D���L=�q4#İy� � �M��~T�aAH�/�K�Ć���㮨��[�k~2�^�$k�:�c��&����m%x�rD"�q��p��q��ݥ��p������=���Z��D��nÈN{ x����G�Z�wS�bp>z̻�?[�*l𝅙$
�Af��i�+Z;�B2i�R���N,|q�~Vt�J�V��_�&�VkU�L��5��Y3�¯���� ˷{J�d�=�����m�+	��@U{�%��ݛc���G�+=k=u��U6��g
��6�O��NZ
t�+P���Ovy��]"p��Rk���|_�k�N��,�����2�"����`��p2@F�wOe��D�]i�HG8C���[���[B�۽���`��|�S뮸 �
S�nHe������YD��P>mk�x�2;�e0�����I�B�Z&ϰ��a
i%��w�!�_VD���2�r�Q��O൜8�����m2���c�K���ݓ��}�)�1Yh�§�\���r�F��Tb���� ����+"[��3�;��%�K����a��J�$=�~�z�,-����c2D^����E'�7����4�:aX:v���1q�YӉ��IE{���k�Pb�>+�y;d|8�@��Z@���9rыsp��l����Y�0������Z�e�\; ��&0�vki��ƈhs�W� HϹ�B\���e���� ug7�5������7|���u�Y�3�V�z�j�C�T��sȉ�)�Ci����SH5�wsCdα��}�O�m[ln�]����Z��X]��&�A�#ˈ1�W�3�<��0�	�K�1zp�?ӑO�@�[}��@���g��٫_�,���./��S��5Am�
�v)�E4�5�9��B��ڙ��r�'�~`��4�3��-u���C�.k��Ǟ0[R�7��'����=#H�1�{�)D�}��[�2T)/YH��܊���y�O��a�Uv\�aI`�>~��Z95�
�Ƹ�	�ε�g�n�x�3�/�+�q2L��%�ل4��X�?�=��`���}�.q�e�e��q�W����m��wܩS�N�np�?J��ʽ���#C -��2P%����6���[jϦ�]��R���"̾������e����� ��Un�*��6Bh��0���%���Ѡ��ISS]"u�S��n -kT�A'��Ղ���@�Vy���֨ľ�	�s�o?5`8�S���̀;�@p�Rn�����
���{Ƌ�*��~�`�Č5Y���|5���`�0B&ke ƅ<:�O��NQv����Gmg^9�HU�Ң��k��FW�ǒ�4�ƣ1L�?pж�<m�$��.�3Z������O�\��l���Nګ&S���Mj	T��\QM�c_���+��z��b+-X,�$Q��i�o��u`������/�%[�I�v5��O>y�ԅ$��NXv���U�8mk�5 |�5�8M��.dǓM��Iy*K��v��Q��e���of�<)Қ��X99�Y9�g�؂UXe}*�DZ���
�Zq�[K1 ��!@�oԫ=���u>
^b!9B��&3����ht�S��\�����o1c�Yq����jB#*ϯ�\�� �aH��	C�`���xo�7�~<�zhY�X�f��9���ކ�o��5����Z�C����m2�Cu>2}��_b���-h�����yt@�������^Bd7�bV{SY���DTS��7[�g��I���+ݻz֌U���&b_�j7��w���ZF>Hו����q��N����ۊhb�ZR O�+%���Uq��Kfd$(�U�&2��}�jR��1�/fB��fj��P䋷4΁8�V!�I��#��5��#h)u)�|z,g�r֖�m���xv�)�.�7"b��%��������ÿhi1K�g�4�'�Y�g�����C�$���f��,�0#ކR����L��!i��J�n�jz>������	� �B)4$���w��(��j?27��4Ǝ�_=,��L��$G�3O���EW��P�
������AjX�r��4A&ZԄvhb����
���>}h��E�������[1$qpJ7et U�$(��)L�������[���.�t���-�D�����CN���1,K�O�NM+"������8�Y����&	 �D��s<@ѓ[�������� ��X�?��uK�����<�E��tϞo�q�5�5���i���% �`V%�0O�i��	D/�Z����c�A��%}"�t� Px����{Ѭ��ˬ�7������̩逸���^Rn�m� �=�x��_��>�����W�ܝ��i�B����]�j2I.d�v�Y�yܲ(�?��Q�[f��# �.)�?�`���Z�	��+h�[㵶4z�{˧A������*Q�Ն2���+�iH�mK �C\<��Q�m�A>��w�k��?LzH���M7<�@���1�Ny�`��N,8��c'Yv7��r�����WyGd�s=�L|��~s���$+�E�+��`�~�*n3�A��M�ތ��O;�'�����8Y��^ �%����4�o
��2�j��x�L�Fm�Wom���o�:�m#۱���ǎY���&����
�(�̃!�=� 1���^̵�e,Rt@	�A��`C�:�D<q�=[�h~Mםr\���騞������nMM���EP��P���I�gI�}/�e4nQC~�|������% ���3�ۋ�_��ѹ���9�����C�(p�g��0�W��@�[�m��aEXEiG�wT��ԋ��VB���sF�]"w�����.�^$_B��|v*Q�a�� ���W���b��E�����f")��?i�S�Q��Ͼ���������O�T�>C���=����?�䂳O<�h��*���k`�W�U/��s�/�*�G�hVS;	�ߕi�b��sK.�û�N��}��Hw+�PJ�b�s��̫���[����q�";�;X6�$�_4ѷݝ�|�4�$�ژ�%�9�_�q�t��}��k��}2�Z�0�y����
5a�	�Ͻ�񈱂�o�#������NLvmhپ:�S�y�����%V�ĸ�+ 	fw�B i�Ta���)��� TQ9Vg���ΤE����rHq:*�Q����,��N����׍�l�����ƸE~�j�fʄ�e�Ȑ �.}�i��m`���	"�����B�W�/"����{s<��/]X��Z���SD@�/�f�(����^�ٝ̂�H�b�m�9�|�@�J���r�i���=ӹ�8�ֱZ*KR�.0
_�>��mb��j�p�	����⾭��'!rK�H�KC���e*���g+P��=�/�y({*�����M��"EG��Ļ��80EF��ڜ
���������%��9��1L����߫s�1� ��T���N��^������N�N�x�O����}�&c��L�|�ؐ�Id��#�}�}�~���R��]ܙ�]}��'"*��b2�&��?]Q����s�O<�Nd�<+s.��NŽ�]Y�ϕi�d	��|�vl�C<>[��}�
� R4�r����W��ޡ݄�6���G�R6NUQV�"�8[�ƨ�khP叼�.��{rk~$�,!��l�����5�T�Y8\���;�n��H�-r�D��櫟�b����y�����3�Vp�6���ض�o+�d��{_{�P$K�{tU������t2�����υ(�Z�;��[������\�"��ѣ���͘ ��_�#�ú��?s����oH�>@n�ԷfP��7?*��5�1��a�eO����.�C7�fm��c�ݠO
71,"7)j��=��l��R����E^��.� �v�D�tS4�q#�}�*�x;�Sd7s?YG^��?�w��2p=��c�ڬUkI�������'�U����X��`�-='���;��1�ou��5��!����� �F�j�"r,z^EG��#�?[lv���n?e�G9Q�]��s��_������t����f!D$�Du��z�L��l�������<�ŋ�����m��q�Y�N�O{�7_#�<ߘ����u���6�o)d	���vi^�H���$�����&s����t�<�̡Pvf���� & rN��r��ox��hx�����/�v��"����C{�|�O� i^}8b@q�,8���.ִ�Ѷ1�i/�֨%���;u\'i&n��n��nm�Z�"�}�^�|�8�W�������\عÊ� m����t��qٔ��.i��^��J�B�ai�km$.�崳�:�0���g�:�b����EK� ���K6�(*y{O�a��Wu�]\0}��Ȓ��t*Mc�g��� � �^H�	��gu�V����+}+�w��5oud��`�ń�DE��j5[������H�3SP�?�d�i���ɥy��?�6�p:t������V@D�=3|+qKZ�Cs��P�6�r�?\�ުlhaw��o�N����Ŗ]�A*>�P�{VD�b)�5�֪N�z}���hd��\�u��VI�!�c��Z���u�o���T��+�0;����c�����Oì�1���S�J��W��=PPf�^�g&����~������!آq�M
B#i$���?Sf_�~ڪr�7�<S�`=��2U#�L&��8&������V�U"�^� �x�#�;��}V���o���n��t�O5ׄ"���9���T-U������m��܋��6˚F}�'�S���Fv|�ēE1$�Ǐ�xI&	���T���4#��
��xWV�77@���2������8F:6��*����66��~2�v����Ӑ!
�h��s���̪g��"~���dS��7%�4�L�ؒ�#�)<�pR�ő��1�`e�e��K��uY<�AP�ɓ
�!�|�}g}�g/��/�8#
�Ǩs��[�T�����ܥ�{t�[��P~�X( �z�����q��F�K:�~]�L�|�A��r_�E�X�n���
��y��e��dy��*��7�rw���l�V��R����C�3����B���zBy���f� �;-gU�{Gc�|�2{�Q�߉O�}����nq����U�i>�z���p�IE����[��0"Kޠ|���ީ���.��h��D#:wz�R�(���s���r��U>c{��o�W�Ƃ���u�$7��޸םӱ������~x�C�s��٠�a{-�������Q;6��A��2a8�5��o<��DF鿳ׇ�?kc>n1b8�Q��Pߛ;���!��!�H;��z6~���ӃdF�MU�������hP�Nx&��U����3�j�����+�xa��%��]���/��2�4�}�X��'H2}����݂�3�}m�Q>�WP��{?o�S)zP1 f��J��1�E�����Q�r�����j�̸�F����~u�o�+��[)Ŋ��/χal�<���T˺���?���^�4ۜ��.3��X#�N�}�����E
4ܙ�X)�T�P5�Ex���yT�ޤnT�lpP�|��e�zgJw/'���I>�u�*���g��+8+���ewt�Q�Ϩ!G�_Rl�,�RЅW�=؜���,�;Ӓq�F�;��'����5����ҍp�=*�-ba>���:����sGŀፘ8%�	���wru���{���y�;�)?�e���W8���;W�-����i1����s�9�	Rی�G�%~yH}2�ԑݤO�v�Q��x�����0L�bW�8qzR2�S�I@�$���E�'�o��_h�,Y�#�:VA��>����8tWh/���v ��+�0��z��}R�x9��Hڦ���eN���F�d;	����o�w\t��_T"���3O�@~Z{��P�&ܲ���$���Z|� t�"��͓���ظ|�n�3�7>b�K6��H���*��,�0.j�U'����?��R4��Jj|�HR��jW����݀���#<ԑq���������f�t��z/V�h����+�N�tIh��@)Z�:�-�o������H0�oOJ=<�s�O�,īs�^�.���u�Z|�3�>q�|lP�q�����	o�`�U!���?;#�MQ0u�������xCZ&��|5���bf3�،��А���yq�{�#�9�(�$	�MIN�'	����TI��Y�ߒm�Z���Uf)����/B�y�Tݮ�����J�)��؞j�{�E�H���#Bȹ^�p����p�ׁ����mjЛ6�7ˎ��F��)2�ȥ\��Au�561��u%ycf�6�����S�7��(/���
0�#��ƥ���ٺrz�/)H����^�)QJ����N��W`�U�?dQa_%-���/[?�%��.n���X�*���
����Ѐv�p��]��+��a	�4���������h��`��8���j�%h?U%�h�Ld�ٵS��Z�;H9��j�@�@An�fԣO��d�@����
�Q╮�+~ c�w���E�8G��
�t�rx��+V�``���#H6DZ�t�7�.�|�N;@��=g�l�i��K��#ΉM�j	���Ӽ*�F���*ۧ�=ǡ:(��rH<�\cR��ᑻ@C�ѣ�E�N�qW��2��X����U�Y�$���_締cC熎�me�#tz��^.���	�q����n^�a;�ӈo�,���!�X^��,�=-k�7�g��:�,TCc�\+�VB���nnM��ٲ4��!-b���nF��KWl6���ӽ�XF�xe��]��i˕�n׺�u�?��}OVA��'m�<h�{���t��hA�%��JO�ٓ�R�H1y)	�y�څ�H#�+TUW��\�&�ﯓT�':1�]X}�,�܎�u�6�� �&�;(�7/--�Sd�����ԩSȭ�c�B�~�9 ~�znج�������O:l�◬�ֶ���ߢi!��5�
1���~����jE**a&2���DUG��	ՃkNu�Ԯ�]?*WĿ���R�vضm�_�V3k(Ғw�B�$D��?eC���Pη!�'<%���$�D�'l4�5e�~�N�'m��Lz�ڊ�(� fP��ޭûM<��)c�m(���倭_j�K�J�_pѴ�$q��S{����P}�o� ��hA�t����3��.{Ĝ�<���<e�+$;V#�4ʃ*O�X4�1����ȣ���
fBM9T=�<V8*>��*fK�#�������%J�K]�6?R�{��E�+��wY�̊+4�'&Ĩ�l*"A�A�!�՞��ڨ]lت��y����6��k����NC4a'�p����,��:���Э}:��Scc������7Ssp�;]��MB�|}�VI9��w��x�V �ӛ.��?t�~���;Q��>	Ћ#���U"/�x�<�Jn��b�9�w�<f�f?Ǡ�T�naSb\_�X)j ]�����E�"| �|tY�w�T�U�5[:�/k���sc��O��[��{��<�+4]�ޯ;'@[]�/8�[��)!��AA$G�ri��!j�!R\Nɛا�\"���lл����\�Sy�Odզ��M �eȓ��	-�ȝnG-��tWη =��v,��MO��; 6c�#�(�rcǪaz�����qH �`G�+�m#?3�i��Ӟ?�rS0����,�'�|lӕo�f�Y����DU�v����-}0��ʤ czמ�u$<տZ�:�ֺo�,�Pk��I�_����2���*�M���,c'j�,&!J��2ߜ	��]�U���"c��~V��N��f`���K.6x���=��Ɍ�J�B�Ԡ�]�*��BʁdZ!v���	�&�������!�	8�\әLb:6h�c����W�7a7b2���]�9,�-�1�jX��%!&�X}N�X���8A:.���1��L	�&��	��C�bb+���4m6
��&�"&�T �a>��ʖ:�G{H�]�}��c���>#GA,�z�	�b�l�P�����|o㿍j�D]S��~G��_�� :
�^ݭ�!�0����K8�[��5����Z{=Lc��u��碡�3:�gФA��c�=:N�1rb?|C���gW��;�xQ�C^#߬m��?�вDڝ�RE��:&��]R_!��KB47�Ȍ�I�[������D�9�Ar����&5�-�8ǫs����ޫ��k@�s��E*Ĵ�����g��S�ϑD�z��4���,���c��ؑXb�>1�C��E�ӆk��!��Gt_�xO�t)�]-��5������Y�K`I�I�O��B�J�a9��������=�Be�扅�e���i��o˹la8o��L�� U��������},���?��}���3���#��k���b���3������asc���j���7�61�3��ƺ?�u�=���R����a�沓�0����U�b�5k�p���%L��RC�;/B�}-�mr}��<��Z�V��Z>�ֹQ�W��,��EM���`�|�X��";��k���#��m����@_$��vbC�,<��"ֶ�8ۜ�ԯ<+a&�s*�A��#��.L^d��;������1��L<���c�m��C�.]��|�2 �M�9]:���Xi Gc�[W��pe�~Ʌ3��Mi��>G�A��Qt�L��j	�Z�n�6�om���8#wl��V?��&	�>$*cyCGOl!�ǜӈ�^��U�����?��W@˅�����(���B��C��B���|�~r�KZw?3t�M8�%N��C`~��Gx�ky;�1�Fʼ��5k�J���8IbK��j��.��3�9�lSF7���)�֦"�wI@jL1RV���K�R%���ד��|1Q�$/�`>�	�0����m�U�����/>�d�F��tcç
�W΢'6��PMИ<0�`�Z�l׌}q"��F�{k�~�^�j�A�(t���W6�v�7>�J��������2SGR�g|�����P����6Fu��3H�S����-�[*̓M�8�S��4Ra2�򧂮-V�m���`J*)7�]�t"ʈp��@ī��+�T4�O\�]��k8lRX���?sR�\yg�#���Z�?�`0������Ӡ.�tx�y}xY!X�rf֞A�tlq���
_����V��ΰn���<��" +�;1L��O'K|<�u��\�%t!&�n�;yo-�Q���k���]����7W�,��d�J�p:�$�KxӘ@b���lT(b�A������P㟶�唃w����X��S�|���z9MK�C�)��9�0�H7Ov��+W���.��u��H�@�{�2~l�<����g6$���{b;	�i��~>�]��y�Ɖ��9��!�t��h�3q\/��8��*W|`��H�+���ɠy��R�	�?��:�S�����(�ҍ�!�Lo��J ��c�Pv.=	�A�wiM����T�5eD�!�N-���Ý�u~�����C�Q��Y�V[��Z ��@D�tM<Ǫi�L�DUg��l�e�Z��dp�a7�p�B�l�&3�]nZM���*"�#�J7���5Vݠ�� bc�pP�Z�FN�k]��h0kl��w.]^C��L���ȡM8y�S?H�wn�n�:�L�6@_��Q�EV浸5�[�+�D�,���^���Z���KC6kH�Ep!{���Է�ׇLfC�H��5�1��5c��6DT�+��V�S�����l��5�Yp���ۤ�	��� �b�#���]
�����JѾ.s�H�}\$�ٽ�=X?��(�6"�V���h� ��
��/��M^crA�v�-pqY9��DG�Q �7%��g˹��K������qK��� h{[��G�hp�$:"^?���Pg���]ckԽ�_���%�.4�r�߃��ٖ\��/�L�֤\�
�?lo���}���@�d7P�\qi;��} 5��
�*�(6��ɗ��~�l��諡��Y� ���zd�{ܻWE����l��CpTs?8M<B����,`.�Q6;�f\8�A͝ؤT�	PӲ�|�H�i��	n4��m:�|��R*!:�=ׇ����n/�{O ���K�V3>j�8/"�}K`�c��n���\k�6���9���`;.���,�nyD'J\ٵ�g#7s�ƛ���(���.s��v^4�^,���6�I=���&���t�"��E�Pa ��fT-�5�^/[.m+��nR���%ГK"��{�4+k��,��'D�=�v�	x�2����MV�T�6q�[m�������`F���ˁ���n�\�C����)��X��
4|��i�@�"0{}/���bӋ��[����r,���Eϖ[�����m��o�ꫧ5��)���aQwX�F�aC�{�(��@� ���f�#a��\����3�_=s}���̫4�%#��̢D�
l���c��`��*>��ǡ��sƕxݍ�������G� ���Q����`����t���;�����s��Vr�]n���g����?:��z)pF�$c�&�-ߡA�6cp[
��$[�H��xɄTZ�P쫴Ϝ����94�G�H�T���u����+f�1�Ml�6贗WB'�"���@G�N�����C+���!֗��o��M��3Xt�nn�nx�]���{����x�c�t���ʌ���ة�?<�Y�]e׼����d��"�(�d���/��3���zL�qs1;l	<�Y�d�k���x
�Y��g�;쇀�6�h۫g&��iv7�&iWQEh,�
5<�J�i�9�ιR���p.Ŗ�(�N��ʵ)͜cL��f������P���}�'=���*A`a����� �ǔ�5�t��jϴ+ʱ��!����7wWPσ,�\����b�^�ŏ<�5�/��([�PyG,�aΧݙδV����jSˢ�b�AM���b�u=��8����	��Ht���>�\ʍ��g�	ߊ�H�?L&�m���ԃv���xJ�`�
;�O��9M
����5"U]UŝWU�/�`nKM�J�Nf����7��{��&�2>([%�6�����g� a����kj���AN���5\)dQyD����?u`�R:���@��0�U�@Y}>V���I�����[��?9j��o��cG��}b����:��7��k�/*8���J}�\��%�@�VJ��i���������|��cf�d&�����
9R��b�u�eu�qGM~>7#p��<e؈�sf�7���>�w�D�m�����Fr"z+�� 0��R�.�ֶz"�nTJ�d���t�L�=��t,moQ���i7&�9��nU�E��w0�Q��eXk��� 3�]���B��G4\ʿ=���[�>�D����v5%i��	���#�d��n3����^ˍ[o[J�l;nW5�������=i�/+
�ɠ8�jN��g1�m� L�1Ƥ���ɮZ��QD��\�v�M�}��t�v�JV����Հ��C>����u�2����}�F"�pZ1���Jh�Fؔ�a�[���
Qp���Ĺ<�5<>��UV?*G"���L�L
Na�} ���lx+�X�*�uZe���>�<!R����f7���2��&kA3܈;",�����Z��(�˩ø_��r�&��A�(�y�D!�����|�͈j���Ǎq 3���4\���Q0��T��KȃΈ�۴>���_zR�/��	��I�q�LP�
����&c���+y0^��?�yEb��s��_�n?�M>D�Z�P�V�t�!Sj�~���e��$��������������gV�F�֮l/I�7K��s�� _!'�[�H]�	I?����; �(	[�k`�P�C��|U��ʈ�ۆ��M��_z"�%������.���C��{���'����"1@J`�7��~����8H�2�b�Z��X ǎ5�xCL��(��&��q��ӡ�O�N$	�j���:1���x����h�#��V�5^���T�w�k^|���V�J�E�v�@󪺧V	�O��iNA�$�frᣮ���,��bͶŠ P�(�E1�>��c���[
�%���&�@��e^���K��\߉9O,h�<�+!�g�ŷ ��-☦.��">�9E������������#���*����"�p�_���ڜ4+
�X��3%S����o�K���%1�^:0!Z��N�SY�2$�M�%ȸ�*�x�oKVe�>���	|�ΒuwH�������?�/�`�~�_�b��>q�\��.k��[�>�f|�7&�;�>KRS�N�:h�5���*\��цQ+Z_-��HL�w�+1c�ж.�'M�殪�����@� ���Z�dr��:+�2�TNa��`�u~J����7��1��q�@%�z�h\��Օ���q1��4��HS(�O5ն�M$��FVf|��1��Y{�E �--G��.:���H߷DV\"���kj�@��DnZ�27�V�L���ƣ�\�r�ݾ���V�`d��T��5��a}3����Ћ^�;}���<�$vʔ�R�q�� �Aiql����雭^s#�Lՠ!@��2;{8�p.ם8��lY�{�2 M�UT�Hc
��i�o�X�±����ؓ-8�:c����y��� 6zEc�%ǃ�u$ #3��ï:�l"q�z2I�)h�)&����s�
TEFEC�|	���r& bSؕ4���r��y�]G����iK��yT�6O1�V-	�Ј�d}����z9�ջ����я߁�W��5�`D���\��l��>�=s.R�|��ɱ�����Ϛ�z�j�6��02 ��J��Id[R�.��vfk9�3 9ѻ�����j� =�6�a=�h��]���� l}S�D_QK�oq6؎�<+�ں�²�1�5\�n1_[�����d����9+0��û��	^�����)�� z����$E����Y��rf_7k��g�7Ky~��^�y~^�`�J��.�`�2��R��t�����FUr%U�+�&5=Ho`��'�<Z�$�m�"B؅	.�3�Y�n=Q;QL�e�I�ǀ�k�AL�?��lO��=���I�aQ0f�����@��x��Db��
-O�8��y��L��
%�5{���:�Dm_�������ϠN ����>�S�{�~��9��()n�4\��jV�^�/��t�nIG�ZpG7hz@�a���c �:��o�+�qEe\��<-qD�&g��%�M�<B'&����+�����6,V���$.C�X+��d���i}����\S�6����iHJ��rf�<��S���:��
��qr��!��P�:y�}����;�H_}����|���8fk:0�Wl��������)��Y������6l���W��a�֑!�2�yqy��"}�c��7_c�mU�<����d�i��1�B�%�n5���@��/��.��O�cx
��A~9������?hcr�,�КV͏�֤.�t���_��RD�ɐ׮Pԅ�9)C�v�`�/'�x��gE�3��+�D0���k��+f�eс��8���]H�����q5�$�p��U���W���S�e�^�8�+#>���)��th��M�t�{���:+ӆ��ۇb%�]h	i�1a��9s�W��y�����U�!>��ӵg(�u�:���a����M�#Dhw�xPϪ�	Z�/�ly�)e��5l��Dj�� Ȝ� ���!p@Y9�9_M�
K���u� �(hj��I��]����% �Qe)�����ٟDE6�k��C�f~Ѕ��4�Lׯ��Z��2�&�����[���e�3������t�:� 3����� ����ᇎhf��T�G�^����m�^F��Q��)���^��Nx�F�MQ��	]�����̶Q8^/D'[�ۊ6jb��RW��*<-ΧΏ-ϩ���v�"��W�\���'�P��k�dP�OQ �TW����y��>K�سdZ�3Y�5�k����S�_~J�:g�F&�Uӣ�oȽ�>쏣��͚��E��H쨯�L�&jVi9��i���׳��^��y�XK��5�#y�����_��fC�t%=[�8ܧL�Ÿ��p:�{��d���ây_�o�����v���b�[��j��~IRÅnVU�.9�� %1��?a�]��4�S���n�ڳJ'�g`#�E ���"�9���Wtve�%/�|X��'V��-eՆ��4�IC�	V@z=�Ğ�Y���:9�T���N�!1�����__�u�}~E�I�-(<B��l���[��`ZJ���z
���vȄR�S�M�#!&�\�����^oG��K>�����HWБ�I���꺆�Ñ��4�IE�5Y�>?m��ˆV��7�/W�e������(�,9�%L�8;�ս=Zp%�f��w�38�"����it7���[6U0����L_v�]v�@�9�Q?m����5���(��d���L��Z|��VLoRii�1���P�T��z`(��ޘ�Lm�^p�@�BW5j��qh{V��+����.�&C��Poe�nm+��U�� K��� �����%�q�u9{�w�����Ӣ�S��7�G�81c��-��� ��l�Q<���Ƈ�a�����5x�ۼ,��Ub����[�\��S�	�E�'mG��jՀ�V�yb�}���.�k���z����s�/�r�YP��'n������Z�8�(1�1����|��8L6�-�!��Z��k��sɐ54ť�Q�s�
�8��-��o	�w�[$�֠$��ZCZ׷�~��6X��j�ٟl��+ iܸ����Ѫ�L�� �B�#�s��X�c�ɵcK�1j<%��u�y��M�b��2�<��1G�.:��t�~d�ΡA�p�,�x@`������?���W-|��	E�r�Si�CS��k�i�1� vh�鞏��m}5���
)��-��y�9	���
����|]&�S,�궾@>����\O�n�	�-KF���ډ�_�Yt'}�א
~���ݦZ^J���WjH!�с�z�i*
�+dy���#�Dw[�S���*�ƦqǻI�.V6t�R�H��HʢX$?!wx~���K��s.��h���@��݁���4�~w�A,��^3��~oM�}ƫ�uY�p�M�8��hQf=%��q���`oA�T/�L��.�6�j�Y�܋ޱW��sm��\Q�E�<��Cc!��	!Y�rt��Q�gke��^��X�~%�4AsM���_���'�>d$����	�B0�����N�ѓ�2�W���H����g�[�d�����#M���tT�����*� �j*3�QGҺ-m��v�,���y+�E��?^ɥ�3K�ZfLh��CD�n>K�[���j����m�"�j]W{H-m�7�p��w�O�KB3ݏ�[M�� ����q����~dD���~!�����K����3-�ފ>Ł�t��$\[��mS���"HP��
����H2�ټ݊��C�hy�)�"�-�G�[�LB� r����@ة�c�ľ!�oYVI�Ƣ�z~3/Z N+���ńk�5'��ބ
�ֈ���㷏w��Cc���m��5o��?��4;x�?4��]^?���Or��ډl��e���@�(����$��Zb�L����ee�˧��UZ%43�
��`�Ĥ�vgtߜ��~^p+1O�ACM��um�2}��~�-iO&*�c�"i�xA��߾U��ӷdԓI�^�,��|�L�?8��>�x�����RXNXK�c8Y*7Bʂ�^�����`� R9.I���V3�� F�{����f�|6�=g��#��^���u]�Q�&D�Ǡ���Z$��{W`��U��9#�CR�QmJ��nX����	<��LH��m�)�+e�9��Q'\�V�%��8E�r�x��|�4�O$�k4TY����M�������g��^��Du�l����Q���e�v�`��_v�8����Y�d?�C)�ϐ4+DPv��1��,����w_�B�*dm5~mL$�'|����f�=Ƒ�!�-����L8 p3��/�Ho������j0��^C�Gi� O?za�3�!��e���	�e������I��>��6/�����6S�WW�o:~��A�85�[U�֌�M�]dM���%|��ۨ�!�l��}�z���< 	%��U�4Up�ڗ.Вv����:��7 xz�I�2���FC��\����R,9b
��Fn��^�� ����y�:(=dk��#�+?�ۀn��1CBS�k'^r4a�� �
3�$�؅%��>e),��GK��8��G�A�ً���"
&�����v[�y�tS���)d�%��o�V��TKOޱ�xJ��k��
J:L>���G�$�}�l�A�4�~M�-��8��i�]��s���}s�髂ng�Qs[�Wg¶��?ƿxI���{��}����~,�D(JA�<d�^H�Z휡�\�(�K��'`������/�-��OM���]�!jqH��1�����G�fS�;����E㈩��,l ͌0��<X'�.0+?'��P�`�lˀ(\[�x+��ml���(��~`\:�}�C��n���?ȅܸܖ���s?�0��\%ۖ���l��Vp�u"�:�X���kl�i9A��GV�l.p���9�=W�N�8�|��^����/򁜐�~��q`|��	�?q�Y)-��c�Vh(w�L=���pL ��[/5VM&�g�|�ў��S�ZjN�+��=A3b/ɽj,��W��:��G�n�~@�%ƙe}PHd���Y�ZDH��UQ��z[g$O��;QD�D!�bKe\��Ѧ��#-n}g8 8�Qhr���$P-p���δ��<ª E\��ڰ�5i�W٣�4��r���NkL�yU��E�y#�m�uBS?�Xc=K���oݫ����y�,������
�t�L=��+��G�l)�.g���2Ow��J>�<�z<GbK��x�!�ζ��,��+�8m���q.$��=��O� �d�u�.��pf���?���q�� HwD4�
��C���*��aX N�Nz���j�u���O�# �������s�6?���%\���\&��ڔ�����r���>JoCX�Lz�.����Ϗ�ꏛ�q�x2=��$�xG�&h���0j�E㷜8Φg�b��d�"�h1�9Y�_��S��\�ԗ��{Rk��Y�g���f/�*8��r��۵>L��OG=ŊX���aF{����5U)[~�O�,N��y��� ?�������lҩ��WID�qtr�g9D�τ|��l=M�k�\+mV�vn�G�y�X/>�'�X��бz�r��0��=�Ԑ �:cC�ɑ���Wx�L��Q�� �$������뜤Y�s@��Mrcx��ti�EE}���������;G:�����I增8�VF�@y�@r�V�<Y*�t�V~�7lQ�\��~MM�JļM�h�I�Mh�߷Y�JG]�z�ii��.S���Y���{�>쬃�X���pAq����բ���Z@���Z��CSE޼d=�R:؇�^��E{E�.�m�Io���e���ryi�p̉�j���b"�_�s�ni�v*���UQ^+�UԶ���t�s]rv,�%Zy̕y�����:^��bݴ5"=�����Q	�O�&� ��{(O�,	�Kx�O����Kn��Ԁ&��Ej2��l�v1�� ���v�|0���@�f�R��E�MX��;m>Q�-�:���[�D�<��F��wⴘ�Ylq�eR;W|�oe8y���dU�ƀ�6���6JDۧnxч�4�R��c�����ژv1�1�vK7��+(�$E
D�m)2��tX4`;A,��{w�Y����s���Kd|~� ���$�Օ�ם	����������9���� �cC���;*}3�Gk��ԦpsD��".[�V�����Q��+}<�h��O������mhs`B��8��X��&��\}U=�Py���B���H�m� V3ut�/ֺ�O�����#cR�^!'�hU��X�ѓ� r�D��"�6���!���ɲ�g�~�!��p��آW��Y9�_�������3���[KD�/��]>6ga��{߫�Z�_P&1��PaS|A�y�H;7�E��Y�xk�vG�g뮝�ug����\ �
�߭��j�'�}��?5�z��>�E����p�)����I��bN�`B�9��)T�Ǜ/A	*"l.�����)Y� L�_��T�Y7�_������ٮ:%�Lо�c����zo�\��]Xծ/�~K����Z��Kz
fO`<hY"�#y�U&+���kNU$�N�|{���叜�2�(ɿꟓyŖ@��A����$���t9�g�f��[��z6�A��7G�{p��P�Α2]����&y�CM�4K�6�f������Q�) ��}*U�mnf�@������7%FY:��sM�~���c^`�Y/�VeNEI��]�7CQ7/�z d$4,�ñ,��:2�!:Jݱ�Ff��u�E�v^�g~CE�8������1+e�&�'<X���ͦ�W����B�U���{�DX���Q�O3�Uo�(/=Y�iI������#����o��b7�Ŵu�F;I���{�׼��𝶒�r^t�ޘ!uϻB�jAe���b>}��R��>���b��?���sy�<���X����]�θ��q�MLL�9t�}�r:�������c�:I���=z�ok���0y��=�*͖���笁�����cH����LAd��a�̉'.}�9�D��lqO���H�O�9��:SQ5�~�q�gaJ�E����^L O�Q�e�%���F�i����ȵ��� Uv�(�)�K�����������M�芍l�E|s7��>M���CMH�́9��~I�O��8FM!ew�E�^��j�~�R���B��6A	X��5�}-v�¼�ߩNompԜCf�0�)@� �v�Wye}�/���6T���E�+蹾Pr�����`���[���O\�]�v������elR5����fGJj��m�*��!���(	5�ƙ��ū�nHN�6�*���B�3���1���`��0>lp<��xڙS������׏u����� ��L�﹡�	�M3 �/a[�"˚f+��ި�� ��7��z�c�.~��Pf׽�Hou`0"��BKV8v3�zV�VYI�T1ag��[��;�g$��H����� !��]���<����q��H�,��(��|D��
d*,kBz����8�6��_t��<u�D�> �����ct��v;����"t�I�־��}�z�ԝo�
��+���~㈽q'�yis@eW�#�c%O��q�����X�(]�vtmU�\���U%�*T+L��ڒ1ޭQa?��6	dL�X e���B���̹o#�������h9�O~�d��G�'�����'oV)�Ǿ2�<��3���!	��(-� 4��(��7QW���AN6��V��M�1	1G^
��� 桕})��,�1A�,]π rQ���,`"|�n��\�,���r��ڶ<'�b��!砩o�Ab��[�1�v�	�P���[Kx''��a��"��K��"Q��"5(a+C�e}ś����|��m�q���#�۝w�j"�N�K�Oo{b��� �H�y��^���[�L�O^���ҒY�}~��3�f4�bp}A����FebƼ"N �b{:����Dt/ĴJ�{am���.������~�F]��s�Ŏ���b��Τs6��Z9cz���W?�
>�5�I�pX4t�@2M��+�Ȏi�f6����C�.�����M�
�W�>���m��H^�'���7��H��o5!�#.XU���:Ej�%�Q�m�a�Y0O�<�=��۸K�^�i��r�J��cDК<u�ߤ�>I��~°�|�Ud��>�f�b�Ǟj翜d���)>EMς�M�bK� �≍�z�Kw�m �������V�	��3��̅Ur�_�ؤй;��VҶ{u<	B��v��۬Q�K%jF�(]����� ���U��l{���{���Y%}W��OY��G�w�|kK�%�w/!��;'A��.8~�w���t�Lb����C��AT�l�մ͸�q&R*G�LX%���aX7F�2?��X}��ipE6��6L���ym!\z[�K���]�A�����Hׇ���\��Xe�ߜm���o[�����EC*�h�ձh�e{c�aGd�mn���M�jJq_��nI�<I%Ҧ��5r�e��6�C�{���C���M�^�v��������ˡ�>]bc������;�w)�.�g��p���!�_xv�t`��[}�v���h�X��Oa�|&����Td�v���km)�<ZP���A�����v/j������Ӱ�禣�)�1��E��n�,C��0k�#擲��q�o���ܞ�判\��?���Lo�1���A ��=`$"�]��4W��.rV3奕��6���E������#�� �tG�+-��m�tNX�8�$:ٕ���s�R
ՌA\u��}ܤ�YSwɝ,>DPԠ>h�do9�޻#�qj��An�@��x(hQX�8U���������N�\S�Z��6l� V�@� S���3���y~~F.p�!�b�`	��P�ԣ��P�&Ys���?�;ڑ�xCQ�uF�8qR����i]	I�����k*Z�5p�����X�
��HW:mMw&��#%k�ƲE�P�_�~�a��N����@.�,�m _�?%��~I�'��i�g�Tޡ���$ɼ�n�G�:4U�w�)̭��b�ҟh�S,#��%���[���L,��\�/�r��[L��>���
�Y;C٪�	�	%�O��P�f������/{�1�ؓ~�Y�)�S��Nj��C� |~�}��e�z�jm�"N*�X0�=�� 4E��iF,C�h�O<r��j�V���D����~n�Ix��W�:& �4��^D �38�*�0U	�]�A��|@4/ļ����7h8bN�����G�C���������o�n1W�{B�L1G�3{�{]-�!�/���h	�:����1
�g���ȇ�p���M/�e�I��d�6@3V�ի�h��ϰ���v��Jj�}��х�Ԝy�u�HŘ��ۄXg_]-_y.��|����� �0%�5q�=�������⨺Qg@��kI��N�A!,u������Y#���x����V�hT��,��h�W�	9�V�� � 
Z}����0V��PfR�t2���	{����O�V��Ɂ�-�O��mӭq)�R~B���.[���U���ci�V�!B�T��r㊂�⬐;�fq�!�FrO�(�M���΢[�]&���C�9�^�	��4&�5C	���lɽbi5E`eͥ�>v�;<� ���	�����cU8�������;��4��T�}��!��dE�09^�k bqmG��H�n����"0��lЅ7kwU⾳2��%Q �W#���s)�,/	�h�3�"��t�n����.0AOǍ�bn.���ǥ)���� �+�[n45U'�"Ȯ�I���ayHf[�.�1j,ɡ�<.9:�o˃>��N����(Ĭ�	��ҹo,��h���y����"��)��S�ӠN�����#B;<���7PH�P�����+�#��'�U�R�|�r�uh3��N�N� u�rtqX[��+:_Dф���b�U��R�f��I�sCkª;�↸��-<β�`�)��eI/ߊcd!,|u^�b��=/�������L���x�3�C#��[6Ywn��{<s�P��;|�6\t�"Ώ{-s��kO��&�?IG{�K҈���
���n}�;����An���6.��g���2�,x��?�u�"Ɩ�&�������/a���~2u�EǨa����4$F'�i���n.��/�|ٜ
�+��^MEV%��z��N�"�k�+܅k�� w+/,l���t�8������5 X��Gt��t	~������N�L �B��W�W ��&��H�Շsw��]o�څ��R*0�-�+�9(E�����ތb�ն�d���&�lm�k�ޏ���؉���&@K8ydW#j&l"ܗ�z�%OS�K^���)���a��s����վ:p\�>8u�i|���z�0�z3��<{g�K�9���4U�
�&������U�k�L�+t^�U���@�$/NGTN�����O�����	�`a<r`��Ӱ�/80�xՋL����t���P�C3r�-����[�2�ues�&�]�7��#?�j���G�扳nA��UN���N�%7��|M�t#�_��ۨ���f�	��߇�0 I5	9��AK�K�BR���dn!���:���֑/ 
Z1��;��t��%F�q�����;�N/���{�̥ ��[5A9K��\�M���F�����)Ć�l�s�M��8@�������i�^o��a/�5Z\d�J�u��"��d2����������$U�r,��������ڸ�%�!�D�@����s�r{�/�Ǩ��|D�;�9U�_ʫv�F�fc�����]�ԍU�S���F�%!��y����IA�'Bߢ�؛�
}Bz֮����;+X7��7ѵ���&��ꀳ{�ĎQm&5�?}�hÓ���LN	ȧ���c���x�b�dg���� S�Ea���E[�M_ʛ�I�}�:6[��L&�!wD�ģ��%	6��-���O	J�V���^�S	(�|����AZrF�		�B��b~<��S8�%�z8�=R6�e*h���Ӛ}�{�j��7kp���e�W��,N��G�����2�K2�n��嬖����Z,D���E؜�?���#����JyI�f��.�Tu��U^Ag�$�׊�30��gC�<��j�S	/����L ��`�ګ���\	�ό.�|baՓ�je�>D|���^/T ���w)�+ؾE�@��� �Y,@�6�����O�(;�5*�?���|3�|;�}E�� @���A���m�|�: ��e����1sWXd��,��s�'ݞDP7���(R�����w^EtG��� ���ʙa/�"9+p���мG�SzdyK�.�<�v?zN{o�գ×&nԖe����ױ:>�(����}���[�A��m1O��hVyMp����RZ����_�޹.qIѕ��~��aJӊƔ����Ƞ��Ķ�*W p-�$pǙF��"�9�N��!K��>�}�a�h,Y����;�Kr<�s�/t⁊e��I�B�%a��*�V���b\3�Â�����E�/��A{Ŕ���-�k&�+��.Z��9r�V�/�f��ǆ���OV�V�'RRH��R����+ZR��'��|zr�@<�F+���d��/���n�V�Ը8�j�,�B���Q\��ɒ�*��Đ.z'%�Ӷ�P�m���V6��nC����M�G�P��� t���5ف��(u�,$?!���c7Q`s>ouֺ�t'��іYp�r�Tm]�z��\���M��'®|�7+yhN�inߢ�"���W�f��c��"�KYěi ���ߡ�:�LH@��*>���&S�Ǽ��)t<�����1y�FW]�Gy�h�4���^���0� ���F	Vw���H!'���g+��v�E)��yLp�`M�eN�(�F�<�g$	Ҡ/V��W!B���Ew��E͓��{REVФoed��þ�uP�4����,G�X_ ��:�S��+��R�8�;u�0|`pn;/��?���<ķ�S�!��{��6_�$x[ѿFKS/� ,����SQs4�@;������8��y�~��%U2l A/���|�o��/`Ң@N]�Uê��%�QBX��z�c_�~�~��28*�H<��C���L�V��!�5�Mfz)UW4VWB�X�w���;�?���k�A�G�����K�}�+e�|�'摄c,�;�+�
�/|��v�h��p�0�Bò�<��(A߽ri���PV��d�j�,n-N�^���(Wӕ��z�؊-��b�����p=�J��Ϻ���9� f4R�3Vɣ�J-�Y�c�����@7��+��|��a�Y����W����}S�V��p`K�`�}E��T6��W8���L����";����Ԫw���%ʹz;��!è'?b@� �n���o:o���p�g��|!$������j�B�Rf���H��#fN'���26/(u�=�o�?_/W��B���&6��=�~���Wz��E`�W�T5����c�Z|��j��R%�;�-�-�*[���"���ћ���~o�A��|$hfrE�/�l&֣V��c!�`��M�ܡ��}��� �� �e!ZR,�����:t�������ن��C���_���0������7I�����'+�P
�����a���<�p���S���rm�}���jy���!�"&4h̚��-H��Z癠!�����5T(�5z.�X0�R��C�G���G��G0�B�0�'�Z���Z�l�}���~�&(���mR����YF����y�h'@siV�7Q_}Z����6��V�7*U�(�BaG�tL�J_�����U�	�Z��/��>�O �MW�o�x��_��0����yg�3���Za�0$
j�2~f�V�0(�,I� y���E�7�����}7�bx�۳VH?:�tm�y	�&D{CZ�e����#G� ���[� Tpm��"�ƽo�$K�L!�tY�� }A5�Z��ڜ�I��F�l,�C��x��{+d5z�c����sk��9��9�褐[����i3a>�7L��F d?�t�����C�@ۮ��EN��P��ܬ�5G��a"�|����d�U��A}K� ^����o�k�k[xu��;���\�/h�Z�����5��*sNm��2��5O�mG��p�e �W
P�=-�d!y���s���FƱ��Oc�t6cM�\jH������p˓�*���Fŷ��<��ERN)lt��d}FWV�ŋ�����b7�~�H�K�Lc�����$湆���괅\;ew�	͍Gq�xmT���.'e����P�* L��*�k�YŀܶN,�v�٘a�Lҿ�~u��7ﻔ�n���"�r��{{��ckΧ:�Sd%C*(���jS[����n�~�aW�2z���F�`�y�W�@PJW؁���$_�k�w�/�'-�̍�O�z�5n��"���.��~K�$�?imA�����qa�5��[3����Xccg&�wt����5vS�R1c�r��,a��Lʹi2؍�Z]Z���G����\���!�$��t��������`P��ՒU(��+=||��+�3��.�y�SB@(@�y&TN��ĩĨ���G�B"���kuB>�P��L�G>A�@�,d�ɇ�_M3�=6c��&@��M�L1�������_�--��=��� ��g@trz���-So�G]Lt����$�Y<*u����G#F��q���bըO"��d�����??�Vt
֤N` �U ��Ȏ|bt�ɼ�<@��G��to�?YĊo��`onqL�iع�~@}];��X���L������>a�~K�9y��~�q�&* /wُ�C� (G�݄e�PF*�(���C��$2̒s��A1�O�`Ҥ�ۜ�+��"�z���< բ�F	�(���Ƅ����?	B -��uFn���?�s:��p��)o�	�6M�8p8K��4��=�=����'���2Fj`i���{QQ~堡F��ۺ���E�h'F�+��ɢ�ns I/�h�ݯ��v4��>����و� a�l�0*Z��N�D������H`�ۘ��G�`�m:�j��h�����e�  ��j�)���é�"@S�#����9�uÐ��4FpM|���H���w���{^k5	��`>EX׫�h �|�����?T47��6>��ٷ�?y�[J�R'ɿw8����ub5+�X;�|)��#'c���ϫ�R/�ί�o��E"�3�,̨�6�eԲ���Τ��i �\s0��N*-
�T=Q�O��L���:�<�(f:U�/eƜ��#�4��1����u�cY�5�߮��KK�Y��N%uo
c�`;F҅��R��Z���{����EU��/���œ��Z��f,�\��������_ǠT����.��+&��R�R?�E7L�_j6�;7\�gD#�n�Q(���T��@UA�_����J�U�=9��)�:r�Yp!bs�Ȇ���W�qhr�Y�gͣk�b���Vk�sr�c�������~:ɦ��T��uq�����fJ���m�7u�*g����:�	kސ��ihX����p��!��1���*Ţ�fk�WS�9EC��e�*	S��@�t� ,�'�bn6�i�� �ag��g,0�y�%�J�$���!f 
�p�^�D��EM�9^J�BX<�%��A�P�e�n�V
�+�Ƈ�������kY���"����n玞!3C�l��Q �S?/�;�e7z���Y�b�K�n�Tj�j<�/�*�QR����A�C�j?�CR���F�D��) eXyq>t�O=|˒��(�?�S"|�?��ʠ�$4�%���K�xrƲ�I��e3
�P=9���_�髄F�Wը��g�:�G9��b��0�.A�Z������6 ����{�pm��I�ȨBb�
���e^��� {��K�a���Ԫ@�������tNV���0�-l-NL����Hxy:4ԩ�%���:�1�y����!N�c��&��J��%@frn�Yv/A��kz(��X�#(!:�Kj����'F�W��YG��E�$f(�J6�L6N�4XJٹ�?ߔ������k_��;S�`I�U&���"r��[#�u�(�w��p�S�T���LvB�>���AȄ��o,�q���f�H���_5g 6&����@��BI.�";��QN�+1����e���v�^i�r�Xz�}�ٹ��/�ӌ`��Q=qH�{\�/29T�'� Ѩ�RI���-���BZ��?���y�b�z	w��#<��[mͫ�6��8����׶���G��vA���o&)�vf�D�f��{�2^�Y�z�OL�?К�V�o["���b��L���e,�a6�j8V�8d̋�>�̄.B`ȟb��Qh����Dj��8:M�õ2��çާ!�Y��'����"P��m�9Ŋ�˚����.������!���I4�Խ�h��&s�x]x��Cd�`3��s7�=�^v1{�e.�/�~G8f����w��ڏ>� ��O*��~�yo*�N�4;����W�xxS�r���\�<���spc�k|p_�0�3���u�^�^:-���ftG�Uas�����O;M~l#���>C�!!��,���?S�\���4� �x��b�o�r�����?���DdY��_�	8�=T�q~h#Gš�R�-SL�_�"4pگgYJh�G��sZQ�Ӿ��a�_sH�0�i��m{{�*���{�Fj�2����"#v�8����Cu	�hb'K�����,��L"\ID%W�QG&507�����MG���6�Z~�a��/���6���˓��@�9��u`E�5Q���v�Xw7���R���W�����UN8�+�a6(�ʓ�~��)�SysuO�D�xI��,i���7��,h�5�qz, �L8�˃�H�s�R��F6*l�nR�<T�*)>�F���x�w������>��}���F��!���K ɯ���%}�>襅�l���~�(�ӠSȨ���?q��px����2����S ֝�q�7aS����&����c��A�,���jP���{#9a�ےE�]�wwH���P�L�4HЦw�|��%�ۉ+���^��!���p&��"x��y���x��}¾uM-O��_�"a2���8�=+X���� ���9��H�^�'��j�h�}��E����BG���;*<qU�W����!S�6�Ĕ�i��Y�Ȥ��;ed�d��*�&�ˉ��M7U�H�+��e���� �N�TT���m�+"�s��W��;������c����Kg!���d�ѓ1M܇��}����AA��^@���;e#��Vc�d׉"��.��#��R�N����R��a[(Ċ�b>����G���jN�,�[���>��5"�pO�j�7!��M^�^�۔��kr))IQ���%�6x�J ��nP�rD�L���#�t�gdU���%�6A�b�<�VD�0�YWm	���7!�8N|��]�{�R��� �q'ʰ��hPf��[�����JoZ����/�� �8�0G�p.c���� ��_ݭy�r?�<�qr�������IJ,���I1Et5)�JΚ".8�66���z��9�����ћ��wf�lU�A�S��J����,'}<����s�8�9<�Bg��1�R5Zo��PI��>����v�9�a���úMLnV+���mT��3�Vy�u���a	���[�%�95��ew��������)NMDY.�O�d�!Ă���!���{h��&�(��z�����(��$�^xK������z��ӤFy8I�$ş�������(@㸥��#N�� c�����6gv$����q�J�1̪ �L��W�D����G��n"Z���Ǧ��7�nV�����������HU���/��J�t6���ߡ��o�z�� ��R�����z��4d���`�p�����T~u�PR���Y�X����N�S�3/��u��'�lvD��[�� ?B��#	��}��� Bd�p0��萯���pt�O���Zw%_��ȥh� ��<c$S3�tZ���ĸvx�G3`��[/��}�xb�S��o➃\}o�Q�*A8�ہ�0���{���y�g&��`,�E}��V�ٍ��u����L�\�2|��4/��,3c�^��f�`(��*a�Ԩ����3fr�]�d~§��������n��|	=�+x�B;q���~���M�qU~nv-*�|a�K���/4{�\��6(��y?b��/�����8p���~F�c��n2L����	݀�{���ڛ���$��晴�\9�q���=1~?�8�-��(+29�`:5�NA#e(JY��}�_�H0K�e���(��ݛ�*�U�����!��J�I��4S�}��[}�[�s*� �iT�,!�����B�+R(�g��AnHT�{������r���jh̺����&��!��7�^�|� �}������g�º��[�ſ{���8_5���R`�֯��ܜqk�19����h���.�	�����v���6����Z����D�.��(��퓜�t-�Gs��M#9�A0���M���qc#k0�����3]#�����nU�{8U����6Цɞ>�4í׺|0��۬�p���[ZV�tfSJ��x�ްW�?����{_�$r�޸�7�a[���s*HᏉ�������1�H
��O�-ݻ(ܢYk �-L[Ys\�I&��j��ϩIE�}����L�n$�mz��a}�(r�粋P��ڀ�N��J�ģs!�l���/�0�e1ƞ��&1����D`kϙ�����	�=��T�: �����8A'���C��	�'�OJ��F�qu%��*��l�0L�C�.���!]���żW���q�R��E�,it
5��o4��M!a飔���$�V����'���q�ȜoM���}����J�F���ހ]O�6�m����N����1��w6 u,�f9?���qw6�3�m����cv�[��+a(����Ϛ,ݧ����2(dc<�R�ߒ*��#ݎ11W��$O�8��I=4�C�H��XϤȠio韢��vb|>;=3��Pw��1��="��������[dcU<{�_+�>yыL�(AW�i���� A�3{�i�� �g�6����//�'�
�+�������^�e�՗Ə��p�RV1��VVf�CV 9�.�`a�G4����G�R f����虦B^�g\-2�ͩhŵ�F��T�u�0���(�ESE5��>�*�^M��wH�+a7b6�Rbf�}�v�<p�<2��{��V}?��(K)^���si[�2Eߚ�7ݤT;�_myh,Ż!� �j?�!ko\t�Z�Kۻ���v�{ΰ�%}{�mw<�pJ_���k^L�t�AK%�dI�16y9���D�<���Ze�����\�G�\ȵw��izgW�R�K���e�b)�or����E�Y�_��y��u�c�_�x�+�%W��gm�&wn��ʵ���NL�sQ�1c��c�*ࠔ�ْ=[|(�&�&��)���lX�IF���z��o���������\vQ�D/�n�Ȋ���M���&��6>�-͏���qlJ��5�zz<AU���xV?�ivUD���:�7����f����O�U����n>p�X͠���)/��*����n��V�S�����=O?N���Y�BO�U#���׌���{G3� �B�&��i�н:�_��$&���Ҁ"r��L{�+x��L�n�3����V�o ZO=�r*mwǄ?{�Q�Rݴ_}�2�&wۙ��qb��@���-I4L ���}䋂���Cx��E��-gn��g��3��VT�뒶����tPk+��.[���źz'�à�씕�&'.�S�d�袕TE���\J���������������XD��(��s�D�.�g�q�!�CZ������zw�-3&@�a�)��Nfpi�iKsCY$��	w҇�+퇢w��m� ������;L¹b�e�����E�t�fF����������?@�~6)`,��T쟇	t�%ΰ@^s�9I�|i3f�>�.,���|�'Q�ޡ`�����hg-w�M���vT?��	Cki���K��m� D�(x�4����@{�jl�A��"�e�������B��&<Rah���w$������E���Y��]��|���HP��֝D���l(��f;H2��v���i�B��v莪�׃a[�#�L��vhsn��!$�\Xu�j�
S��~��?�k"��F�pV a��!n*͛\p��(u��ck�Nm�������TJ�F�Ǵ�02 �����a�x rx�W4�;p�Ga(�D|o�zy�k$Au�_w�����Z^�4x���y>l�@�ΐ��s�<�R���w�����!~�Qyo%���qA]!)�Zs2o]�-�W`U���cέ�fot�w3�Bv���l��M�4��O^Y�1�`�2]A�����"G�w*��]��_k3��Yd�i���g�Ȝ	πf��������2?�T�8#���`^*�L,-���@��D��T�gp��rWgL��^�m��,���5�e�o܂�{��1��^����S��p#z��]C_�M���'�Qj.|b7I�>��*y\�v��FGg,9�.5t;�>�2�κ�X�>=�ag���zB��ʹ�p�J�m:<���7�hЁ�'���j[UY����R�d�a��R]w(P�c�V�zj������=��`��`���{�}���c��f�AU��ǎL_r�S�Pp�I��4���V �Fn�9|�V��⌗9��A�G���x>��(�}�m���-'S
]^�ɐ�$[���L�:uh�
�0I���牋��������R&;	�D�5���t>~8�G}�s�{lݱėxt�1�_�Nя�e�	�G�k#�l:����^��s+�$cb{@�r�*ߋ?��E앺*�)ׅL�@�b�����ƍPG+ݽ�8:�p 6fo����e���Eq�~:�8��V�����qD<��n۹����:� A�g�0QX�WN��.���d��m����Z9�J��� =�̼%i�$&��.��>s�AC/��_�:b�(����1��d��w�\R
���
�n�U\���b�*�GԤ�b��0�4�:=B��Ѕ��������q��bd��,�*_K~P�������L��lC`����!��mD�W��,�^��3�e�o7b;�E1\]V�F14�_Z���,��o���Ɲ�<�#�ٓ���g����)v�9�Kɹxg; ؘ��
2j��\�Q�����w���*��n���̹��P��|������o�� vD ��`�ғcs�Q�ݧ 4t۞,�i��ٻ�C-��_��E�n(.ح�qk$�)��i�H f��[�ʌ�n~�� �`�e�ݔ��m�ʻ��Wh1����D�����I�+W��pqE�9�3���HeqS��;���[0i,4�ݑshx`��7��>��$"mIH��u��8<���;W��7���`�{��?[�y�`.��7Źm�A���A�.�Q�a���_\^��`I����[�����̶� ��d��=��"�~k��Z삱�t�]�r�v��a.=_¹s,�B9L���c��#�|�7��ͮ ���Ã)�I�v�;v���\Xd7�9���W����w�@qZ�8��s&�|�F#��ӾuX���/��9�Cª��X�`���!��)>���%�ݜ�ٙ�kd�#Qp��l���U�� oB��?�|��gR:�z3���b�k(��7� ��������t��4Yv/��:�* �Y�I��f����pA#�@l�0��`(g\0�wW��f@�9Q^S�����Az4�^�s�ofqz6�f?�!nH�w�F�C�j�VM9���{t3�2A� �R ;�$�J�@|<��Ks�of|�(�`}���Z] A'��B�E�ĴL�-�wi�1�}�J5G�v�}�Η���� A��;�}_ܦ�6z�	^��SY�UZm����`R�0��γYF�#$�ZN�g�.>��5ܵ�O	����A���}��Ab������o��*�m� �����.�-��զ