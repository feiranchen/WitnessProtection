��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��x���y����H�z�������'��y���m���$�d"5�J�ᗑAë 
� X��I��*��OV�����Sl��)\ w0Z��'�Gt�XY��ƿ}��ڎn���������~�X��G9+�8�-<�Uc�Z.�)�Y���b�����N_��U��Q��?�W%�k\�x�H�7�|�\a7 �!�����ˊ�ġ�Sa����*3��-"�����#�NҪf� k�)Ӊo��bg�[��ld`�^���ҽ�S�4�͍2��v��Vۖt�V�� 1�r0+�u�A۳���	+ߘZ�F�v��uS"-m��/�w56:#Qª6bզ�o�tt�|�ˀ1���u�\�m��$��;�L����jt�Y�{�����_��`�m6V�6kD�6)�rI]�Y�>3���?[���2����!��
�[�_D���v��k����������3�`m� `B�b??�br1ʱ����?�fT���$���d� S}�8x��L����S�b٤�b��d���mLo�D���w:O����.�e�1E����-"��A����Յ�0�)�U�<��M{����5KH��y�ri=|��+ !h������jN���`N�T!�!纇��E��3�?�@ "Q�nؔ.�͜JX�D���D��J�ή.��������#*���j��0G�I;^&A�\��aL� X����%�_��P�9����l�QofF�;������i�>���s��T(�v|�|Ij'r�S�-�i��$mmC}ے���o!�:��Kǀu���"�`G%��J��l>�LV�ӛaF���>oh�Ͻ@���x�5�w��z$�I:����씸��#���a6���?$Q��NDY�Y��b�XR[� ���"����%~�K����J�L#� _�O_�6���ọD�Iy2�ih�Qz!Q~ ��{�4��_z�}�`VC#�=¢Q��k�1�F�$3j�9|��x����'�X����dP��S�[�B�?l�VA�|�!pj�.��&wњ�TIu��A��ϰ���k��Fׇ
�<R"���v�0��2���?���5}ӭd�"��Ca�Ux�:�! /K��Yim�z�T��zmO�HqvZA�Ʋ�za��x:n[2]T�-���J�o�Kki6o�Lc����z��p{H�|T��W�5���e�z�N�/�COj�坩�J�;ϫ�D��P��5 �;-���uᢉ�mWV�dU�L����A�A�c8�ֺ���"T	��:sbo�4���9�4g�����.b��/��㒦�W���'P�(�~��z<
���8�_�4�����cB��$	�Y@U��m�r�|�_v�j�*~�x��֪Is����Q?+�-��7�₅8�0�:��R�O�2c��v�a$�vY25G�&=5�"�V)�����ڜ��3LF�{��v=Z�C�$,w�?�
��NF����w�[ʹ�i1��-���s����t�z_�#��Sc( s9u�'�Ş�R-����