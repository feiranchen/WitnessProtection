��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\���=`x�����[�m�r�WPp����}�'�{7r(����3=~aо�~��ԢF��*���o��/
���m�Z�׊z����a�u �js��
?�4��Ry�h��W1��S����Cf6n���d���p��'�^Id���2AZ�����Z�!H�H)�P�;L��*�9_�y19;��.zX.&0R �&���T�n{b�j#h$25A~.ɮ#��D�Qf�?��:����; �F��ʰ��1b%�	����|��-��'�/O5����w�?���S�%-��C��L6�r� ��J�|�r��E`�%���E�[�&H��	ĸ"@��o@����mc!�����?�$�t�<�G�f+0:n%��<�o�����He:�v�3������̻# ����Ep��%�S����|�۱����4���{;q!�fFw��ߍ���ɾ������bEl�yЧ���w!>Ҵմ05ٽ����h��{Y�^�C��I��b�O�u�.������V�����P:�+=U%V��w��������;�n���d#S$)�ǆ��G��o.�� 93RY�J�4m��7�Ыt_�,$lE��]:؈���T={"������H�u�p�2N_@�ל\�����6(����A8E�9=��,��&���*r�M��*��.�Ef�����9y˘����M��X� ��#@b�G��ٳd��m�k�H�ŗi��h�  �i}u�n}����pE����\==��L.'�gѿ@5T�����[�[��t��[���ѹIJ�'����vrK�Ȁ��
��EO�A� 8��S�<Α,ً	̻����C����ꩢC��|M*繼��
8�UnO=����%��"�w0����6��7P���V�3��I �}�34�)�F�dّ�K�
�n���(��9����:� +�g�ّ���K,�^��ɋ���^JH��ۏн�~��	��'����F��|�sm�N��'�S��T�A�N�"��{�빑7r�.Fbw����(r����[H�.�	ǃ5$�x�/AaEj��LfG��R�R/�r����'��c��H4�o?�3�����e&�!�C	9Oȣ��'�ZXNeu�;��0�C=;f��X-��P���#F^�ͮ�>:-���Y�����o_'X@����{����M�V�ݥWYQAg�a���z��{��JQ�!HM� iFs���
��M��A�>��q:5��)�Z�i7	ِ���7$`�Z�qq�+�><�b��s߿[�ӌC�b"_Be~]B�r�a��x�-X�\ד����R&bp'��ϊb���ˤ�U�R��ѹ�nplD���3+{�CѽQ��(e���?�	m��M�,���=
9��끉:�C��ƛ�k�+��OC�� �������o%a����j���x��a%Ne�d^6�b;7���}��X�S��f�����Q���eQ���+��������g7G�S~��㔏�eF:���=W�-�2�R� qR,��g����y�5���	rdl��3�ր8B]�D�+�ܫKV���Dtv��?)[�ʿZl!M?
����n�N<bF��<e�툩o�d$���jݗ���o�� 6�rW��� /T����!��)��1ג��i�%;�d�����曉r'�s��Qɀ�,������O=81�cn��K���|B`��S�g��������y�L����i�����P~5�Z�E�`�Q Cm8�I�2v�7>��p��@J���I8�qq%�>��C,�6�z5������DysqϢ�᥻ͻ����`a�rT��Қ�w&��&�����((�I>��#T@�M�O�)^G��d��9&Qo���L)3纃�P��˲�z�+������F�pQK�a�BOM��-�vb`�8G�j��&_I)��Dr�	�w��pF_��O��a��G��܍H;��k��X�,��h/_wx�$b�X"�U`U��=�C ����t(����>Y�r��pU1�ݓ�4�H-On����} :zfGQF�.O�O�Z-6ܒ�*���ؚU�^���R��"x��t��	`y�Xw`�P�`�_�����w �����{#�CxW�x<x��dO�D���TZ��#���Z��(*�EN֧�=�A���a�'XNPjo$C<;b��N/E��`4��Tڛ]�b�3$�[Mr���ʇ}���2E� �]у+l�*��Rn �,���"�o�|��kj��9��!vZ(Ʊ�<�����k�n�?=�ٿ�ĨE�8�{t�]6��M��4U��I?�8?⭊;YL0<���
i�����n�u���Ӹ��%*C�Գ���C��[Y)�/��qތ`[N9�kh�kέ�儋t)��'�A�������`�F;��T��8m4�c3�v��-����	����8AZ�b���i�#��;�Ǽ<�܅��^���yI�s�ݸQm�:pt�=�W��6����{��?.#ڡ[!h!��W�>8� 
���~mѹ Yo5������c�Id"�p��A ~���&F� ����%"+���E�i[i����<,��w�E�5�ЦDi��R{�B!��r8�vXp��sv��
���o���s.{i B:�;�n��_ ��꾀�_*��੩����d��ǜPX �Sh�'�M�{",璌�AhD��P��UBN"�]7��/���X�Tr�)�
�
��g�mkDa�5����(����܏�+9q&pnjO۹��Qs]�"��1�Y�i�Њyyo>Ʈ�r�i�>E)�e1 k�C��VWZ�a<�/؟#ܹ�c53�4�nM�yMW;ܐ��I�`ᮀ~��ܜjw���[j9
S�uN�ϙmw�]j�V��.a��N�٧��hXJ��9�4���r�?P_�~�93�t�E�a�RS[��*�i�:,ϟ����\ɰh��
x�u,�ǱHϭ8�o5lv�����;�I���IM��.6e#�>��ut��z��3�Y��I�~���
=�h˯~��#�I`���z�eh�
Z[�(���;u�3�vo/��+�y�98_l� �=6[��ɱz�.O�n�(h�V�LK{�0�E�ԊP!�qV�ט�"6E���Sv����ٶ���%){��p��>|�H�d>�0��T���(,����i-Q����8Ѽ6�){�Mh�"R�}� l\*W�N�����������p��ڑݩ�ˇ��&|| �߶^�������n{L�
e������Io#z�_�C���,X{���;)"��c�g4y��?�)M���4@aRAĘ��wKt��b汸��"!(��=�~9�����鿵C��iD.����T�!{i��g�c�XK�T.x�z�
��'���͎�c�Ekbum(g���<�1�[l#�'ڌ	��?1����4-��#y�)T����X��0�+�3	�/�\�e�j [C@�J�Gft���vJM��-	��ܹ�sU�_�,X�����׉�����vg{�{u��B?�M:v�'�.���f�ʣ��?������˭�����X�P_=_���'?x,�׌��U|�נ�{����F�w��^>~��l�-�gU��>�x��sMf�Zc0������|.�6iG\4xW	��!X���Dy����-��(��E�<`6�#íc��Yw�V]ȉ�ܗ^�,�64c��Q���1�\聎�:�P�函��u�Y}&�V~pg�J"����i��P[�E1[����\�=�sFYE<�<��dԻ��b�g3�����]��tq�R�Dj� %���b���"w+_�^
ǆ�h�%����K)k$�0�A_�����F�����cܼ���AZ��}�bK,�U���T��m]}��MW�lRR��K��q�U�K �s��SR5��'�_�5�/�#�u��	��w�qU�(.����Y9�:��dk&�|R���Yw��{�$xb�(�0�ǚ���mw.DԲ��!���`�q$���s"�Cيw�]��0��֧%�5�H��.������ �fKP9F;,�wf�<���(���w���i���iPB1�lńb�`�<���JR�&^�<���[������0��ti5OP�MT?@�L��{�1�
E��U�%��1��x���Mm�he�ݏl²�w�\����W���r�2������<d��z8�miOӿ�܉�;K]�M�^X15$�zʡ�1D��B��
Y��ʓ�H���D�z��I�NR���`7�q�I����>�,��0�A�Ak5���-S��h�;�Ũ
�'Rhۑ��E���+V���,�Rsr�}���.Nl�t�˚���S((�'�1���̥�n�
��[NC���4"cq��.�7�����]_tM1�;�g}��pj�ABvIH�j٦�w*,�#�U���	����eg��:����E�#�j�n�Tg�{��-����~�����XQ�]�M��׳�ӥ��8��α�]�7{Z��c���n��r�Rx^���n����5� y��X;YX>M ,��o��K�'�f25����5D�E(\В���^L���S�ռ��H�̳�b���0�/��jvYP(۳��)�t֚�c#-Y���<a��s@�j(0 ��Dm�;,��ϗG��#���θ�xSP\�E
U	o�b��M�΄�����T�kBV��R]֘ԦK���X�#�6���=�D8{�y�0W��1���!�4��i��0�:d��y��)Bׁ9�(q9E�(l���騷�}���p�"X ����>e�q\l=M�Nq��$�L�$���^��e:���m���J P�RɅ�=?t�sR ����t�Ŝ��P��T�c<JN�W�������Ru��v ���LU�9��{�-	�-x���b��OW�ABל@>�7��b�B<��w�=�����1��Ik"�[�X���/
�%���0A4�2���'?Kz��{�ѿ��ck�W�!đw�-_��6��㫕4{"���[^_�ru?��H�o����E�%�H5U7N �0^U�z���n"����d�gȖ�0��f���y�\^JoN���S4R�*�d�P2�Z�R��%���⁩7衪iڼ�Ҵ;X�SUl��L�$	�!;G�ƍ��~�G46�u��V���S8�8�c�pO5���e�BN��*g��D�q��ذ����|����lM��[C��*-�����('|��h4��i�S*����/fO�18�&��Q�(q��f�& _����q��� ���y�7~yц%>�U�/��}ܠ;ג��&ֲ=2��e�x���
��1sb�X+�jo�.�:Y�E������*�*`N�Ǻx|��q�NZ<½9���o���� 2jH��M�*fj�M,������^�_+�;&3~A���3Jt��>�xC1�~��ǋ��e$�7�?2_�J6�kթ����=D�*T(?<���e����[H�T`���|��^qA�5�&�$�����8��t��L*��})t+~��B٫k�	�N|�rIxkG�T���3���CN	|��asá6Čm��du�}ƍ���� ]�"��W�U�����`o ����Ԉ�ye����H3��?���S�/����	3�ŀщU���;_��'��S��A �
��� ����`8#�ܓ姨��}k@{���6��t!l�K�����$���ث����{��L��_�������^6��������;B���G������1�9���^�ܺ�\�N��:���>��p9-�A�08��$8 ��$>1�dޗg�_���m�#O������L��?��,d�s<�l���'SL||-��(��g,?q)_ւ#z�b
�|;��I�� +��[�k.���[������N*��� �����0 H�ǻ܆\��eX"*�"�,��&'ЛSߧ5a��?/u9B$��Mws��
���/�	۰�nts�4C�)��,.�V iw��T��(v�&V��
�M��қR��љs?t>+�
�A��L��m��]�rSTi��`�WvZ�QR<��?�(�Q�/^>&��ad����ȍ����J4*�`*�9���W�%fZ3�U'��T��a�4]�'�����_+k�+H��r����s. a:(\5���ʕ��DHѡ�C���(��0P��W�Osڡ��i
�!�����z�!R�.8�{��q�'[?�M�\;��驕gd)1%�r����!��b�z:?�ͅ:i�ٴ#�<�!wh�@���	2Ţ�k��# �[�u����AtT[.Qt#�2�?J�X��M�G���(�G�{ڀ����O�G�}��W���w���ݢG�EL�%i��-�&Q/8�O!�ǒN¦�A��-�ǍD_��h� Q������b�������9���٭܊���|�8���	i�Xp#��� 3�C�I����aE�MF2�T��k����#l�\
��~���I�C�o�$=�-$<��:�;����3�]~c���[y���k7�����w�������F�Y���`z\v?/~"���#�5�fY	�M[F�J��%�SC�x���\�<�l����g8+�����ZNhj3Qɛ��J^n<�;>�3{����_1����N`,�8bG���������F&v��a�G�7��E�kݏ�#�!��������mjX������:T�M�DS�/ʹ�ʧ�c}�KlV;ia��'i�A}�>��j����v��N��ն�k]e��DG@�FםM��,���0vWo^�:%�w66=�K� 9�U��c�������e�b�ty塼�Sv�L�C���Q-ӂy��9Ϝo�9�蚱��r���}k�0L�cJ�Z	���U�$�-Œ}n�J�ƭ�V,A�y��?E�/5ϭ;�����l��7qabc���e_�eϯK/V����LmS��f�Q�YMNsBK��� �o��nKb�Hmg��!��L�wr��p�q!L���K�Ԑ1�l���B��q�����S%�Zܖ-�
��a�)�@̇��z�G~�Pul��V�F�����k}E��qQ���3�Y	7Q���K��EĆF��(������e����8�3̇ll�Y2�-��ol�����>]:)��6�}���5�B�~؛{ �b��q�T|���c�4��6�9^'��:�g=w"��v�x_Q��������+�9:U��ק(\��"|`C�.��d+�1���_ȔO�����X!Ֆz��0�7f���-��~~��Y��$r��'��ߎ���*)Us��݈P� ���U{�2}
�Aޢ�wG8�����:�� ��"�6�0d=��a疕��o����yd
��
BX��/�S��F�����+)������<9��ba>�ӓ��!����4��N�௡O��w�Wߺ��;UC|���@�����$�cE���Z(8lE/l���8�+�|�|�`R�S���*v����� 	b������@T2Zm T3�\2x���
9��1�4H�n�SR"�~�v����X��#�s�Wm���Jb�v@̾�}��h�*�?a��  ���Yա�{�Z~�<�̋V�w��!����>��[e��ʷ]p���f��L�d�6��B�׉J�`��O��7k�1���YZ�?�� ���T�T^~�dbCő��_�:�U���P4n��~|�%떾��=n� Ut헁�H�}૗�辡f� oG�,��0*~�+d�����d~ߞ*鯲X�+eV
茿E�$�s��{�KKh��m��]�U���t�:.��"zsC5ob��Z�!���ݰ�7h���~5�.p�)�^�wI���n|s����k+ud�$
��*n