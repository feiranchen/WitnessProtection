��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?���e�F��M#�=
i��
�l��~,�!`t[Ҁ%()�֪�Ч'����gF�ڨ��̌Xs[��'	K쏏�͑��ðƕD����FG�y���]�i~�t�W{�1,���^x�шP�L�X��ka�Lg#i�]'��r�/�rt$��)�}<���#(���#"&���6��G�0�IV��t����fC�[��2q6Y���^.b��|L�r\��,�&�?��_���~���mI������?��G�ص�K?-��|&w���Vz��Rl����p$��Ԗ�Tȍ0�/����{��Ʊ����ͼK��۽��w�y���w -�c9�h7aL��5#L�ы#VJ�K��|	����O�� �p-�����m	�{1�O��;{c�*b �p:w�]x��PD�'��������=�,i}���o�����<�o]���lC+-#><Bs!dz 3K���zA�����5�"���|��몃�xnt����I�D` {�sx��A�4�xp?�i�<�Y�[q�iE���H~���B�U `	�����x�z����pѓ�uY$27���1���*K�\Y� ����rOpͥB)i��6np�%;�9��^��|���ֳ .f��6��!H�"���N�)�����{n S%��唼�W���*0�ܛ$ٜp�χ�����x�B�͸��iښ�̝����1N���pyf[i?�`J��Q�$ֶ��w��,�A�>wAa��зky�-lp$�sZ�Kw�����JU�)��]=	�5��&I2H�j�<��#��#�D�E��P|�%z�+�xgzZ�o��T�%j���4�rj�˃�o��N��&�D!��_��8��L���j&���:r�}F~���4c.ޡ;�s$]z�Hg��3}�S�Sd�+����SP��g��p�1"��|��vF��w�Y���vŮ;��i��7�eyܜK�U�[��f ��\�t�5�zX�����5^h�ܓ����������]	W瓙o�,&m��\t���"4r��-^�_ �n������z�bА¹]��c>?��Sƍ��S���Ϟj�榐B�D��5�\�`a5�(�L PJ��W0��0�3n�~y���@�ʦ�N㘁tyB��hP����qg�7��S�M߮E�� � ʴ�Q��mìhNO�3��4��.�f�ʆ+�F.��:Λ	��K-�z -*��i&��2A��W��U���b.M��cb��2�'��G=a|�0`b� 8���YB�r4T%�\���ｉa!��o�����t���(��6�c��K��������;������t7����G�0�&͕*�*�DP��tQ�VJ$0C��g�`#�Dff��n\�_�=��Z��zo���=G�-�툱�8
�h�yu*E5��jR!A�y�=iɝ�,�2�Ȧa\��9�Y#_cnO��b��S�;Ц��^b�=��ZH|f֔]�[���ks�<��U��}���q��J6�"˚��M�^��r6W�(j1���4"E�iwp��qx���~�|G�=�N�8���Oı_��r\��^;@�����BuT���rX����-�7�c�>p�I��K�Yi��r=xE]�@����x�q��0Fw��M:���EЇ���FR�zd1��N��}�����g_t�A��~ۋ��I�u1��$�����Nաwy�����xLJr;!t�f� l��ƋS��Gp�nMV,���ۆ�\ e��Mq�a��'��]�����j�d2Ǌ3�KR��&^NV/'ؕ��jj}�C�N�
�6�fH}�4';\� dS%�r<�;0�q��J�wxӂ_3���j��������?²�UX��ʡ���� &��4���8�IU��q���`�����s>,l>Qb�JP�_���`p�/|u���L[���v�q�h�$� ����)-�(�
��.�Yh-����d� � G�UҼ�a����Ƴ�s��Io4�*ԡ	�pli�K��(⒕��	;k3I�i�ky���xBK�ӟ����_:A2�ȝX֒᭏����C��Hf�pL��R�P�	��0����h�_�O)0� E���۰��ĥ�pT'�]Lxzos���h'���|�(\;u�w������N�7�,F�No������p�=)�����y�+�.�3R���_��Rf��~�D���θ�	�{Q�B����rD�N�ɧ����tveY��[�GE3�y9�%[� M�Y�GC`��.Ǎ�b�&Ґ���2xI7�UX0:��Z0��{�zFbU������rA��T؇�cW��v��"�������U�=�^R%wF:lÈL���0է����v��#���{�2^,��	zt��g�+g��{�qM�Q��WW%?��DKy)$'WG\���@��r�X/�}����� ����Am�I�����)Lvs��/�����#щW��iCK�a��(u\����y8cԕc� ��,�E���@pM�1��d`FZ�߃�5�����R���ı����E*Au�,H����T�;5�'8]��tڲ���]g�5����[������i⛧�Ŏ��=���f��R��C;n�.�V�Y�tqU�D��m��ST�L�eR��d��<LKY>��0)Nf�C�z�Hx�T$����%�4B��>u�\&�(�c���
���1-��/��(���9�e��0y�{����j�?X�i�	�
���(�%؝/��02DtO^:ws��z۶{���a���#:B�5�z�=0�?MG��a$�MX�?�!�W��~�G0Ϛ��ӆ�7^/g�A&�;�y���M�v�6��X_��E���m�Aiϸ=��()J,���@Qyix^���h���U$��k�w̓@6J��Q2���k=N��^��0e�1�䒎z��%
-��Y�*Y�v��6υ�!s�hw�	 ���(\�X����	��**��y��]`���b10�݄7� �^�:��9sc�t���lo�cZw`S�%Н/��@��Q���Z;=+���`���e��2�ˡFs����Xe{$�jפ1��e.K��)�8��� ]p�<s"gk���%��� ��^4u�Y�(.Ա��Q�zN0=��i�r�<��B��QB�{D@+���M$��@�^= [�L�=̣��ߞf�@1�4J�3�N*M�3"zKލ��S���}�rS���̸��8ʢ��U��@JI�5�TWϫ%X|z�t���1�Ɲ	�7�v�o8�HFD���'�����q.H<9��V��w=��0����;C���S1ߎ��h�1b"htƭ*B��47����r*T�� rzꩊ=W�N����)�d��؊Ǿ���e���ݐ���NKv��ubaҡ��0�ԫuYC7�e��*D��>�Q�1�������0_[;*�y!iW�0��(���}�6Q���<t��j�|�z
#�AlD���-E�����3�.x���2��|�d�� ���&9�qNjNm�.P.��TS'����Z���fTLÄ ͂<���P9�����E�UoV�ǝ�4?�<ɻ`[�1�)hnc;Z?MQY����U��vs�ʷ>�$*�y]��n�C+�t��V�m����5�f3�l�`�`B+�t�������+�C����Q{ٞ�Oqn "	w��ځֻo�]�d�	ϳ�g{���7j��!n�c��ɖ,b�G�{-�*�:O/���J�`�����ye��C-����v����mմ�|���)���X��D9�52�ڸo��ޛ�����}�.�4h�P�n�#I�-P���92'f�BOiѨ�N���+�hB|��0'�	�vb8����f�䓆��{�;�~T����U�M�4bMh�&�TПJ>��S�N\(KT?��e��z���U�����u�^�!;��&�W�n9y�sz�&�|��<�QY�mo<��JQ�D�6!�+^�OT�gg�h�uY~�������*Ȍ�_} �ࢼv�����%�A��D���8"���잮�D�&����.����H�_"a>&�\�^�;m�m|�@0����@fdy�"?ʦRA����{"؆�L~�Z`�c�ITܢ����[��c`�g�峋KWW�M���L[��5���1GPs���=�T��1%m0@���)t7g�I��+I��X�&�E�S2i��u�1�����.�Vg�)s���4��Y��G�����N�pQ�bv?
HJ���cD1�>J��3������4H�̥+��D�| O�QQ��M��T[��4�ޅ�|��R0d�T�+h��������2����Ӎ���Q;^� �@�3=����d7kT��(������,�2���8w�׹^}Gg$�r��˴��XSŎG���w"�"P8�|���[�i a�Vhй�`��E��և�[�P�o{0l��~�c�M�*�#ѭ
i 
�bt���[W�Jt�9��)�(���8h#e�N:���5ߑ �_ ����i�׊w���������ex=K�����x�y]t2���S�%��)\��T?Le���<E�''Z>=�^����ƛ{U��KW��j,òD�՝���y��y�Gs�X���Q���d��I��{�+�i\S�E�|�V�$�*��V���`��V�5q��P�x����ݲ��>��5Ւ���'$5p�j��U3�`	�c��!�5��@ا���ŚL���uP�-����LX��B�I/�I38���4+�?�N'lJ�n�������w)��"�q���K�I$Ōf����Z��1B�T�FB7!ު��?��{���o�w�l9J%�Dӊ��$>��k�/g�g
��p3fmK�j�xDԭY�2�w�#S7��(e�L����-.%�<��D�GS&<%�|Ç !�O#�f��(��O�.l�o��l!�eG�:i�5�,*��������3����1�:���7�xi3��g�"�J�`��
4�(P���j�SUx�>ص�=� A����X�8vY�[qŤ�-Xd���~8��<��3cv!�k��Z�K�b"Ն����ͪu�����!��T��eL������5�4}1]?{�}G#�#��@�p���̂>#$!��_fkR�`Fk4�0���\˥/X7ߑ5�A����i	"{6KB�`��k�q����Y;�=1��WL�����A4�ks/��6����\�HHK�7j�o=�(3�����0m�HcO��ʶg`Fi��ﵓN�d��K�ak�~� ��7��(�(oN��(���P<y�hq�f�E�Nu`���T�P�=%�P�6A�����<���cL-�����A�����0�LM�0v]�[BG���jN%<d�_8��c_Oz}+��[�~�|���#�r�"�$m�}��6�����p	mN���癢?�XL�}���z��	}����<(KXf�4 pT.�r��mk����
?}%��B-t&��|�ZF��Rt�5Ơ��i���V%����{~^h[��&l��$-��/<dh,3D(���+x@t���t�z��L��om!���/y=!��8{�響6ʂ�yH�5�ik5׮��&��Ot[ǸC��]85[������� �`��Y��|�.D�.�h�'�P�6twb�[�����V�����EF�}���x��.���d8w|�=���<88��˛�~G�&��8�V����b+�@�F�	��[�]��J���
�k2 �g�J4� �<�ꞟ����/Ll�I �>��z��
�=��O� PoI�ok�g�C�]��'�-T_�^I��f���W���2r�p��k H��W�66����iM�s�ndpzQ��A���!� �\Y�5JT�o��'~#f��{�'X���|�8�����q��#v�����T>nI*���*xH>��r*��V������VN�y�1����]�]D�ov�^��B���Z�=6�X��f�r��k�C5��}Kr*X*��7�zϡY�u&��Qc����O�z�_�ev~��H-��� �(�P����]�f:�K׻��4��{X�C�w�i�˔7^>��`ٗkA�Ұ��H#ߑ��p�5jTz�Pi-&���ʢ7|����P�UR�S��1Kc��J�����9�-(�E�cֺR��X�2��2�½tm��w���[�
{6�r�Y���RՌ(�;�m�Mv4{cgY���og(�n���T��"�Ƿ��)�8
����TR��������
��,����-�S�+ʜ$Jw]�*4)��x�="&
4�>����q^� ꒽��Or����;dp;:H���"������r����B���6;����b��8�+��p�A7�C��/�ϩ�N#n��g��@7D��2OP?���	HUXO�jU
W}tc?�N)�{�����z��;q��6Bt�ρ1i��d+����B�{���V�a�$R%i�ٽ T�K��
�}�_�B�a�J�,�>� 0ogM�GY��:�;���L�K���Pz���2YzL+?�J�)ڄ{�Hu��L��l�h[ǧ�h{�IX79�w)�H)��?z�&?�&�@�Cp�hk%v�`�+��g�-oBCnLO�&J�۫�e$�U����tr�7&z1�47�D���K���<�����;���^���WPJ��r�7O v�K�����^b��w+�_;�j�NC�����$ZL��sj����3�����8k���u���ŧ�~I���*�>���hrcL?fϒa��z~��i�i$Q{�\�-S�6_�m�@p()1f�����T�ͺ)C��{�UC��/�v��I����`5[��m˫.]9��󏊳^��Ð���,̲���������0�`�}�Bg�Y��/Y�P�h�K����L�K�yR	����2:)��{�y@3(���?|���]}�x�c�oXjF���� ��"Q;�*�O�1\@Zt�j���q�WBS2�	4��i$�_�0���x�;P�	I�����eśL�|�|}*3P�G�Z��S�q��qhzGVCP~3)T')�"Fs���u{R����A�ى���uga~X^B�(A��룿򓂇�)ZqJ�8��"F�7�A�1C�e�,T�/{8���Če1�q���#"���s5�<A���ٵw�k�``}�RY��0�yј��䵉F K0��7s=�xA�-rV��QC��y���K}d�d���W�`
��C�v�/��g�d����ϧ �L|��_h\��Nz2rF�ߒ�\=�K�پ��>�BT�{t��)�ö�(�a1(+3&���Ə����t�%R�X����x��/��Sg�L꽹���w��eTo8��pR8߈UjO�K~���{�tYNʺ:[,�Q��{�����GpQ��8N����(�j^��%��ƍ�k��w�(|�E��[9��/y+cֵA�����3vTx��(�Y����]tU�zo��L�(�7�sMH|�p$�l涍f^��{9��HÔ��0��]�U�$U+]�G�`������n�C�Z�#M�==���]88qZ�2"�ú4i��>�T��m��V�Y��ň�Ke׏�E�GlD�C��6Z����h�Aa��K��>�}X߲���.F��Z����C�m���5z<í�͘<Q����WPG��J;����5�����Z��F*�E��WB��`�΃���;�[ׅ��'kS�"��W��&��o�O�]!ق'oF�ͦ�P�[�v�\uG:iO��!�`�1�\���kwo�J�2�v��1*zӰ1Z�б2��|�ќ7T�
��;��k�h)�"�o\��<3&+F��g�^�=��;A=6k�v����@�Ix4P8S�̪V�6�M�bw��d��z�)�z�8��F��&�m��H^�y;[ا:��/�D�	���Ʌ|s���mų���_�B�ճc
�%����	If]���_)�t��9㕇Q�b�c4�dyV��@����A��Z��E���i?M��ɏڒs��{ƆJ�L�ږ�m��2��$M˗  ��XoH�^��	������H����|�K�+�����y�GG���g����o{��� �{;�kY��j����@}�/�1p	6��Q�snr�mkچ�6{�Ŏu��е8,!�ʝ��[Z�az��h�]��b��>��:x��W-�000�ލ��*�|�h�a�,��#8AW���Bq�u�L�4�U��Wǳ���� �=w�in;� ��6��/���
B��0�I�꿯�IS��nU�QR��⑵6���+�# wy��ͺ�{L�}� ����m�r��H��n�͔%��@P;�����~�l�1�X4@�#�kq3,ϋ��;X�G=-�k<@�zx��L�"����!���	�G��4u��D�ʰ�,�gC�`:�u<�D2�(�B�+���A/n��	 "��Y���PT��xN�YsD�Mǘ_ʣE�Eg�S��W�&�����a�e��턗--&u�Q�Tj%,�b�ѹ�;���=�3��*�S��%�ăZ9R��fbT6�>��t��|�������^"(e��P%�7{�ۆTNF&r��Ůb�{Xp_�̓ޫ9����k�@������]��֪wh.�I��
�so�ޙb</����(���W���D��{h3V�t�"TB�D�m!
�L�	[&��cS=S[TB� �� �a\M�_�}0II�/��I�M�ݟ��h*���O�ي���M��[���kC���V���]�F�?�F��u�y��=�w�	{�[j��iG��/1�-��}}5�ft��+=|���k��K���X��82T��^HAn�e�.Űfy'$�>P����1��������	�LW����
�<�� 
�:���EZw��p�X��0qT�HdO����g�J�p8�ůJ>�E"��h�X��ez�k&R���i��3E7�=��'ڽ����6�H�Z�Tk
���Z��m�_ʁ"t�|j!��q:��Ўv�3\=��£�}�B��g
e�kHH=�_R��ю ��4�ZrսI��ř���z�`��}�x���eX�6�¿�����TFf�F��?OK���'�uA]|Wr.qbq�np�~��úr���=�FV�=��X��E�,[F�ٵ��&k3���<�����h�H�z��*
����-^z�T{����^j7C��x��p���'/�˰�Q�2�o����Z$�������u�����ULQw#�-���'�*�D�9ٟT@PEI����_�磌�5p�����7���̀�/��Z�7����>1��`�yu̦{�8�x0n	�k<�_i��S�*,5�%��KA�[(�!�t�5�$��a��_�<��kB�Mf���'ڧu�O�E�iS1��������`��yde��۷��B��h�DDf�҃G� �w��q�߮�wHZ0�_�����@�?�3@�3�Keu���N�e��	6̠Kw������p%�
O���H��f,�*4��ƽf�bXɩ2i�4C=Լ��5��g�P'���V�]�|��@�:�`K�����!�-�zw �9^CZ��R���R�a����A�c�՝t���o�{͛�D�SF�����F�J/������OK���ί�T�`6��ʼ�,���|>G�6;�~�7�M"F������2�̣}埪>hv�1���H���KA4�/�j�$[�ʞ#��CRt�٢��X�$������.����*��>[��'*n=)ͺq�&�㛡����l@:�fV�<5�NU5�#��S��TV��s�0��3O2�f�����%�xi�;�4_�P+�+����ob��/�e����uZEx�t���'���8�;�Nj����Gt�8����}�ͬ�Q,� �%)�b�ezjzx�y��5�h5�8SV�Tx��o.����4BS����j;��B���~b�~�e�����r;yC����G�8Ko0p�nW�
{aBmBB�5	cX�A*˫&����JBۑ6'(=$�&HF�$6���d�Qtԁ�m�Q���&��Z��N�Rv2ur *���'�&�uB3a�ET�Pߡ�Ŧk#�qe]�v��W��ENqx#�m��r��j�k�Z�㚟��N���O�ҿUj�;��9e*&�5:�1Y�M���c.��sXG�c� )s^�t{?l���T<����,��v|�=��f�m��
���=!r��y�;�M��;�|q�0y�M&��D�����[�T�z���+&
�K*4���&�.�a<F� ��{������Ȫq/Ւ����&XN�.aڃ�E�������P$���i�f!�:�S�h��y��Cups��8l�E��(5������+��^:/���tj�n�v�ۓ $
�?S;��T��C�/��,א|4O7�(.���!_�p\j�X�9:x躴�-̅ovr��7����؈I;�eƕ�u~x��4]�3�b.���,��LS+�-����s䃦7~%�ek�.������.��nnC�j.5�k!-�cl�x��l3���L�o Ș�F�U�#��ͧ�lD�#ܿ���i����QiO���G~�-bت��S/Op��tY�g�R	ť5�}����oCɼ��|��F�q1P��&=�E��wul�ES�7��dyk�A�D������6��m^ �S�9�t�����m�L�b��Y��;��+{���Ȟ'�R��3L&�#&���3���:y��Ј�m�$ĳ�DLڢ�����L�#53yb^}��@[��&�&��|��s���:D`&��FU;�&�ҕ�d�)\���M�b�
���9��4V_��$�&���2!��>�ф]ݶ�4d��hhv�vq��d����"��rd��	t�>�B�>�~A�|�#
Or	��8��+=w��=�٦^�HE3��C=6�R����U9�6:�hyJ�`c�3N*�`J���TD��w��u�I��E�V��t@D|�3S)w������_�/�4��Oߤ��L%o8�l�Q���'�~���(M�}����0đ�Ri�D��:�d���]���ɪ�sjy�?6{�
�Rx7�",��U;Ek���u�o��V������p7��&�d*䪟�í�=(n=E�[Q#�~�W>�M
;��F�F��),#e2�Ϟp� 5n�����]r�M�\�t����P��n�VF7xJ8M���]��n[RǬ�2}��|���������iۉ0 gc���J�:i����Y(�.d�m�;3�]���	
j�[���RHJx�=`3�+�P�OKJ�*#���ƹu��!�f�"/���aVi����u�p��h���.f�9��
��U/H�/K�ٽ2��s��1�4m�j�x�h?�Bď�35�U�ט��:m���bi��x��pͲ��d�g=*�j�_�	V8��������j�z��ժJ��h�p����z��O�7` �iDS-dFP���j�g>�����+�'Wy�]gv�Q:p�	��E�R����5���d�as��dC3���C���G��Hߋb�w�W����iZ�L�}pQ��,�_��?|g���5��V?w�Zl����[�h��NY��b/���NMn�E]%"�����+8���y��gK�t�����)M���?�(�i8�م��	���0f��(upz���	��V�hM�,r�7�H��?�(��j҄3�����YܑFOE ��ꁽ�$�U�!�"-~V�[
�	���/�|Ц7-��$;zš�i��l	K+XZ\\�J�o���sJ�'f��!Yh!�c��5JF�7 ��ǝ�ٶX�*��+���5��|��)���A �0��T菳M�!X���/q�H;�@-ۙ�Ҕ{>��%�7l�)��[�T��h�u�tz$&�����πp�d}d���+�4�c2bf��N�p�v�\����0��[�ki_g1�i�Qɻl��L�XO|4O�Udo�od̦���'/D�}kP	|�w��Gt���M4��-	3�5fbI}�[h�'��r�ћ�j	ic:$��`��j�ܻ���NUY��A*��l�\��p}����l�>�y$���7��JȖ�ª��t>�}l�$���N��[��2������� }Q�C����|��a(C#SY��6����e��gTC������2
.�݀�Zj�z�K��x�&!�򀓑"��K^�w�jO������R�OB$B	B���-�,qJ��A���8��j�L��E*WI�J�#yD���PH�>zd��r�R��T�)��#*�Q�U��än��^�L����N�C��S�k��k��cu����������`Q�S�O�=�X>ZAԲ�U�+.�;U�"��3��-�^1T"
�/�+�G��ف�7��/�S3�Cre�6��\�Xj�p5��Z]�ۨr?��䤿eWr�ƍ���J	���VWo&��0=ܸ��&\�)Qf�sgGvڨh���)�eγ�)�
��2/Y7��b#j�8v������}��ؙ��W1j��aˠ5��@�f��!'��nw�� �~'�=*�}}]s���Nc���u�|B�i9$1�2�e��Ԭ�4H�k���ɓ�(P��;�,���٣�J�� �x$��{�	x��F��V9�Ne%��`���W�8Fy�_��I�s�R"��ЉP�`�� �@ E��*�1ٙcǷ0��1�*�a�����]��,�L�m(r��g�D��w��X�bm<����"A���+22���z	V�4��z\���B���GL��K�9�k-'��s��NMG�xf�''�c�(�čzD];X�1�w�B�އ�MPk{ćp��+qEl\/���c�]��+oKH2;I�3|��T$���CV��F���ܯ�:��4����w��w�?��n'g�g��6�"�D#��֜C��j�%͜f��u�=�Ι&�����~����7v��A���F~�ZEU��D��w`(�C�M�Yg^���m��Y�,�;7��Yв�)H�^���N���\wU��A0h3�vss
�}��Ň��Ѐ���[慧��R��
4z3�=}�핾������_�]a$�w��ΐe����r��$A�928"�Q�̥_�+�\ ����O9٫\�:Z?�\G���쬇>��'�l:��o��2Lo_��oC����q~�'��04� g�ëъ��+>�Jh��vBh�IZ�*�_u�H�g>��ۑ�_w�.V����9�"S_f��܀^��`���1*w��{�ά��o �Q�����S��I��l�����aģ^�%:��f�9�(��o|�&�x���I峊F̂c6��C3z�g7��f�~��%�o��9��@Ӟv�թz�V��#o��OS�yQ)wB�E��B�8J*	:-]�A�7#���t�Q�pӁ�N]�d����9�f�ꚨ�	S��d,�%�o�R�ƚܱ�,V�k�kЎQF�hno������꿊])����/�+�ׯNK��9�G�B_pkX|Q�ȧ ��x�Z����M1���73�:�k�P���=>%ǂ�]
K�3=(� ��M���+��ODOJR�0�lAf<jP~}��@|��E)��b�ޜ�t����FH2m��A��t�u�Cy��������|���Zc�:������
8S
������M���u��ɡ��[��VI.;�=v�E�w6���jZ��Q�p��ֲ苈�S�O�G��>�F(��ov��9/��j�js�_º�y���~��������xW<TS
��W���0�`�ÆV����/����%�V�IC�>׬��,��6��$��µU��*�c+w��� ����b��_m_�����K�8��6P�¶n���:!����<M�2{o%����eK-�e�R ��y��A��"e$��d��L�}H�F������y�E�l.�_����:e��:�����mu6�J4U�v�F�ke>c�k�,�8�Y�U�GQ}�)؞��}���m��_C�9��ղ�v��X�6���%��>�h���ܩղ�B��W������C�~�*]�,�����V�F;�k	�����	�B�ӭ�?��9�q��-¤x˄D���iv_L�E2�ui�T�3r�ht$�Q�+ys�ØK�̑�����}���� ��o��P'�;�����k[X��32�4<�/)Evd�I�Άh@�f�*$ O ���l6`j�f���d�[}&�
����s*���N��Ru��l#(��ҷu7bm5�=Һ샱��%W~��f�O��;�Yz�b�uj�Nb�	�B�4E�ʕ���+��m��h*�]1���)L}�yrJ�sn�Q�cVYV1S���=z�r�֠�m�L�i�"n����!B�]'��2��>��B�[,��J���ci�+b�z���n-}�n����g9�e>�ת�P�av�ᤤ}�EK�#�����-7�FI�~L�8�6ƻ����lE����O�SD�!�Dd~M���Z�V��/���J�!Q~߈fK%,/8�>�G�{~}�d`��տk�7�"�">;M�x�`�$�*����8�5�$����$�I�_�X�dN!w�3T�1��k�xF�?�(n�Uh[��(�T�Y�s�o�%�	�`����zf�pJ�7�	�p������9���o��|Ѣ���,|M��b�@XW 9k��h�v��2����U�L��a���a&a��9h(��r
��0mgj�E*�I(P�# �Q�<���Y�����h+X��I!S�"�3`� ��:�������7���I�"�Pټ5�Hɓ�A�P_8����0=a�L���X_�?�8�v��`�r��2K�� @y���*3;f�@�/��NV@�^������[n�i�'�Wa�Z008� �(�O���o,���-��(޴}m���l}9�W��N�`y��|PreU����{n�m*��?�9���[+�3��S���_4"8/q����T���7N(�͍"�j0Mk篎����_��%
����*��Qm6
l-��Z5C2�h�t�l�h���q�D��rvj�x"@ˀ�� [n�G-K9�em�8��ly#bY��j�*�S��J��U�)���?0�$�+�v�������^�� L�
�!j���%r��6[Z���-�w��aS���ex��:S|�{�N�q��9_�{9�$��6��X��p*�cR�O�B�}�������NO��w-��m��Z�S�4ϴV���-օk42û\-��cI7fV���)�]�9C�5x�WO�5لY�X���(��F����U���b�N�zÃ�|���UXV#��ͤ�L?��-Ӛs4}b��:(��;C����v��/��mh���p (2����f������5ˋh�&��fV�1Tx�;`3�/��,^)W��?��Q�y�]ǆK]҉X"�3٢�:����r�Y��X͊J,+pd��ğT�)*g�:��6��,����JQB��������l6��F�8��o�Sr�$J|J�`�E��LVQ8�W�Q���z�����`���\�����#�������
DAp&{y} e-�&��`.r��_��!�Ҋ�����;/��e��)�b���M{�E,�H���嫲�c��\����`^�ÍY�{�����Q��d�.4dɧ8����׼�Qڠi�U����H��3�
�\�a&�J���!��ÆLM(���S+��Ɲ~O92u�F�s(������y��.���<���G�ڝ��Z�#֢c��ڂf�����@ްU��m����Ktg�I�����\s[����+n���S�wDTz�Z��@Z���I��f �"���H���U-����b�Cx2<mK*.��P�����د/;$�Wb~�:㇔\\��#��F��	ŜQ'��f������b�o�_.36�7��v
��</�WP>��g|�U⥓�rXL���U�O
�<m5��$3z��$�&�Ck�����p�uu�)	��	��H�~2�*�K�T��M���hK��<��.�����	ʯq�t;��R�
�X���lf�k�8��T�"e��vY6zqk^.��������r��kׇV3Jy����b}��ϧ�W3:�s]2.�aa��',e(J|�F���K�A2�v2>�W4�R
D�׳G���oh�q��D�j��,�@
;�t�Kע��@B�Wc�<2͖-���4�D�p�b��$��EY���יƸc�M�t;�M��mY����Hv]����3�7�g�!?�$�l�|��&yZ������t͞h��������-�M�'��j)|�c;��V���Q�^����4ʼ�>/���+�\~��� tb��!|�aq�X4�=]�D��"�s�j=��׈����Fe�٭w�KlT����g2�����7���ܜ^m���'�m�Mimo���Q��H,�92$�J�i<ṝo��[��A,��L��3F^�=[Ӡ������$`o�f�;�|S,�,�,��\p��uӛ(m�Z��js\X�G�:�UC�?I�l҉
���5��#@��g��6�\Y�i��HE���W��5��Ф�P��SD��me-�pk7X�O��6��3���Ҏ����;�� ��r3�1�B�� :��;o�,�%����q^�@��ʕ���]ev�MҚr�?�?��s��wR&�N�܌���ڢ���檈:U��ɹ-\�d5Í~F@R����{B�8�,��G�ܜ�^D���X��-����M/6���j��V*E�kU�7�&�B�z��x�+�?��2f����.���9���� �j��/�`{CI1;g5P%�h�5X3�-6mq��oƋ�}>.���)ߴ
?�!V���7#-(Oj�O��?�/9$Q�A�&<[��J�iI�<�;��WR�aɡw�M�N�cS��<z*��1�Z�Dd�26Xi�j�8�S�ܟ6�"��ѡ��K�z�s1�O�$����9{��;� ��Ŕ �_؅N���Mz���ع�;��~�pq�� ���"�s"�r����Q5nc������"���*Se^�ÿ������ ��)��֥�%#�<���5�c�(7m�u�3�m�v�Q�[>0��|h�ϥ�=�>������~��@��z8m���̈́��v��Vnު��X�Q�O�}��΢��v0��HIz������̏����!�y����ّ��=���P��q�+8��i�NC�_���m��2�"���H������ֵR������'�"������L<�Z��4�Z�ǖlnP�j��
����L��$d�8�ı9�ˌ�9v����`d��k �g��1#�TH*�9%��N��b��/s�@��D��h�B���<�-L`�k�{:xL?���#�3�6��F�[��B�r���h �2@�a.&=���8|2��3�P6B懷�	z�,u.�-f�mO�7��lM$����en���0��W5C��$���A+�d���GC�;U�c;�P����ʣ9��5���Q5�S�Ep� �6���юpY���Z��m��y*�ꗶߘ�����4裭��XBDe�K
�~uI�Y/ �Y
AH^��p~~���6���:��SQ��}���wY�u��;�&�S��A��\��e�Ҝn��Λ���V�A��L>o��aH���"�1�A1l�� ��U�7p[�6���f[��}�f�WK�x3��Gi.8��������hwށ����$D�CuԼn|�F'bm�N�}|���UZ�B���m1�[��~t����~�˱*9ؓ�ps�>�Q�6:�R�V����PM��I�ܬF_4�RKw�~�7�S㓃�2���(�	�&3�]�#�k�Oc7�)���C���T�UVNɔ�t@�� �Vo��'�|¹ھܯ_Ư��UIbw��94q�w���+����1�^ݺ`�S7��HD2q�&��:Qǂ ��|����4�7��u�B[��}� %M�3�W/��lEɬc��ީTE���zsg��j�-`�%t����Β�IAQH�v��,l��	�ʳ��d9Zv�{�7����ZL���#�����ee\ْ<K/�m�#���W?��(��}_K΂�OX����E��U3�Q%40SiA2� �0�񴤥��^r8�`�H�����e/�Z����K ~ݓ���{;�8�T�{��GFAǘ����H�� {�( с��4�*昙'�*�3u�`�.�n8:+��������/���k�"�b����ӰU>������M����ǖ�-?p��{����Z��i,���Il��#��(�T�t8�4��U�Xn'.�����	h�?�7q�嫋\�m
���]�k tA[ݢ!0yO��]r{H6K��\�1��f���S��fo Ar��1V(
���_����Lhw�hm�ot>��3�Cl5M�d��(�������7}	���/�ÕY���J���������=8��,[��J��9/G�־R�S���]�TI���T(��i��Uh��/�s#1�yS2��d�#a��ba�r��	�Wͯ�p�P���B^�5k���ge��Wj$D���$r�c"w/�}��s��n�""�]~���A��1��	@���#��U�|n�Vcx8DbjCw%��;|��ʊ9*��<(tp���+9����di'ͺW�r��N(o�x�_��`8�e�������#D�V�C�ۈ��X��&Pd�Z�Y��ߒ�L��ǋ����yæs܋{�,Ճ_�&9�D6�lBS�P@9bhb�?���nf2�x��24~���ȣ��L��)ѳ.�e��s���ňK����eZ}��A
���6�gC�W�+@�Ĕ�d�k>�XV:�z�U>]���jiv1�*z�)<G0JK����t�KB���#Ul���`�����N�<~\WHQ oF|D�!�/�R3V�h@�}x�9�+O�u-9Ž�' �������E9��q��q�v�g���E,�_�5�5��.	��}���[YU�&�?&�1��5H�$���)�"�=���:.�!I��HPy�N(��
� ئ�$��R��A�����5��^��i*��o�z�B�p^e`m����"�ܔB���g��#Ǝ�ZBt�K�*l����;����N�yb=ϐ��>�a8T�8h��D ���@/@�W8�ݐ�X�t��R'�a��X�u��tnz��ed�hx[~ݷI3��Er��pD����.$p�S��J���z��&�zY_�K��V���;�-��=�.�N�![v�Z�����h�c��Y��-)�Ժ�\���(X��G�N�{x@�_yV����,5��Cz�;���x��w�*��&�!Q���6���V���!x�nlſ̨>�Egb�O��Ol����ϽԳP,j��B�TR��|Ǘ����]��[At��=3QxuX�z�G_�4'@��Wo?�Ǣ��G����:�#�����{�h�@���k �[<),#�����G@	�V����a�#))vO�I�̉}���g>v�:4��>8���˺
\'��u���d��?`*�ڣrAS
��M°�,5eed��9�\v��;	S�/���v{������8�aH�@;3�	i+�W�f��Oqr9��$�h�V��AO�1ȵwL� 
p�>����X��cn��2�����w?�:�+�qp�E�D��z�Kl��8�9k� 	&[B��ü��?�x�����w�p�>)c����?����tN�1$�p�w�=��������[�I�$q�6�5�ˁge�n���� m��KsQ!��>#D`^Ix��{ͮ�g�]ܾ�v/8^�R]1E��E-U��`1J�~����^WB3�{��f�T�Yi�S`�n����������ڂ�����A<��1Pc�y^Z�Ք0��TB蟤"�[�t�dMVb��'P$hKa�~ї�r�}��,ACL:Կ�za�&�b�%�tl�~�z����0��tP�z��@�.��7\k��#,�1���/�Ukv��=�~+HD}?�]�{@�`�Z�����4����$�	��њ
��XO�_i���8S���)9��g��C�֏]���z�J���"J��q����˙L�Q)�%�A��E��u.N��:^݁FvI������6��h$O/4��ͷ��lo,��FW-���� ��� �� *E�
��l���*lT�x�⎺� �b/��NZmA�\f���}��9�rĚl4��b��R$'c��Cu��ɂb�P�[|1��7*�{s]�G�!O����?q[c�R�&�{�=�O��ĎI����2���+Q���M��jy� �����>�SS�� @�Ba�s�^DD�>y%�a~��T�f�VLp���S��{Y���mSD�{���"��z�0���3��/�g�~4��X�ԃ�ry�y`y@/^�'x�WD_�XM��3��×`�gv%��\��}��������-��S�}6a�<�Fi������x���/���i�X%��(�C�U�_���b')
��[T�A	�	�1�h�6����E�zt�\�Q}q���s�p�0�ʀ4#�cM"0�0G���@x��&cФ��F1+A-.�^9�_\���Xr;6�=���uP}�8�H����v��u���1�o'.C��)L��0T�|
o�נ�u=s�V8JC��W_u\�o����!Zn%`À{�L]dJ:]�<D�s �À��$2Z9�OV�#x��mA�+�Z�ָ�����*Wz��������?���G�P�Z���Ƌ�xm%s�q��ʟ��U~t>����Z*�8���JD~}�4�_�	h�)1+�J�-5ᾑ#�$�ǜ��ب��VU/�g�D�y~�7	��T{�H���$��a��\��#�ţSvrP��*�ݙ��6�jT�8�/��lﭛ�Y�;DrHW9�x�%�I�A�Xaגz�?C�*` q���q��匍u#���@:�y��]n���~�&hJG�р4*�pR���HzmQZu��]@)��!��:a��L�lq#�i�w����(��~)]�tp�tn�1��Ka:����Ib�6��G��W��mf������E�>����H�&
��F���Y �F�F���$?R��^����'̹�w�D��=���ug�{�nS���,�v�Z�v����'�Mlp���!�]g��U���"u�q��|���v��:yA�5��]���Y������ˎ`YG?��£��1̻b�l�9�Jv�@�z�r�4甞^I����:��M�Sd��`�. �.Ҹ�� �m�>��fM�`�������d�q'��$3('��*��W�Y���(y���>�����S��u?����C�w��`��dA^q�
��K�=�h���<����H��^*�L��M?E��C���2�w������V�bd_�-�;�~b��W�x>�P�?�a|��?_m�¥���Q��2&�)�R���[`��/��ab{/"�8F���U~���>�g�&��Q�=L�P�S�r�����(C.��1�7Q݆�ڦ%E+ۨ�0:�S�ot��c�"q8� ���=��
&Ul����&۷	^�a�0��ڂյ�?&����E�|yW}eJ�7)�I՜�c�f߲��p>3�`�ew~�q<,�]����(!����)����,���h�/?
k��A��q�y�q���]+��^��B?���!��a��7���"l��j��U||��� b��k^�3�L�!rf���18{��8�B��[N���>�-1�泼fQ��T��o&#�>��\fv+T��s�iu�<�sZ^[�윥�#�S��}�}{pt�Q��ѩ��M<�O&;1A:R���$sʦC�/�՝J�����b��I��8c��K�`�M��38��l��6y�5����εՆٹ��St'n��$���.<��^���̶@gˤX�G�1��?w��Xm������J|�ۗ�28eV�~��[��C��-=^�%45���u�`39x"D7�Ul</"`�aX�Jh�~]�O��l�=��T�0rq˝L��]b��S��QՐ��U�&*��	4�5
��|�;���U�!�:<�X��_#�fj�~�Q|`X�@�&�3�	܍��% {)h��H|]����'�v��Y�q��Ɠ��������0v����%����� oO��H�Lb��}����/r[�^�KH5�Ԁ���3�FL��/���X"m�0�����+�Y�7#k"E�ps�s���
e�]:ET�b�CYS2LC+���2�<b�v)�NWv���g����EN{���1�JnAګy�e��PU�@:���b��"�0�"�^�|n�y��t������u��.�)? �@��j������ezpP4~Y1�zc���ݞP/�Ћ6�.�3���S( ��YP���<\��e_�3�̿Y�U�@;\�g��/E@����o�l��N��K�2�ɣ�k��RL�n6���1v<��E��N���H���P�uSg-9��D��� ˤ��x:V��k��î۩�!�#�k�/��ZrU5W��1��V����j�d:�C�i{/t�@�$+ �p�@�u�	M�,��b���HtE�ZR�C|I�^>~�S�U�����@F�:��^�^�7����8 ~�$Շ>�k"�9���,!�)��Ɵ�r_h�_2\@�����Z�m.ثV�A�'��J�擶�����KnS"��jr��iC��� �x�~.�GQ�B}�z3>E�;Ӗ��j.�Ţ[����O:A�|PY�"��^ߓ���&ǟq��a�����_��|,�r!LWU�@g�?:�����I2:�?�*�M�E?������^������yNj R�첋����D#֧l��YW2-�~�!�RK�9����Ĝ��i�FǾw)�-�81s�_�����B�X����{�a �,4�Aj�h�ʃ7Tj�C�A7�OO�(��:���&��tw�f({w�dx�3&5��}��0(�Xu�&7x�WK���1�Hi�6���#�CX���L�8��/��T<����~^�T�l}��o'h0q��$��[�7� ��լ 꺉kn��L&��LV�
p�`;��"�Y�!+$d*м����f$:n>㟁�-^ހ*Ο��ΩI:��&�nV�9ɞ,�x�m��U��ם��O��!!U����w�ʳn�z����e��q&�Å���XP��/�_���_���r~<���5��R�_b��>C�����Us�fA\_��l�6������2(�R�!#"�.Vdo�=U	Ơ����զ��WP��|nEPy-7dh��]ʬ ���C�BO_9Tc�G̋��*@wmg�c�_Y����@��J�P���k�K�D�Uǔe�@
�u�;�4hji���(?&�)X�x�GTR�
֜�O})��N� k�nJ޷No�W7j�����*��9s���;3
&�2Oq��j��s�g��*��)ś{B������ս�鶧��z�������P��Q��G��jtӿ�a/գ	��'��� �`6������9[ex5�E���I�=l�i�و4�~a�A�!"|��������!��|�sh��~xxr�D�ޓgP
�Zk\99�