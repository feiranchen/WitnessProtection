��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�hd�f�B���o�y�;�>Π�B~!J��/����n�C:��t���6�l�������I�����[���T6[������G�!p�冭;C����(7.�/~9ی��U��~t�-����d2Ebꪊ���I��`�oǄ�A��*|�>��Jl��q��7��ݭE�p�B�w��v�ƯY��Դ��l���gl��D�t��S�ʱ��@s:۹��t�`4�0��E��G�j�n�<d^�G��Ҵ��I+��zk���\}�#O��Ho�}'����(�k��-u���HV��寲�6��Ƒޜ��z3ڲoH��0`|����
�D�N�,��r�De��"ء�Ul�M �3�S��s�V%P��~J���))D������n��<�Y��&�[�~�Z[���4�X��Ũ��!������� 9�<���Xo�?���t2��.޾�_�����*�^r`���%Ǵ1�=k�RPG�?����j�ʰ��ʢbT
N��}���і_����س��=f���0f��x7��}����f����MR&*ҍ�K�,�&n��(���W�4x�&�У}��L���च���+�5�y�ͦ ����R\���|�Xφ3��+(�J獒������6L1&�Z�C�Q���{����W�C�Kg�P��#�	���.���p�_�7ÎsV��Y��'�+a�C�mV�o!{��q��4x��cĲ�x"+�[�{�yUP�Id��p�5'�ci���Jx�:�n2��KQ������"��p���G��yŝM�/�X��9fV���$m0����a��̂4T%���#��y�i	��(�W�Q�Xɕmw0����o�����~�@ ��Ȝͤ�1����RX7UJ���Ι��:��P���B	����x����#6!#Y: ��ytS�~����a�ke(ʓ"��]����}?rIv��e.��8S�����>#1�ذ�
���[�'P��Q
6!��:-��o��.5�| ���Ź�#�?�*Ơ_2����==�����6����}��l7��i�&�d��YqԔ�0�ȵ��_G���t���TZ>�6�*H+�j�T]Nrl�T�\��|UQq����{-�]�
�8Q(�߸�+�fK���C˙b4�$>��9Ic�+��pB;�G�̖<.x�)O�®k�.藍QE��-�e��s[y�����8&�|���Jq��H���N��bPCAd:�������Ø��!3�0�#=�=��IX�� ś�k'��F�5��D
 5�8J����L�0	y�r浄R�������Y�S�%Vz���J�ul�e���9a�Q��c���=�fY@!k�j~�X�`Z�M��%8�>����3)��?ǅ{;�Pr	:��-h�e��3�.S?3�%�#�&����+���IW/���e����y��Ԛ�9k�jd������{�	qX���\�B�56��8�c*il�֡����������呋1��(�%h������"R�K���K�/n�R��]/��?�[ ���<���^RF�sL����0'���#u�B�i�b�d��mwbّ�:���DbV�ނ�(���
�����%����ߦ�Q0;9��8Tt�vqx'�;�}��`�[��ބ�w
��$QY�u�M�E#���T`���
�1<�"���'�)�.�M��n���X�4��V���#�&�*O���p��wF��;j��;�u�V�*5ٱ���q�i+������̹��
��l�rǵ�J:rm��8��d�9�[w��v^�0��렑-�sd����k�=�p��Pv�~@/��8s	��B�C.�`��[v ���R�%,��cJ�Ϗ�vi�5�K���z�04���P'�jb�PO8�a.���9O!���P��^5.�%���{XKe��J�մd�Sp�@-�;.�N�ע7�g�a�<c�0�`�d�f�B��U[9�,&��R������2mΌlIbhr�a���8���@��F�dV�w����P���7��]���
���1��e�@�l��(+�LN��&ae(}8��?���	 нp���W�X�#��c�y�G&x����3	�x�r��V�rJ|�_r�|+��Pt�݈���
�U�-Ѕf艸u��̮z��D'�-�^T#��]����x��h��!�ZQ�!!���G��X= ��K�X<����jBǫ��т9����:5zr^y!̷ش_7{>���!��s�8�>=V˖Af+bf��@�_Y@է�������5:IB�OǿlS�^&�o�V�H`�梬�#�c���^v�ݩ4���L�["E�cÅm#�H"�`�sW�������ү������#'�ܥ!B�VPҁ�v����H�Vd�����͛f�ũ ���D���f��6�n.�~9�bï+��%����[V&���{c�������t8�?8�6D��1]���|T�-����#׀9XѼ/�~]2�΅�"mD�+��~ڨ�7Ex�s�]��vr�t?�����4��=a�;F�X���A�D��Vw<�c�ih�h������(�3��O���o�n�@dP$F~w�XN��"��O�c��1}��|1DG�ڗ���T-��Z���H]+���PBi3�ݰ��Wց���]g%�������	q��K��(Vo���&�eipM��8G绮[a#�E��f�+]��3�V&�d��).;�E��}/��Ԛ� �<u��5I6��������(��lo��r���1���nJ 1 &Hݨ6��-z|(��q��9�Z���w��b�*#��7@Q�{�f�Mm4&����k��_R�}�4$��C��Qu$2)����B*]��? ���~�@mضh� ���:r����5+�ʕ|�p:)�+l��9ʢJ��[�v7.�o����m}(�o��U��P���C���f�Vh�����A�]YS�A&���ȹ�y ��ĳ2A\��ƌ��o�%���4CMέٯ��Ե�V��riQ�Դ�����3�\޻1���K �\�,�<�#����S>.�����Q�4Q����-��Ŗ��ZV�Ku�q8rQ��:'#���.�7L�J��G��|{1�4HR�Gԟ�nI��߄69���n��<�ڒu���Z��!�kw���T�����AJ�Q8{�3,�����;+1�+�AYd`�JEϻ|tKr2 ��A@��֜bR�9z�G񹁨��C(\w\����.�l��c]�==��|���a�[�-g�*�l�߸"I*��?�A��ہ��F3�Y�I������!C�,Ȗ����.e�o�5�?s�4-ܘI���3ڏ�H0�݅��!�$,�@���%��N���������@q�7ț��9���Ɓ���UI=*��a��ٚz�և,B%}�{��t�&2
�G�TT!�����笮6c{z�V����r ��ȡ��� 8�c@e���#�^��<�l�œ���m�!1˧E̵��tr>����)m>�&_}��fa��=��똶(��qJh��U[�;�k0��E�9��XS�����j7}�A�ɡWO�#A���!a��8�4�/�SKz<�~��������;�2�]��q����9�9M;�����u����3�q�f�b��D!]��)�Y6�s�G>�Ilٹ�V�kp5A:���H�q�c�|>�BE[�]"i0�7��^*���$�F�1
��0c�@�YLlh�'���C%��`���c�R4"&��K���+�i�03��Zh�H�^��eYǦ��������v�?��f>�9iv�"�i���'[͹����}�J���h��K�\��`a��wOzg|��s�A���B�
�;�Y��v�T��fJ.�|��G\�pQ�����3���Y]��tD�JKz����	�]�g�Ҕ)�4�
�T^�F�!���z6��Kbkz�Z��u��j7��3��҃
��HZ�z�rZ��0z;�q�խ�t���#B0Y��!� σ���2#�c��ת��`�օ �0s��y������P�x
�'9��aO�r@�pm��6SF�""�޻��V�z��0g�Y�;5��$�(w À#V���A) ����~�q���8J�l����Np<��n��4�EsE�%�2�s������v���@�����2��A�/1��j0@�W�;��)��B]<dr_ s5�O��|TO1t��p�7�N�b��ৢv�l�)�����i�8��MCگj�b��:E�2g� �U��D:������l.
oњRM5q���\��D�xG��ēZZo��	�|~~_��,�p�)I�H!f��5��hw�}ۗ�f�B2��?��>���w��П�σ��`�����C�C����/�9�&�F"\�K+�+���f*&��bw����d�!������Q�im��-�8�)k��t��S#<�OY�wTx��+7�o[
��ϼ%����pߵ�[�-8l����E`����?�e�{#8�&wCFuu6t���EI��cc�Մٰ�\.�9�S�|��;¥�/t�����c�Ԑi���7z�kt����p3kF�L&DѲ���G�с|zߓ��'�cV�A�������%����nC(
P��7"I��+�k�R��SB�ۼW�~V�@sg�d�� �&�������x���1$#�s��0&Z�$N���iԉ<��b����;�εq?� L�����L5̥ l:ҡ`�r���X'%�����k�f_�F�ִ��J�v�g�Ґ��pg ���[RH��y��\�~z*M��ye�=�z��X��QeץeZ��i���Rm뫚���!��$��	��<,�m>]7��7Б)'J��p�"��Z��e�H��kB�C����h����,����MYc�T�]�}28]��l(����%�휟Sc��y(�~�J|��A�EIڱ�ڳq;�M`o�C�=Sܟ�7�LV�?���3|��L���Y�zw��;��v��PˋC�'a�<�NܪI'\r?�_�X�O�f�<!¬^��kC�TniD�M��+"Q�D��B]�����?����X��,�,O�}�[��G59��Ln@E����U�LB@��}!�Zb�X]З�z
�����Ù�^��@��7*���V�}]�O�`�.TPb��[O�m�$]=�ǻ�?Cl�����jLc���70�^X�Hm��]7nVQ��Ġ�FS�n�E۰!���%��	��4Aa����O��-�N!�6+�����,`|1�aw�NX�ł��o"$��`5D�>h�F���q���8i�,U�#q�][잎D*e)r�y�l?J���@�:~J���$G!�����KR:�rrQ����įiq�>9����*C���|��c� �7�N��	�T��>���?e?6�����j��}R�wA|��sjL��P��j�D�h���_��s�r�3c4tkr��ja��L.;�����@L�ܫ��7j�X�Ǎ+������~�/�E��ů��qz��c6�_4W�)w�h{�y��;��#Jw�0T�o��2Fd���8�}5�/�KM�N��H����\.X��$���}����h��ڇ�6x5�]��O�/<@V�لd1Yu�/�&�o_x�a��:��০܄e|}�*j�6�Ф��J���>Ŀhċ�sML���,Y����-t4�����V(�T�Yj��2��*� �yx�^U��L��*�H'1U���)����l��r�0�d����i#�߬��<�<K��v�������bS�P�a��������&�b�x�?�QҪ�a��G�萄膶��WE��ǎ���w���eyGBIk��JE�ǅD���6E���d.��x��$g?��7MEBW��KѲ"��+PK��H�"��r�j�������QM�(X���~���n-q1���T�F�
��{�L���-d��fŭ�ʶbX�`p}yd��	=f_��N-x51_�Z��
����~m>
���6��[
�ӡס���ٲ�^a'����g��*��*N��匞����#K�+�I�%i�&@8�g�Ob��m-r�%�2�vNQ���h�-m�8
�"���q���r�7~��f��\����oӴ�֡��J������0<�&�wYL��ٟ-GR)f|��?�]ǡ���)MD��N����g�th�F~bfP��ɣ]�l?2@h���g��ʲ%�k��[t�Lf	��߉�]�CiX/�0<�ў��MI��X8G;:C���������l��1`zIƔ)���z�n��h������f�U�)�H�Y	w*/�l���{��lB�z����t��G��\�a@}0	��+�z4��F�2πE�v�.Z�^
+z�U�ꔭ�p�\�x���"\����}�:#��;5(���K��:8q="B"�`�|X:RG���Q��_��3�[_���̸�4�a/�9�Cʌ��I���� �W$я9Sh:�����'5�J|+Ԇ��m12���������~�ʨ@�"�6Բ�A���!!��Ruo�,c _���������W����T��/r!M��.�n-�~�^�+u/��[��1��Z��B�k���ZbJ���t�����
�u|�*��:���+��qe�V���6��������0"�/����AY?�����@����}z9 ;-Ŭtx�=�*�R'k��_�xp�:YG&�g�`�Y+�Ӹp�n)�]%Hʚ�����ȯ:غaT�ke�iu;ɼC�G`fi$#�����rnz�[�Hv���h���P�+�L���S�[pE-���g�}.�`����t8�DY���&dif��z��;x��=ܬ0��.]y���4E�J��,�M�,x]R�=4���C[�u�	 ��� ���*v�XHe��={�m��v ��u�ʽ���
�Z�U&NyK�v}8�꼩'�!���<+2�ƴ��f��BI��d5�#�d����3�*8�x�o��2lLi����khAx���5:��c���п�3ĵ�`�,E �D4C����"O+��K�?��A�ը�H��pR������8�����sxt ?�Y�����^��W�y�9�)�S)���_��Zl��P_p$�l�����R	8������5M�3ZX�><�;��u�^f�����>��9nL$՟�ƶ�z!�9��jH(���h�ӽ��Q�Ȃ�ɹ�����M�9ǠE�3�O��h������	[A���e0�������%�*�?=4���G��OV��j��h��� 
Q5��?ЅL.�0��O}~O����֠�^ J��3��>���)�]�l�PJf�Q�N�[�q�Ѥ.��Ok%ͽ��(F@&�d[<�{
��,���rh"�]Mq��x�a��,��C�{�Kg��l���G��#ӎX5L�ʡ���Lx����8�9����	7x�N�`�d-�W_�[�#]�ɽS��L�w�#�>���2��ף��Y��?i����x#���n�Mq��8�zn����YJ�p.�t��@u��SC�q�94�Q�g:�����ͩ��`��z�~�wa�c�x"-m@�`��Fi�[�{�vX�fV�
��梦��ie��[��|
�҇Sm3�F-����z���(��������i�����r#ծc�b{f�v�g�]�4��>��b��/��P�[Zv��i:��(R��ˣ^�c^����(��ֲd.v�|����4R���Yّ"�b
��������p�v~<� ����4��%�
^Y������I��T�
dH��b�+�=���`D�m�AXz�u�L�S:_� ���TBp��n<�ي0�K֌)5㈃H�Ӿ��8�E,:��v�H�k�N[�:x��.�qI<��#O�<��}[ �
Q���%������-`�(Ȇ�#/M|7�e5WT�S���������@��uh�o���b��1;��wC9�C߼4�#�0P����\Q���@�،4��QAE` %���4ه� �Ŝi_���	]��P���l�����9�ەo�=2c{^��`$�+��Ct�i��{X#�e�V�O���H�"�Ij���p�s �>�����l�vɧ����4w�uÓ!�wI����}N��E�q���e���zo���$"�,�x�¨gI��'�,��K[F@���~iR�����f�a:�}\�<i����j�� �V���;_�DJv,���D^��x^�g��!`T1�vw��r�����O}�}d��!E��\U)��2��[����]��J[eؾ�0S�D������``�d#�{QcHv�A�e=x\K��jY�͞���_=� �}UT]�����@i���ɠ:$���L�E���.�����N�*f{:k�C#���m���{ޟ�H�vdV���'�s3�b̚w[��տ>���dـ�n� ��#"PJۃ�3��{�Ԓ�����c� 5�Ճ	���@�J{����5���:�7�
�՚�����O�`��+�>½W�p�?I�Wy���}�3��#s�ߣ��������a����fku;�p;e%�M�~�BU�S�+��;c�"�VO~Npf��/a�92�F�P%�9��ki�rmF�酋A�a�U�X�� baph�}���M���$)��(��1�jy�,�W��scf�qA S:������p��!�;�a<��9�M,Z�u-��e��J�y�"�)���-I_�l;�ǌ#�/�(�|U��>N}Λ���'9j�i9� `�t�@��Va, ��U����U?�tt��|�>=�����ʞy��!��z�u�G�!W�V�@Y_�kZ} ���H�<_�|̂ה��fh�ʮj~���![������)��v�!�@`0�a Z���>�=�u�{]2��|<�#V[�'}�3�����U��,��M�\H�):j���6RΜ����њ��r�)ʛ���4>}�S�YF��p z2�m���R�W�~%�]%y��}�SL����kc��=���?�-��P��m~si��11y�h^fINA�*E��C�i�1D���|q�9;���L�4kG��݉qu�8N�hJ3����8�AvEc�rU<~|]P�%`N1���?b���
�����|m�Y��',�t�"p@r̟S{y���\>u��Wi�6�.���L���c&ö/!Dq�l�pp��o��X5P0�4yO�)���8�':�2������v��)�rK���i�`9�^���^<J���:D/�}�>w�$*�2�X�6Ux������2�.�|�o�w����LI�Y�ﺴ���x+EV25��w�]�J��>�����|A����k'�}v�`�j7���F;��C��� �a�~��N�^7u�3FcY�<ȴ�<m-F�PR�������-��$�k�/�v!���F-7���)�3s^r#`7J���4�g�����:8�]rdVٔ;d/�`�b&�Ŵ�Bc����/(�L|t��q]܏
��@�~��ι�L�qҭ�s/o}iZqN�x��5M�*�Q|�x����Px�M�nk�N��UR����P*�����`�RaK�G�
��������ں��)�Q�5�:�[����� ``�o�%[�oN�%���F�2:����
:k�v��Ś�����>�)T���TL�VC>;_��4"�_�r�6�-���ͦ�Ou�0#�r���u��B�'��K�f�f�E��B��c`�s�4�	-��f�K�T��?5�i������اS����4�cl}�>��|D&Y���F�T��0��S��45oV��y�i7o�n�p4WG��Sl����E:X��S[ɑ����d��A�9�����Q�!'E� ��+�����,R��)���(
��J�'6��zKv���3��~_Wl[��8Ź�-<��`E�y3 e�g[@,j>F���/d�P��2�5�l���@b�0�ޮ��+��Tl�bO���4���A,����(I����gil������Y$|I)��%�{���n杄d�>���c��w'˜� ��qE��j��Vb�r�u%%xq��ʘLF�d��.7�n�d�I��2fD֢&yD����M`����6��B��UE�v�
�F�#GI��E(�Z�<��W�,K���͠BX+M�Y�a�0ZeC2���3^��o��Y����m�E�F�D-�.�q,Ήۤ����A5 �0���mNsG��4�^j-^p��1A޻Cu���������p� 
A�H� 9��u1��&�	�Ԯ#~nG@����L'�����D\���(�&�L��]i� ˸���|*ߜ�p�D��դ��hz�vn�&ַ����$1\x����~D�ܴ�����PIbv^^lK!;�k���(h�e�8��FxҤ���M�2���kP�����i�S�P����^x=t��E"%#��jc��6.��������w,�rո�����=.�~k�,�u1*Z�Ǌ��)_�%Hʚ�:=�uɀ�K�{����+�S:~#��
����B�ۻ(��L���I�x��~�fn1^,-)w0��	��R�}�[�L���z[�M<��6`���Ӽ���[{�J%��5�m�KEa�nu��߼	�EO�L��i_�D�o���C��ŻiY2Go������,D�韀;d0D�^}���:]g�#�5���U��b��Xʚ��t�'�)�	�>���6�+�V�Q��(Ku4- 9Z9;DQ�>m �h�|�i,���68�����!��[0�_�/[y�f<g��Ӽ��l�Q�7�c�Ϯ8�&��]��7�v#o���*[K�P�K?�#�nb���c�%-�TD��~�8�G1�{�:f���~&�l9e��)��6�3l�&D�n�y�J8�i�(d�FMQT�z���LyU�Dx����5vX����V�۾�>HOI�	N&��X��߶�rX��"��Թ�e�[mxOt1�[�� �Bg圗�8%<@�Ns�6�??=|�<X:8-��,m�F��nW��a���z�����`zEt1昜+�|���>Fc��B���+Mc�d)�α�F�Z��z�=�H��z�Y�*�/��������k?��ߗ�(0���Ij��f"�L�g���n�A쵪�ne�|8��0�'��G��`9�(�+5�����	S��M�0���t�4]���d��'��%w��iKn�td�HU�U�N6��{Q�8P�9����t$��2��5+bv�?�+
�P���p��.���Z6Ϩ0���6�v�I�X��2��)��i�=j���_Vx�;!	MBX�*W��͢%�s"��"��{�j�jo�eu]F��Y֯(�cb��B�*��MX(2-!"��7�r��+4��dO\�,�Z�j�@\,��B_}���ȶ�1X�20e�Ĝ���lT��q�cl����C�|O��+l�xKM���atVb4kl���^(Pr�ޖ��A���$[���lT!�n�����,cr�{J�'5s�a&B��#Lñ�*g
���5}�M��PI�1�@��KG)鎦����?�F)�F|k(�׉���b=
�zG~������f���EX�lП���mJ��C�H}Sma1{�W��lF�v&��Yp`���X�%�c��3���|PXR����V�zA�Ǳ^�70?(��f����]�?�������r��U��_�h�����&[
�eف���tp����w�Ej�Ix�A����g�k�5��:��s����JI+F5�0�[r�S�!����1ǭ����E�>���i�Ej��1��%�gre��0TF��U��g���ӭځ[�8Dd��	a�2�S�z�FNDp�ob���s��s@3�.f�(>�e��>��bK0uU��H���e�����mc���Uc�,�G�?��C�KT�% B��8hKa�҅��d��r�Fc\r/���rr�'9������&���d����"X��6n{s09�����!��}�@PC~���;-{�̙�z�}Y��R|�B}p�Y�K2�4�$�2��&��+�(��@���#K;=���툛_���az//���=s\�
�T��{��--_z�"���α��T��5s��m�(��q��`�B��L������J����p�E�M!W)��z( ֬�2����^@�#汋Dm�T]��N3��0�{^ԗbD:�&��5���.h�[�fC�"��3��ta.�=�}(��;��ut���8�9�Z�j<p���2`��l�^�wG/���G��Q45�LB�w\�4��I0�C�d�ld�H&�m�� ��w�>���.�Z��2(f�,����s�iE(?|�C�&�es+@X7�`�mO��C���tc�X��ԤJ���4��|�����=���n���Y٦:�Xl.}Wq�
n�l(+�Sԑ�믆p���~L�:��܍��f���M�q%Q��CW:����� �xMd�ݟNm܆[��jy3�j��&}%*:�fЄZT��-}�K8} ��'��]n��
 �rH�C��[�
�iE�c����
}SE����T����{r*��VF�#��S��hV�ݳ"z�+�ߙ�

���~�6[|pc%c"*��!ug	���$�@�	�vU�{y���r{�D�|T�^�&zZ�d���ȍ�í�h�/�)����9�N9��È)��B�	*,��"�\c`���]0į�+�)'��3n��݈��:�:���V&R�/ZT���xO�8��X�#��;�DMeC�@N��
�|7%����z��o-1���7ڼu�(C�ާ�B���zu�hg���ym�%�i<K|AR�����S{��[��<s��b�d�#�"0������%X�+p�JZ���8Vu�dD1�nO�ۏ$HD�q�*�
l.�-l������"��������jێ��w�Y����<W]6��i3�S����/)�
8�ƪ�U�K������;�o5-?�y��\�m`O�Fxf�����8��;�r�u�A�Ǯ*d�O�)]s�x��(ɵCs�#��l�O���\��}�}�ו�s�h��WP:�>��N�jG<���h���	xb�Yq���Rz�gi����f��|��d*�_pW���;�h���\4"��Μ�;!Q���~�|��E�����OU�of7<\~��Tʡ�ve��]�m�o\�_�m<cY��̾�VW[�򚻡�,��f<u�v�%49zt����(��ɔ�{�¡��=�a|=l}0��z��
e��kB���'�<�L_�_M*=[����޷�Y�%�apB��wΤ���yWi�2��.��#ܽr�}Ѯ;�~�{��8���]�La����T�`#���S�ūh����Q*������н�Q�ld�5a���7�I��ҵ[r@O�V���}E��t�R-��x@�͉�'&�tW���9��VO���/�-��Zy�����g�����U�Z��!��N>q}�<�Qg�^�zp��}��pt�)Q���L#���=�����t1�@�?�,CHf�����@�^�7v!�)�]IE2�Hw�JM��C������-Q���
�a�}��R���*?�uG�����AK?���ܖƅ_��f�>�L6�"�T+�$���}�IAj3�X�C4ޡ1�쥲W�j�7�s���3�����]���%I���o�1�}]���=a�?؄}w24��y�������~k2�9��zI�<� l��x!�p ��{:h'�D��o��i�C_��<U%��Qpq�����,��rl�-$).x��uNp�*���_�y�1/�LS4�v?M�by����Gr�}�a���ڊb���!���H�G����ESg������e��Md���-	U�	=�8��2[UI��7r0/��܉�*K\���$����JT}l�w�Q��f���x0���b��mϾ���~�9����X.y�M�̶<�f����C�	�Y�f��JJ�i��o�UdN�8��B�㒫�3��u�_�S�/��@9��sc�9{���`�E�sS->P�{��W`)À��v`�,&��T�驏=
A��Yq�V��6�N�Ƨ�ܖ�b�x��²�6 �gՙ;m��P�@��)+S��u����f��@�����)���x�XC�j�=��>��������X�����tg2LI���D8���Ff�`�f�<e�kyh
Q^b W\��)!鍡#��~�Ħq	kq��H��:��������YX	
�DG2p���2A᫆7�����f�o뱍�s��6�iϮ�п�����P��]6p��%��9Rٵ�#���V�H|�I�����e�����Y�֝5 $����&��#qI��|��� �V�*�$� �����m�����1��W�B�A�PW/68H�jRUZ ;��c3�Y����.�-����B�!��)?Z��������q�C����L���J�8�p��{�����KRFC�7zd�~��Lm��g�uF�%�h38��)�C؝c8��t��]o1��q}���)w D�s�͉��S�>����ՑB1oD��f̝��N�/�o��JTbN9�Tn���f�ˣ.3ˆ��?���A�Ć�ᑑg����lG�� 7*�[ڄ��#<&Z��$�b��8���/G}�kڵ���~d��T���3��"�cX�9%k��k���&��~:`�R�+��Z�B������EN���~�9}�n�Px�EW�����Dm�@2��+a���U���46չ~�g��jo��~j0R��.�F�EKh�#`J�����C+���0<,�+�x\2e0�005���LP �R��-K�w)��=�q��N$�v)<�m\���>*Y����2ZQ����B+���W�i�#ǣ�舢��]����Ҋ��;2��5�3z�S�X�5��������u7]�Ay6��>�C�z�/DU���c����:x�@h�W,�*(O��9U�ZO4| ����vr Yy��5g]˪d�&t���#+1�W�,Γ��(:��q.bZ5�if��c���L��7�3!(2�lx%�s��,����(8���́6*�r����u�-����*�"g��/$+!j�j��Tj��/�^do�I#`{�;kp��gJR!<G��N�=A{���u�-�h���/dJ�,>!rL���"ƁI��c/D�T)��T��!J�r?O�wϻ�no�;�-��uط >pB{#�u�<�si�SR�) ��'ĳ��b��0�o1��C	�gg4<p�UN�C伍�b�im�#@�U���YS��
�&��`�k��A{��ƕjn/�
9�d����t����$���V��P��W�+ᾖ�R�DF�mx�*!�q�a����UE�r���Hk�!Oa>6mYj$����āǱ *��'.���`/�����8\"���4�ba����@\=%�#MPN�Ӏ[���^������b��0:6�-��k���pS�*lQ��P��(�v�aT�p���;��e�"_�>z�2�s0�\IdP�K
5���EeM�2�_��i���Eɐ**rk��zpm�Q�F�;������Cv}g8u.U�R4�[��.�m�8R7�Т�`7yS�4G���$mx(>�4gGȻ�J8�������

������1�2%_�uo�*	� w��2\��U R�sN��e��r|���&Ǽ	�^F��}�?b!����JQ'Ūן��$!I��4�7C&���>Q4�P"�ɣ�K�N���Q�ќ����^���:������Q1㡊P�0���U��]�Dzܘ������;ݟ�Q�ܮ�m�(5���~��H��d���a	"�2��B�nCCR�*�t��K��QE��8�9��X5��}��ULtFo^7{{^`�k�g�L�=�$ A�ӰI-�n��%qk��n��4��K^�D�{{s�(R�tI��3��Ӓ$�S�N&���6w��|�NL6�\xT����$��n�
��=k((�z��F���FK㮅t���z��Na~����7K�3�!�̰���K�.ݒ����`C�B� �:kWZ�1VV*lLژ�!�E���]7����ԣAh�NӔ�әsՔ�����4���+̓��d��W}���cY㨒9_gK#\x�"<�����ψ����%|W'm�Ό���"���K�.�14"y�q��N�!�޸�����.�=b���<?�G=��ެ}�S�\5o� E.������HS�T����^V�@���J
�Z��YBh��R��Uy_@V+27I�����1�1X,�n&Y�Z��8Hr~z�up��g�*8w� �2��גb�]Byf���?h8�Q:��>7ʷv�f*8�LI{!�=��Fj��+���w������D���p�ŏ��d�m���g:o3�*�v�`�8Pc�� Y�(��.R��$E�I�A���M�HV��&����w6�{�l�fg�}V23I���S��R�;�m n��F����u���]��p!�KY�Ex�#4$���4�=����C-c_�1 �Q-��Ƨo�u��v�)9RjM2mo�+�i�[�gy��U$>�F9��IZ&���*�N�0��$5}��>�\��i]&� �T˞j�-"��4j4e�D���z�:��*6��j��0^VT��:#�(К��F��q ��x�-|M뵀�]��V䀓W��bn�\�d�V����dJ�3�UL!�ǃA�~��5��e�����{8�P����(�5�/ܡN@v�����GC�}n������.��}�)��P�c-�X�����I-_a�JWш���91��!��w���&ź!7�:ּ�t-��e��n��j#����9o,��J�gVWy���n��,��&ŞKi̿��!,��xrL����v�m���UݏK	�ȞeR��n`�䓐�Cl�=6�N�}��< ��{	_^���o��t�e�J�/�=~9�*�i2����_XWq�V���W�@�}��B�g&�4,%��L��?��7� 8Ƀz�J���E	���44T�n}����?6�����j��O^M��fH/q��U��@��1�X�d�@�q�)��NH%�����q~��'F�[F�#�<�����[*�1�#AQ9�e�Sk����ڔ���m0\��4@��nw��K�g����@H�!yW��
���}�}�S�X:CIW���?IW.��'�u�6N��k��M�\�@��Z�"Ils���������mo�i�R��M�^�k9�����Н=��,�5JN)����no�i`�n�d,[�p����Ϯ�ޙ�"D�֦#u�}6Y��0PC;ň�n���`a��a�ӚJ�y���  6O��d5�{jE��+���9�x榖|����0n=wr7���].B��fX�Ŭ��������z6�&̙�=ӡ��}�1�{$�J2�n�����RK��/�����OSX���W0k@I�lM;�#d����ʔB�3���G#�Q��9�L.�C�6
�_jj���e����n�{��q��H}D;π������#����Ayp՚��$���k�P!v��m?\�k��ߢ�62I�)�i�;�O�k&��4$�-�ײw�;֎J�Ū�{����u�X��q����A�ƥ���GI�����(�y뙽�Ҧ�&\�Ф*�u��)���X���q�KI�SIU��{6̥��c
X�fm���Y
U�&W&�A��2��n�4�U�\~����B����"�������yT˴�ڏ�R���fT����nr�jJ(d��B�88Λ��1���γz������J.�t߲��.�4��4��)r������<$��H.+~(��A�P%�/� �8�©��`�%[|O�<1�.*2�YRS�r��׬S�E祴�O�l.$�+6d��T��,�n���x�k�h�8`��>�hR1�i��ZW�3�Ѯr�������Cz2ə�΀&�Ī�>��Ta�ۀ�%�Jgv����rNB��E��-��ʱ�$�'1ڣ:����*|��t�����j�K�s��G:KLI�b�ηk4�������I���9��-u�.�3��)�h� �� ��LL��W3E6$,���l#��*���[��Ļ�z�U�d��*D�	�.�}���d R����R�a=�Æ� ˬ��O�g2��D$6&`���ph�s�f>��p�C_�͛�&���y�Ҿ��c�d8�/T�Mޤ፻������L��S��O��Bd�A�9��ü? $h��t��JE'"����>=�9Ոf�?���`r���}qz���=��-!+M��"u-M�i�
녺���H���|�� �!�&���)��^#�+l������s�Yj�P��M�P�{A9���T�l��s��ʺ! __�����{=����1���&�L��r�8�D��6���Z�6�e��)h���aAZ��{L����l�˺�o����Mf��2���،/��������[������A��W���e՟ڜ�P>$�����厺s��tw�3�Qh���S�	S�VsW�R����X��o�%Z>S<�M���nƞ�d��B���h�
������7`�T�k�����;M���_��e��5^+�(�-QWm���K�q�#���,~L��x�V�1�m���'4�)]�'F��U"�:]bkg�Y>�ܔW!�L�*)�1�aء�.җ^1�Շ��k��CB�z�(�|�w�cl8%�9��r�aӑ��R�0ES�rV
k�Ϗ=�D"�b�y�Vb]K��qj���Z\��o�;Nڷm�?!�2'�p�7���$����۱{#(�3ތ�禮������/kD��1h� +Af_S��.�O��m�nʂ�$d���~!mac�2$�תB�Pϛ�K�����o��46#����/5�Ȫ�^���G2P�ߎ�P�������y}��k�X��|�W'���k�VH:U��E��=�4�
Mjq�{��2��ox�O�ȒYh�/3����xE,Ez����Z��zR�}�?�x�G�]�5���0G��)�3�(Io'��(����F;,#nfF�&�m77@�����c�
�Q-���8���r:�șk��k*,D.П0%�qYZB�䉇�
�*"�+�i�e�i��f�?�D������o�\���{+1��I����*`�7�s�Ƕ��{���d�4�!B^)8=xF�<����a�i��บ�"$���ώm�Ve&�,�h0�nu����DU�
ǫ�B�`�p����Uo�A5������:��*�C���s�%Rm��ڹ��l�J@��@����� ��b���e�O�5�M��e�����+��I�#溓8`J�����pSZu��Л�ԕ�q �p���!=���*v�_��	��l���*M��0<�=��&e�k5 �M�z�ӣ�I+��r�[����rc�,mlܜ�`
"2��4kr��1Uꑗ@<�g�A��|`�m{
z��lL܀���p;��^�F��]{��Ë��cO�S�U7����Sß�;b��d�������ٻAE�5����Ӵ˩��f���k8���E�z��2��M�w������x��G�WM�4Y(s�bT��&'���d�Xp�=���|��i�윮���O�53��t���S�xXlHI�� ��7}l��)���o��"?������
�����>�x)/���ݱ�z��B�s�B~@����g!*�����[%��zss@XA�5��h�rc%L���wi`)��ԥhCF�͈O�3�9��S�6���{ V�P7��w��Υ�F?�8�5��~�1�H"k��H6������
�S�ɂ���D��OE�h��|$��"�g�7��]��*�GR�2�g�v�n���9�.e��e�+`�sM�{jkF�R
���mHCt�(�|!� �'������2nn�����:��s+��m޵�3c(�G��)#p������L*2 0V�}�xP[����`��`>������y去U�\�ș,��5����Qy�}�8Z�L*8��)]�b�󲶞&F���[.���9l
�Gp&��;wlȝ����l͢�R�J��2�����d���j���C��#)V�ZF\�-���xp6�?�b!�j��B��������7��N@5x��a����'���*d���j�� u���o����Σ����|�,�ݒ8_ٔ#������bLB ��H
�.�.�x�Gj'�����6Xw؇��v�b������M�@�� ]QS�=�p���y���C�0͆8��a�9�e�B��6���[3v�vo�+�+��8�ꉍ;��`�'���{�d9�����o3x�KjI�3�Ԉ����VÇ��tn��p��U��=�R��4��|�y^'jₒ��������>7s)��V1�,�w>��~�z%1{cV����s����d̵����&F�f�j�m{-^&�BF+���ZU[�s0�]Qj܊3ۑ�b[9D��^���i�<?�����N?X�����\2���z��PP�y8��׍.��?9�	f*�O@Y_��Q��u]i�=݂XX�_|LY�	l�Ly��p����52>>���V"x��jDi
)I }�#��#�,4��:�����i��fM�"�,�j���:��x�b7D�^����H�m�c�0,�=c\
"ͅ ~�����P�sv�#����5k�/�
Z�R�
95/���T���@�Î��뒡yPl�(��:B��x�b=27}�=��{9b�6�ɫK܌h����zș�D�� �J��;5yw�?k|&i��-�Q'�]H�^�$�,��¼
<��Rגh sLI����Cs�+Ep��c-��O�@Ʌڋ��7Br�$��f�3/ l"�$����"����l)��tl\����;�G5%���,&!44����8�%��>�sY��?	(�L@�R�͕~�S��>�$��/AF~fIЫ^�v}�}��?4��N𮞩�uN��R������}i��#���/�_��.�M#�A�^+ �zr;�\��Л$�6�KOV)�V�K��Y�r���MLH�I�pf�(=,��Cx[��_Rz��V�y�]h���i��G	��Q�h�v�p�&��.[�k���ʛ�R�$�}����`�J�i�-'��P�Ԑ�(S#y��~2E���C4�@�_7r��$��)�R!�[��8�L��X��*9���á�?���	3p�dճ��2SoK��be)��ZL��_�ׄj���&CG�V�r�OP�R��}�&��{bZ&>m�xl��e]i%���ĕ�WS k�쇟�� G)q���aٛ��j��A/���PN"x��������|Cwo�|/�t����_�Wҽ|�[��7���F�og"�Q'l���	����H�+��!]UR��k}e%w���n��!Sk���y[�����,˽t^q8��#��m4:�[�E��r
#!�HL����� �e
 Dg��%: 	"�:����pn��-eE����y~ֆ�m�Wf$ixV%��o�[����1_5��������ط�8��x��~���Ba=B¡�Ǟ�6��c��4RL����-��Y9�*�����{4J2�p�\������lԻ��� ʪO� `xT>�W0��"O��p��r��_���O��[��f!�M�C�a��4�e��E'��� �AH�OW�X$��#b�%�=kS*�tiK����*J���F�)N�(py��h�$��ՖP�i��A��F!.�;Tm�[���t76�N(�NG^�����6�ڴ�{V�//&'q!ۧQhGpו�a����@�o���1@"��x�g���*�ْu�RJ���R, �ˈ�N��0>��������^B7�&p��|J�G-r]*��7�Kk���Շ����L7��1<�Pr<7@I#�2k�W��0[)�S�J�<�Nrǵ�!�v��g/Hgg۔��P�=�)3�8�-�4���`���t�����&F�Z�w�˶]T�Yy�lG����[�}+�c���-o�?I��q{��ͱd)�*-|�V!PyN�3�AA�	�����0�(���:�����.,���ʴ5K�����Qm_E%2��5较8O�rX��Cl�gPe��92��<�����<k{Q��y�0���7���1���֚����G�~3�A+�n���x��BVB�����4����[-�� lu'��'���[�'Ǝ<厜�������W
��L�vߺT��y�|�t�V��l؇)���[�e���{ ��ˈ�xw�a�	�=�q���U&Ԙm���N�M\���c[(�}�Cn��(�,<,6@C��'bM�`	�}�Fj�^�T� �Cg�)Q�`E썮F���O���SC��72,�$'Pi�9zx�)����A�\�f͆��b�nr�ĉ<#��AA_s��u�f�q��}L6���8�1��-�AF�X��j-f��}��-;������1-px��� s�z����~�s��3)���WfM���7�r�L� �]-�3zwr.�o�u0!f��KD䬽��ǀq��H�l��;�0��ҳ���9pH�Dy�������.��%gM��F��5>'D�rT<��L����x����t~�Z'��:��	فȌz�g���4�@n�����R��f*~���v3�>O�H��R��H� ͅVސ�2ң/ڵ1�ԯ���j���y��Ӆ�|�������h1��V���I7�g�� ��1W�U����3J	[�,��oN�O�ƴz������>��"Q��/�f� ���K�^4�)R�[��{n�k�nc�[���&%#հ��0K�S���2�?���r��}��*�i��?S��	$��Ӛ�^�[��Hd���MJ���(8hS��!�2��=���i^�[cq�3�����Z��.�9���u�N�=v閵�ײl��5��H��ֲ͉�,lI	�n_Va��c�*�Cz���.E��9���J���&�Z��TK�+e�6=W��|[�P��b�YI��?R+�?'�����������r���t���	�������K�MBm��|�\%��"���Q
(,cX�C�I} [�|�^J��GMv�a�T>��&�Ƃ)��Xa�X*�D�����j$(���F�~�ڠ�`Q-:�/:�%v��f#=i1+��r 쪵=7�uE	����Nt��2����m�B=|��Bk�0Ǣ�9x,G��A�9B=��.�� �:�mJ
�mo�������e��3������� `����m2}a������"��C5��K�<�vJ��@���24/���玾��p˕Jp�k���4[t eKd`�����5�,ً9 �E���Bb�#�+K1���:����N�G)��򮩹�s����-Ӷٙ�6���W�o�&��b���-T6�M�%9^�"��W��a���L�Ɖ'��n��XK�O?p7�`�Bm���nd�Y���j����\��o���HB )�HF��j]�Q��?Q�H�܆B�%�p�'z�T;
Jd�y���u5���1�O^��cwK������yΙ�L||��0s�9��:_�g�������D�f	��|���[���{F[���P�7���+˫��FT+�E��Z1;yUg�wHJw&x�n���	ɃR����ʟ%���@ ��_��H����f�"��b��s��ϭτ'�ơ>{��)��>���ז�9~d�,�֌Z�`�椔	s�Kz��,1�e���>�8VJ��< :����l�¿����FI�<py�<L�� ʁ3����l�xޛ�k�;�'����T�C���̌-*w(���aс�>n���ơ�mh6	�H>s�@/��"S���j��w1exe�/�d�:r����&���-��Z�Ev�����P�����oA2��P�&�(W ����0�Z�,���醈M6��X�x��F��N0�Y��7c�ޚe}�Q_i����/���/�#�0R*�H�2��}/��i���Ң~���
�{hd{9�yA��`�}�:��
 ��P1��/0�ml���JѺ��X<3{�	�M��f4bCb/DC�jD���M�1�P�;��ğ����L������y�$�kU��QC�sZ�Hԃb�g 2����I���."��!�R�I �o6Y�,���k�7��1tj��a���J� �.�Р�����)�&��h� �>`=q��#�2;;E��V1|ts7C�>�(T�s5'���̎/���«�pB6p|4dz{3�i�g 	-R����F�KK��C�S��g�O�Ї��/A	[��#���n]�Q�Ҧ�n�)����� ����
��跍�2e:K_�^m֣���,�Yu@�������>6�jds=Y�^̩�Ǘ�HXv\l��S[��fj02x0b�h>Y���|�[�'�}��"���n���i����h�y$[Z%���5a�/�sG�%��|�������`z0~�:Z:Tjv�ӓx��hҊ��k�~y����V��$9�g��Q3�����41y> ��@���@�eR��[��Kg�R"��pH��1ED���)c  �qy���6f �d0��o����!g��ON���7���	�%�+]�AP���h<���?6�lCJ���PQ��}�U�,�2�$�iH�gHr�G�k�b�/��H{�x��˹�H4��܈�ɴ��,������M�ZhX�㹘��9�m�]��-���{<�������c��K�;+*�z�S��W���{V%�7�e�#��C��^S9��f�z�������i��of�aɞ��ch-x��A<e���o�4kO�]{z���6t?�\oA
:.9�z�c��m^'��AK���<�K	���.FZ��Y*7��O-n{qX�X�x ����v�{��T�6�A��AUR���#�]��A�k�v�G^�9�6
ˤ�a���1?lǰ�;Tl��[+
H�^ �++t{\��*A9~x�[f���uz��#��m��H�}0,��d�Ad43�sv��0�Ub�
\���Z=~�<>�?r��1�	-9ꍍ]���_H�t	+ Z�Q�GӦ����&���֑:v��K�E5�S?���C6��3m
*��F���b��
+p15�3��&�����M-%ի���ك+j�9˺��g76j��D���<hs�ZN^;��.��Չ!�H�.�3��q m>�+�;�ϛ�L�	�?�Мz�k��zm%b�8�n� )���ToGf|I���mI�A�i$��� hp^X�KA"�9��DgsRv/ǎhg=�:����n��6���������g��Y�K�yk�A��ca#}ȝk���S$2�C�T��q��[]pQ��lz�iյZk>>�S�<'��Z���h:a��pQ3O��ٍ�`0pv?�T�A.K���Dnv���Sĭ�I�?Y�'��F�ɨN뷱�E}��cQ��Q%R>H`F���;D�,x+�s�-��T>�_ɹ�ٜ8yD�6�Q�x�>�5s�y�_+
}OW��\���/���	�.��駺ݧFt��`˾.��a\F������k7�=8�j�I>ژ^����	*AL�'�����䭌�|���
�`ޚ�#)�9�:�`H�@�L:Q�tNVdL�h�J{����-�t����]��^?n��APEFx��8=;n�JR�J�-��!bw	���_�X'��=b�������L5R-&����E�g�3�M���<�p��.�P�V0`>�C�(+�O�K�%a����Й\���|�z���V4\�VE7,9�mQU��T�7y�ey�;R�,8�gAR�#�>x"s����t��]_[��
�Q������m�ş�,����୊���g�t����ٗ+��C$CF�+/OhC��?,{G]���	Qdꇖ۱�!7~ᗇ�V��
�����A7K�\1�Z�~�k���J�iB�>�����IG����-�i��0C`�����QY�"��$Ɩ��(�E��h#,�͑�,ڠ1�BA������B�o���a�{��u�ԏlV��߬F��E�s�����Ea���'X䀍���w������O��j9T���b�G\~�!�R�����_�L��3����%��O&�b;���o���Â�9��8T�����ً�]��y,���)@Zf �ta��xzm�=��/N�`,�e�K�fy�Ѯ���v�R��`�q��:�|4?�ۊ��2.a-Y�Ed�,���~o{��/TeR�	����=�`�jV���Ô<'��r��d	�~�>.d^�
- G w��f�����/Ǒ|s]�o�~�
�F M�]�K�u�Fq�����X�(���׸�5�C��5H/�;ަ��P5�yc=~#H���� �Z-��ҟ��q���j��b5~�Y�+���t��\��[��6��������6Jq[�C�h���P^�4�C�@���݁ ],9s���f�h�Q���8{���2�+��y)n㕓�)��	�p���#`nE�̫ע��YiQ��{�������ap�v2���d��̷��5����7U��\�ե��D��:���wh�y[.`کxz>� _�w���'2'�e�;C�!��%pL�Q,
�p�� �sS�E��aS���B�K��k�E)(�������V�y>��o���?���C9���ZTna���s
S��5�s���f؋�|å��Lt�}��
���������]�� �k�d]����װ˃[�r&?Rql҅�����Uz��������m���	�ͬ��� �4�&)(ˆ�%o*&7���M�w�gj����C�i��j��4���$4 |q�ܳ���������M<��vŚ�Iaj"7@�{|�$ ��.�_3�쨔9F9<x9�U�HS;cU	����d�&�������P}����>�D���>ǹ}'9Px����L�a/zV�[���8��nHNo�tV+~�	�e�����{��ۉ��wk!���H�K����O��>��RP	![�Fv�󄎋8�pR �Z���0��4�
����!�7��?d��+�[��:�Q��<�G����4r2��2B0C�k���&y|1���u��7��4��@A�Ϋ�(yѹ�a�����QH�馜��� 7�-Q��\~p��y�s���1|�	�EX�=sנ���*�Ԑ���<�Y�����D��U��%�N���,ʅ�4��ػ�Qt�C�Ⱦ��ެ�i�F�Kpj)!�]��H��Y�,�	�R��{EI�[��eqP��a~T���dL<_(���YJ��P3~�9�~g׽�/L��g��@��XE� ���N ��]�L�7`cpG�~�m�P�m;y�h<���( 
qR�y#�]�ԕE��9ې�Π��Ŗ�˔���'�a�uҹ@lߑ��)������9�u��Q�����Է��׸d� ��Q��|���S)f(<�2�m��跥T�.!w�i�J��9O[^ �>���sf�U6�T�t�Lo̤�Γ7��yn�Tr�_��������`����)��OkHX�Q#^��.�*HQ	��g�M�k�e��������à!Y�AM�C�Oz7�AN�0B�S��s�/)�6����s��+�����'7�����j���ÊIѶ����q<��q��^َ�������s��L�P�2��m3��G_�.�ԩg���EZ�!j89+�`
�R`_ϑ\3u)
Z��V�Z�Y�0���s�fK��c���kZUQ�
8͔m*g�j��d����YS5�BzQ�Z8x�ɖ/�,�!$��k��lCy�bT�F�#?p��,�6�����	~B��iw�z�Q����L��B/�my�-���!^}q��0ޏ��Sr��{sχ*9���֨,��@����k�މ�&�+g6��s���M)Z���|�J��bx�\�礷$hpnK�,ݘK>'�����m��Ѽ����h}���g�n�?�B7bK �$��c����c=�ְ0#l��!�X�!#&j?Qh��`���&9Ӻg� :�����q��C&G%��Q�Ʌ+� >!	ν�.X��Z�qW݅��S���-�ou��H�3?Xψ��vq8��Z�ɩ"�p8|�_�qw�Ԕ<���4��r�������E����UW� �7,5��<c¥��WY�wͥ�#��:6d��O/�ԵQ]�E\���qĴ��!�)P��]@S����k�/v�����_QGN&$�	;�����yBwy�-�r4��N(�����w���U"�E݋\� ?Y��IȻ ���Ey�5/%�i�� ʻ���hN
�Y�^D���DMl�4c��/=����k�\=5i��F������D�O=��ܕs�w�!����áv�-r��A�z��8�&��=<ZJ��\�$���&)�
�C���7�{JȒ|/C肇ZWw&P�;��������(,�L�мltA�2f�7�Ƹ���m�R9�J�N��#f��S&��r��腐BNkDf�A���i��Ϲ�Փ"� �]Cڴ�lum�k��]-91��0�!6���ɗn5�Kc&����a�ms33���ڌt ���n�tm��+��s\=�u��j\ ���?�h���[��NQ��� ��$
��DYa��:�x�H��o3.�4JF��d�e�����-ܜ�b���:;'��i �9�%8��s�A ����:ip�'�w��C�|t=^4����x�wH:����P��\�A�����f��߯����<~f�4V�иd<��t���@Z���k �<��hU����� �n���Y�z��z�[�Io҉4�� ^?��v�Ld�ʐ�[3��� O�_��J�26��H����^(��O���t��Yqk���e@4 F������<��bՊ�
�+hR϶�M 7@��<*�mE������g����}a着��`�5�vc�3o����JdA5R����g���Lo�~/c�x�t�WG�F�ѣtd���w�5Z\�3��摀��*y[�8�JBQr=���!�j�Z�!x۴L��Y�A�w���o��N6���N��x
�)����Ҟ�qxƖbs��+d�]��������������4{�_�Z 0��B���E��([�f2Fsj§r�k�m�{���1(�<$�����9��+��ZC�Vg��soW�ƤCó�.V>+R�9{爉�=C?�%}%"r�V\t��ُ�m��Fl�������n�97�ZB�Fi���;��\�N���yGV� �E�������[�d���(�8�F�ttI�iᛅ^٧�R��`�1���_q�^�p��k�?6�ز��U�[TYv�����Vo��FɔYk���1�_2u����g~;�}ZV���P��n�Ǳ�1�k�M��K�(b<j&!�ol=��<�w
d�-q����O �	���}��m[���+��'�c�Gk����j�~R�4j�� ���3Tk&@I�-�oXߡj��&��d���ήj�8.�|���c��=B֝��r�%m�
�:
@��L2�D��9�6��M�	��NN-����0�唵����Y���N�x��.��o��J�	�J4AGέH�DҮ%dy�>����0���KVմy�)M2���۶{�e+h�\Uf��kk_ft��rD�[�^p�P*G�I�"�S18�9��a˖4Ӷ~p�����Y�S˻��8yyY�K�	�W����/���<=r�q|�<0�9��Ѥ��H���Q�7l7ѽ��^��'E���:����\���Ǽ@C��̞�A���)�]�Q��. ��8���ӥ��Vx�z��JU�Q�V��ޟc2�!zXXn�[�[�J^�j>3���)�T:'E�=��C�Qc�?145t>�j\5H��l����v��ݴT%7�k_��}*��l#�SG7�IW=J���u�H�Ǘe��jw"�X`