��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX���6��El��&u!O~s�iҎ?��}�Z��0�a�i����#���Q>�y�S���q�O�S��o]�L��atS>���}�t��ɿ�@��<���'�aL�B��׺�/���$U�*����}g���o��$�F�Hy��ѝ8{����ׇ	��W��Ol�1g��q��"v�m�w� ���^�t��30)��m.��,�@MD�{T3���^۷�s�L{�����	�@j rb#ַ��M;?wVGG�>�������]���F~M�;~{�����ս0T�)0*�٪^In������L�s�#�VB ',:����`�eY�l��/nXLI������i'�(�-�+[+�BWDg^i|��C׭�;u�5�r�a��g���K̲���ݢ���1�-+}�=�Z�bM���TA���/I��'��#��f*T�$�O"G|'%�6�>Y��t��E��}��$�&�-w�W|P�B�tp���fh�φT���E rXr{���}>UT����W�*����{N��t0в�tԯ�[�ڃ� 2�	j�m	C���R�6*��Y���G_CD�P<�귏��o6{KP��Ӈr�w�Y1��yY)�g	GŠn8����"4�1�h�rL$xpZakƅ���ˇD̗��ep���N�U}7�x�BD�&	�7\A������@��#�}%G��d���|x���pc�+\�p�/i�H6Y�7����8Q���8�'�۞����`Ohvk�=�ϰ�ߐ1ą{��ߒ���Ԃ�~�0|zfj�xgq%m���3�-�k���#�j�Wg!�ꓴF��cmq��'�xj�x5v6�J�d�~, �z��GK���a_q9
�PT��	$��U�Cf�W8|mΜ�|�H��m�L^�B�ȉk���qi~:U�yp{�V�>��rd�}st��TVj��>S�Z}��?�~��[\m�L�Ahu\	�G��G���R.��%9U@=�S;U���]����� u԰��]��Uu�!�`B)��LVG��i�`�B�~�K�m���47k���R!Q�9��?�@��(�&Sb�n�G( �B��`���A*Q��_1�pBTf�+��AqW&�e�9��',e����<�v;8�:�o4��=��q�a��Ҵ�˳t��(0�&	�
����k�؏�{R�Ё�<�6�x�O�N_�H'�|o��Rʤ?�� �'Ȭ�_��Б�T~o
4.� �}�Z��cHQłׇP���R��f�!g�*�~;�FD�u�QM�_�mE36
�r��!^�A:C��
ߗ�y7 �1l�W�O�=��{A3fe5����`��6����'�h:�vu�#��*���jE������='T{~�����.��4<Cd@�r�JT_ɹ��9�;FhJ���	پJ���O����p�ȯ؆�

E�e���AC�@�9T�Uhd�CZ'���w�:s�^X1d��%K�ݛ�<�K���e�JQ�7�j&�n�"�����B�96��^���dw��HV �=(���#>&�U_��E�,,L{/*(�$ˁZ��V��r}N`����焮̾8�đ7O�kU������	IFc$�j�vD)��T��,y薙BűD5�f��>=Tz_�[YD��9H�xg��O�A��B'JfPf���p<
�<i�/�&��J$
A���G�c��������H����E�&�3��N٤��<w��o-NY	�s}mb�PfH��dw��_�^����wo;RR��q����^qI�e�+@Y^����K'''���os�n!\,8�^��eF�K�8W�Ɍ�G�m��e-<��mb�%��Q��9��'�"�7(ρ��D��lt@T�ކQ
���ekO��m|�}��P��OSg����]�H����댫 .������m���81�O1I��2�K!8��\�9�E���|��	�n��3H�v�z=��Z�!�;!��c�i�C�NJ&2���:Y��p΋���'�J�Q�Z۷D8�˲d\ep|�Fn�7�N�FX�8Z���)�
0G?d�i�ܴ�Pm�o�u;��7��_h|�)��%�Ҟ�\�M�:��ߍD���Rՙ*������ׯ��CR/�����3x�0��x���)` g)�pC��̇]��S��Fa-�Vj������o[e�+.E!]Ʈ�h4�km��)��e~P���ʴ��z\ (11fX��̄�.b< �,~��<��i��ä����Heɯ '<�3R�{�?�{�2q-5��:@�
���$�M,^��+��G�4�?d����FG��@ڎ�zڸQȌ���+���R�sux�Uf��^_�T��+�h���$�>s.q���b:��xMM�1`����EXϒ:G1U�Rk�le�K�����*���9Yh�S�	?\��k�8dǝ�[2�13���v�����e��9ً��{���y�hq�Ø�L: �3w�@eD��o/z ��!h_�*7}=߿U8�H�1kW#�
a���nKeC�J撊|�����r��v��N��u�5���J�'������2��=��҇��_�>X�߭
'^(�%���h8�d���Rq��Y�+[�J�C�p~���	A1���}4ڒ��2L�;룛��X��)V�⹋������E 2���-
oĲ�5�B����)�	� ���h���@�pAF�u����VI�$��Y�Wݩ��v߻��E�ǛR�]�F���B|e<�;�.���Z��TrkG�9/+�A"�"��S;��0�Ϩ�o/yv�R������>Q��6k\H��{.5l�j���Eb����:�*����mDy��YI'�vt�c�N�#o_^^�=���T�r$����������}�nX�o������w��S��3mL{�E�0��bƑ�X�T�d��Fڋ �w+e,�M�Á�#���=R�,���AAC�ԑ��X�~8��㕟�#���[�t�w����9��(���÷��P�73t�.����y�y��jU���6T�'�,��b�zGd�����aj�a~ ����L3�#�T���aM?�vu�nd�x��p�D�.���`��޷grJ�h>f�p#j�y�PFc���)�U�'��T�U{=�pq}ԊU�6I���*T�Z��g

\�7�SW��K�?�W�=#�*��ջG,fҒP�9���S��=�K�#՞%���j""�0 ��z+��qx�Zl�x����sIj<��w��&x���O��6�G�&��'	Q���jQE������|C�#�%P��Ҫ�m�SHa�ʦ�'�QG�A�EY��VM��izx�2����`�蜫�j�R�\)��GH7��	ȗ���|����_`�S��c�BD+�3�R=��*T�Gζ�eߧ����33!��{g�\�	��ɥ`�JG$�0����S��qf��k���b_
��鸯u}�g�iI`F\��o�>�sw��v
ԝ�%�1���Ȑ�=E�t�2���T���I��um�b�ϔT3�Դ�w�'�A���5N��7El���6u+�,@d@}%�m����F^���[{^�F_�C%�_�c���pN-cJr�U�٨%�z�4��2m��L��0K�����~��o@�1+�U�Ŋ$�l>܆���Z3I+���K;��4q�q�/�&��P�0��ӱ�L�
J�R�ɔ�o� �cj�����sS!q@꒐���B'��#��j՘�+-������oo�&jGS��d�Y�'��QEo(����`�����������q�;[�`��ɏ� }�
-�eRh"8�H~ǿ>�����vVi#�7�$UíT���wÛv_�6�V;ѰqT�`�}���C����2`��pC�m�ȼhKM�!E���A}���S{,���Xo�_��$�j�[zU�q��bTۍ7��������Ȉ�����o�謉\w�NB��J���L$���Q�����a�w��P.N�/@�Et~�WA��g�].'��-��$�6��7==-��)L��1�A0u���$��������Y�B�VZ���!Mfx�.�B���
�t��µ�-KrT7M��s��wフxE��k0M[�L 
c[� +����f�m�Q��wI�9]��rb4��&Xٮ���G �L�?���(�u�77q#L���p�z��r:�����nޓ�z�W"{�;��E���	\L@kt�M�)�7�BKy<�c6��F�N���&�o+�K�H6��k���F�����l��
]��@p���D���q5�>9H�]�ݞ�(HF����F�h��c����ǉW�M� ����U�e_�������6����{6�Y=�� �*&�~\���}���eJ}6�6�#��D�����IPD�v�`0�qyQ�����.J>M�/|�@�ү�
�¡����B�{�n �RP(=d��z�S��� �jOWB��g1��V7��.^ý��-�*�0���Ys��Q`?��x>��Z���1T�]�՟2
*�2�$���B�~n��=M��6�2�,�Ƽ�!��}�,�_�ޛ)I���������V��x[1X�TL��>"On�l�`�olЌ�οL_d����Z��ۣ�@�8LJ�jY�VGs�7�]PNi]M�T)���4r��S���������H�a`w����W��U�����"�[g!e=�K���c��^�`�?�*�:đ�>�y+�CY�L2�-h�s�*.�#�Igj8}B��8�g���AgcH����~��+c��c�}�9@�o�z�����������e~�K���ϡ�A�u����DT��T�!�7ͨp6���g��x���e�Z~�9�R�\�MF��C�n�.�{4ե��eRo6�b�qw�����Yb��)�.c��i��N��C�^���YA�^g�)m-	&�^yצ:WFF�G���j�hwf���������Wj�/h)⚞�������AK��J"8Z҈Q��noI�v���;���Dګ>8��9s]!�UFr]��C�:��*�l��mi784G�Q���;�5�a�m�w�ZG��y���+�򊷠�[-!.R�=y��U��:
39���_�2g��MN8�����c1�'ʔ�B�\�1��Z�^�M]\D��t�!_:�"�_�Ǯ�ߩ�G��S5X�"�n�3~X�(�aק�&<�C�l��¶ &f�95Tf��T������B(��ձ?VJ�6��u1�o �-ьYi1.iU�����A ��{xjRw�nE9�JFe+�셩�J�c,�������G�����N��I�����R�zs&�CZKI��y�Y�)�*�PL����J�d@w�T)�*��\`ƬkdMØ���Kx�q��UU_ò@�0$}�罅����ä�:���"�Z]f��x6����uc��U�F4�F5!`,�sE��p5k�L)�E�Ga�|���C�z����>)��£�e\˽,��aw'�R<��p�h�~�����	e��U^R����La�G��fDk��BxׅFga�h%e��~��E�52�K$p�G�a��qU��l��]{���tK����|k�,�RN�gn��t���;���Ԓ.��rN���G>wf8��qʮڃ8,��>P�8����xa;����Uee�N�(�t�����}�jB�)�Ŗ�!�q�r�h�{��>�{��z�����y�xڴ����P��~}���`���0w*�EOo_mi�r�Z0��3|(��Z��S^^�����_}� ~1OǴN��8����)uЩ2Bj����1����'J�{�8�G 3�oi:߆E]��&ԙ�`��.���2�l�cđ���d�e6�k���=�*��)���b�(�O�a�ͭMwX�8�09^xa����Z��S�4*���|�y=o|�-��Y�Lܲ�r�k؄T<��Φ=cH��?r���M���C��Q��T��b�'��N�-l:��I�asEɪ�*;U��<�I�u)Gr�����{�?�%as����ֲ��<�H�/:(�;��{�g�1<�$nW���}�\ʚ�d3�P#����u`��iD�e���X�brk������	(�Җ8���4�t:��\���K(|�zM�pا,ze��7��G�f���������ǜ�4O��6��i��"7?��b�j�����r$�q�ޢ�7v@us:q��䅪�z�V����|��)�A�������@���f�$^���,��G��)?�.J���۬G�z�x`G��u�͂����d��es�8�On����N����6�6'i���42�f�������<��8%�,E���~JL>c�T����?ނ����ٝ$�/>B�uV��*�G�V����~��-̳�:w)��$5��3
�L�k���!�1~�Q� �gr��&�΀-|�ǃ�Q�ͮ���^�߹�:�T�5 �c�)p�;
bs�0:��-.�-Rk���V�Ty=�)l����/�#^�lP�	���ȍ��i/]��7�����lL8ܝ�ÁH�NDPi[1�1X,�#@+�s:������ �H7��*���Kİy�k�Ջi<�s,A��ł	��$-�-�_0G�覆2�rT�v��H�\8�9Fߒ ��՞��,]^>_	��|��g�뫅G���	�`����,��R��`���>���M&�U�u�o,eI�2E�3$�'�pQ��-�V~q;A�aeG?�(�WJ/0�,�(p+ޱ��F5U��D6��-;��7����9T�~�����Œ� (p��m�@5ܟ�WO�L�px�����  q���0�4x���/����g�(�yWn��d'��Anң�ndc	�e}8�eE�6u��G{=�?��y��n���	Ʌ�Ab.�ȥ�^4J,�z�
G����ȫYq����q��'��>
�NB����f2�ؓ�{��*�s�̀��n8��?9��`��ivl
�;��Q��'��P�
㍬�+m���I�i�Lb|\��K�Qq��D�>F��Z��Z6�|��70��r��{A�<ݷJ����ZԢ��(H����S8���r�)OgnN������y�cFȺ�i3�-E� �Gd�o,���am��UT�&[wa�����5ǕH�U�b��ߏ��I߀���V����L�t�9ң�}Nh=�6��a	��فO}�p3������-����[��%"<��;��,���[�f��r<���;_/��^���{pCK�sh�!�A�%H��`���>6\0��D��R������9� �p�&|FW�Po-\�����C�_�jf�u\�����8�ڦ�r�~�Z�D�Li�7��Gl���K��O~�|,���ΤvIA�<��P�#q���L��"�at=�wy������1a�Uni��9�5C�)CXw�xKg��MZ�zmoV.���U|�jx�a^aH�^�}��{L�C��}p�
�>O���Q���L�sA��?���xo|�徚���ϑ%�!�l��0��fF�d�sݷ��`�.�G��ѫQ�U
�ӈL)�!�@�����1��� ��=5Z!�.N�m�+�y�Ҳ�2��<ǚ:E�����BAj�}L��2ز������a9`�% �1�y��m����7÷�a֨u��<�V��9�F�:��8нe䁲�1�E\z+�Y�^�tG��W�z��R���|gU,�+��z����*����O7���;4现%P����B|z���[9�.'pm�?����L�j�X�#�2��T����{�
m�[�t��LH��ۗ��8vFQ9�����̴H#v~��/�E�g��-�ަ�}�K����LɤA���*l|�v=��' ���_l?�E Ƒ�c�8��q�8��>d�%�ms���%K�s��p���a�
n:[���A�P$NGUW~�O �����l$�w��K܆֔�v�*�Gj�i���Xyw������Fw
��6s�����n�����U_���Qi��s$�d��UI�J�;r��	����(}�����@��wTk\�Pk�c��2�9O*������TA�eC��N=�n�R\_h1+��M�R��:X���G=�䛌�����
	����F���gY����n8����tBmR��������Cv����=�8j��ck�iD#Eln�o'ک�BT/��F�_���}�6 �ZH�ڻ������*�Ћ���SEq�OVӐ�X�:~�o�R�W��2��~����Z��`y���r��y�5�M����tr5�]
�}�S�Ǹ晜]0���,��ϴ�*���I�J{;2Ԕ|�.<%:]$����&�	�(�(���_)lɴ�G������&O�.��?Wm*�-���1VE�����(�;"�k*�=E�\ƻ�ϔ��9�J�7[��n&e�:�p?��D
0����`(����i:>`��IL�[�Z�O��v4ڪ����=?y���w��:���X�}ࠣ�����c�k��X��H�i��u-�}���+��D��%|�[�9���q'�Yjg7�T�%��bDJ�m.�����3q�P�ٕw�Z@ip�*\�H�^����{|�a�:fkב&D
�,fM�����F�c.�V�X�}��T�谟��i,SRv����o�����
�zW�ĵ�M �XVrE�4CU��]�}_"�t���������w���*Bv���fx��z>�=�}^^UTqXӘãe��ՍKP�1��Lj�X�ӳ�WqYH[�[�c�h`[s�Bn��Ѡ����=��c��`����
��?�ֹG�n7[-���_��t���v�S瞔'�����e*�Pv��a��W�t��