��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��>��/�є�|�5.ƚ=���פ��[J��3�-l}�1��ۈ�C̡sF,�Y?N����'�mL�����́SiPq��6��(��|�+�����_�o����\;�^1E����~é��r�}8�
ÿ<҂�Q/�U𢌾�՛]���>�)8�R� '�4��vV�mg�X�>�v�J��qc�MN��O��e���I��P�uD�6.�T��7�9�	�v��f
�^�;�����X�ៅrSl���łV,0vkI~9
�m�xͯ[�|\��|Eր:2����g!z�S���5O��T�R~���կ6D9C	h��
�6`D�Cح�7�^ê��F�$T�evI�\���t����'4h��&#��wj�&?�&�Y�{g�Te��+�	O;k�p�`�[*��J	���$�~�9I�����e.�AP�6�P:Iv@�7��ǀ�l� �j=��L:� �Z	t�B��#�6Cp�q?��@��AS�m���c���O3�?�T��B>|��~	���e�C��?�$�/�����HZE����<jD��^Ic�q��p��	�:���U�:�?�wv��	r�˹��[#���؋�?�0-�bǽ��Vȹ�2��6��m��>�P��� ���T��a�Q��*������W�4�>TH��.�dv�羚���zZ.&�w�������W��|�%E���|2�,J���B��T�\�t����܂����SE�<(�q�������<��Ö^�	y�o��ӇU�Gf�Eȵ�g���E��rDD�iW�F���m]-dw��zKg�L�,X[銂&:��h�?D$�]Ǡns��h�x�ky2��~�A���ח�^0��?�V���G�?B�$��a�t9����V�H	C����QVq�	�+1�@͵��4��#�
��X��HA㌮e�b��Z���*�d4v���+l�7%O.y�j�r����S�c����'��Pą_��g���! 3��̀����4�4�T׸b3�Ir�ܴ��K�z�2�9�9�&����j�8o���t������gE3�@"u�{N}%+��p[��1��c��ȉz)�z(��t�l��k2�.��;��Ďc�'{�O-Co�4�p��0-R��s����� W:ul;�nX���=�-�M�e�S���mM��]�0bs�M�γ�"� R"[?'��Lx��3z=N�-/���*�v��WD9Z'�m��w$��;h�d�|��3AlJ�S�Uu���4�ٹ�b*��`q��$�ݬ�v�U�����4_��e��+)s�
ш(�u�J$&n���vS��z~OL�x�c	�������Ƽ�&^{w1_��nR��C�~ %�k+i�B6Ǟ�U�^Y�|�l}jBr��;�(ix�g�R&���b���Tt�i�K]�;(fL���q�u_�֛{����zD��7��y_}\k�9�P�߀�S٤���k6��<�JUo�5�d�9�c��H�M`Ywx���1�*��/>��*G���N�7ԇn�h���
D����!<9ܞ�1UsF�ղ�Y�Ll(7��{�'����ʊ�۶
]Θ7%��~�̊K!fcu��6Ǳeu!�o��ϸ׈�'��E�_�T���7|&����/+�.��pS'���xg��h����d��r#���'�A�誜j��"��%[@-_�)/0������~���Y��zyš3֒^v��	^��k,`ru��rC�J�_�<��A��*�gŅ��u B�$��F�S{�*��`[�m.�t��m@Q!EcQ�y1�쟘�I�cy'hµ�5WN�h�-���%���\P�fj��, �4�,�7��;Ks���5��^�͠%ݓ)�n9q �c�����_���F���݃`�%�z.�+G!���"~�*\޳��8h|�x	5�� tB��@��+!�X����5�8��1����-l��Tp�b�C}��q�](� Z-8K�g$�|�Z0�a�1��A�FbX�B#��@�Ѝ��=��-}l:�_���;1�����6F��7h�/�r�%L���'�ϥh�I�kc6B����X��>NJ�J��c64S��t��4�n�^�$C��%*|�Y��}w���ص~�f]��R��v��7��x�9����/lh���5��4]m�}uW�Y�63�����)e�މ��>�m�A���9j6@)��˙�9v��SD�B�fn�Z�*�t�`o���4�:k��6�O#V�̭�
sh��䍠��p ��$���GUEy��R��5�DSQ��!���P���_q/�s�����-�d��Z7ΑGU�d������
�ݫW�����ИѺ��f����iX<ϏA�u����D��'�tX�-y'�oX^����V)�<���u$��'��[}�`���ž�b�������_��� zL���=^�y-�s4͈')��+�S:CSa��%����N�eyZ�$�E���*� ����D�а7��0Un,��]�|��G�7@HG��KѱKB�{�X4	���	*v�⟑�t���t�FY�5	Ht�j��SO9�D�TӇ=��b����\g�r������*�ܬ�U�8꓇�����S��v���S^�[�u�Ot�9$O���
�`��t�;����K�5 ���=hH]!��(�N���V~�����H?!� "��,d��._ $#PJ\jv���b��M�3�.~�G��Ni,kͪ;1?V�}���'|3Eid�p�Q�f�L����Z�E1�z���~���m�b�mVmʮ��I:�=O��n\V��N�A��T�O��i��� ����#N��I��]�f�ق-oS���F��J���U�̀�{em;�9󠣲�Ph�F�Ph�^�.�v��H:�S�.W��,c�<[~�H��Ͳ
����Gw�n���e�`[��z�Z��,0���x� G�=H�ť�qb16��>�vs׶�YU�������(�s�#���d�r��]�s�^o��1�
�V�/�ݍ����ɞ�7�MD&��'��	%'��<�4*���P�d��!R_j\���:�xS����m<̘��?�zװ��k���-3���[��Y@�3D1�S7`��q�(��A/��l(����nT������[HaK8C�c���[�l
�����-zgp�9�W֛Ș����J�ǩF�W��_�M�A�F���q׋�L�N�p���mɬWfY��YuO�h�D�w]C�~v�燛��d[EY��s9��@K��F�;;�Q
�I]���Hɡ���S�7p-�p��'�ئ/���/���y�����E�-�Љ��!�X�I���e�<JH�(O��+�$� TC�����l6X��D�0L�5�Q��x)�-���?���0���*P� �<A��H�jH�}ʌ,��ҩ�&���� W��7�����e�GL�@AAdN�t���8>��3ȣ*#��'��*U�Xx9��u�&'eEz��HI���Ԩ�Чw�EO�}���w�Yr7��~��MB�ӻ�6[�)g4���d�Ǳzq%.@���Y�}��x��mگ�ڌ�RE���<>x�24����BD ��{A��������m�U}�'-��n�)���p�7c�W�t5D*/�Ht�`S���r�U�h<���Xo��$�XW88�RB/!�.f�7��NqX!���8f�@�(<l�c>��m^Hra����K+���R<7��0�iT/��QI1��5����	Z���ip�t���W��f�L��K4���Fh�����z���&t?�x�1��\dO�U��O+�C3q�2��Un5J�e��7j
�)s�@��9�{�W�NcP�W��?0��پn��g�FC���V�8��灘�+Y�^��:y���ȭ����L�ɩ0��6�]q��*T�P�\-�ڟn���.3�����o6�����S/�V���B��Q���Y��=�������py�&��6��Y�z���r��4p
E��Ѯ���G��r�*]Yd�)N�R�f�N�r��w��de��^��`0�L�������<߉'�~Eդ�v�3뉸�H���ê<��������p~���e�n�n��v�݊������H:��Tt�$�M,ct@]1�A]y3�C�Bq(���jTG_�R����_���ʀ�][��~�VA���{�98%F<�.D��d^��Ы>�(F���e���HY%z �q�S�F��o��I{}�<�Q?DhT��>��p��P�`�@�V�IbT���i��덛ͦ��N*���g6-� ��;Fc�	����ȟl8(+�P�x��R�Uq�A����T� �V;\K=w9��.��DN��1:�}�pR��E������1	�����	i����gUR�.�'}H�r�?C"z�N8�$��{�!��[�b�.Za�mo��7M��#,24	 �?,'tg�7�@�����&��8�_OR���O�?�%�a=;�X��[�)�EM��nQF#��w��&�}Ib)���=�嫳����&���p�����:�.а��s'��/n�CD2_ܧdiҪʳ1����[=o�ү!s�������!�*cȵ�o����32�r�����(�,�CVN+a@��a��]k���է�L�PJ\�&s7��CTlҷ;(�85�;>���9B�d�G��.��V�
�f���b��#�D��8�(z��Oώ����g��|���W��ܨ�qָ� �m��٣b-8iLގ&��2Ql��Ȝ�Q��Md=�#H��#LK!�Y&��.2��W4%�݄1B.2���5��Hu�5�Qaf$-�v"ht���aW��0(e#}Pv��n�����M�b�W�^?p�E�b"§�����-�ҏV�\Q�_�藼�Uj���+���Od��Tiڨ�Z5C*q������`�D_�<„"�l��D���̓�d:c�������4��h]^�a�J�#��)�D����Nϐ}t�/=��T"6�j�v���o6�<
�ě���4�� |Z�?�"	���<4�G���-��s��<���;�u�X���s2�(��PT�|��u�⁬k�K�dS87�LN�Eg	���u6bN+ �1i�$��ϊL1Ⱥ?����}�O�yY��L�3��4�`�)��\��_
�:u,�ŚFM$�:XQ0��g�b)	��� �\��҅(�ZS[�f�"����R�P˵ER�fq��Y�1'C��q�,@��i����&�mjlo`��␲�7�I�e�M�۶��dw8^I��a�k(�*m[���Xg����!?�FSR^��~�p ��������crlzH��WE��41�%���gm�ʴ��,�:S�yгY���t>�uc��K���ͣ5X��KA��_2��ȫp^��㋔��~,�4�����"s�'���!��S�*z�ʐ�v?	�J&)hw�ʈ�lB�SX���t��[�̏������LC=f!D8Q�"�[Π0(	�n	E}j,�[4z�ւ9+���V��x���,҉R볾���$���>�n������-U�	��%K���D��p��~pz��u�m�&�/]�*�=䦧Q_	����2�6;�c�5W1v:�n�їB� ���p�pH�|X�C�_U�j�q�}��r��Ęb��(�[~�^�{���P�Vߍ�bg�X��ı©W�d�O��{FGK�=ߏ���Fğa��J$A���$�e����Cv���F[�7l�+'�����P��ϧi
H�<����gaZ�ob�S�OJi0�g��-[��@��~����ޡ���C�׶xc����qx#,�Rh׊�p|?<3VM�lB��2�,p��3��n�Yl(� ZP6 eJ�Ӗ�i��+�	 {/�e	�81E��,칎����=/T���޵�߂"�s�'5\ 4��"���C�烤�k��A'~�Y���� U�)(�����H���;��mh�'�"6�(. �d�[�����պ��öV�|3�(��bמ�>���a�ȑ���˖�a�l��t�S�O ��E�N?x��f��*�M������N�`%"�=��΄�E�
Bb�ʀL��W�1n�yY���E�4J�L酨�O�L1��SY����	y_����s��1�?*��w�w�щ�G�_%�[�n���Z�e�n'| c�M���RSB<S�N����oPM�7`��j�X<���.\��Ct����C�}��4�`԰3��v�_3�2�Nc`'�w�����$9��P�������Ӓ��
���T3��}������y�(^#��=l��E�P��ly{*;����O���ІWi��_�C�C�j郠��w���������7O���~�����e�������&��'k���G{���$q廤v��j����O'
�)�Q
�H����g�:Q��o�;�m' ��z�Q<��d�i���#��~ӟGQg�a ����Vg1���wD�шtK�J�?�Q3x�x�h%&l��9��K�M'���wU=������G�b?�����b%��=�M����GHao[�Gj���՞���,Gᰥ��ؾ�4�.)�ٵ"�ʬeaSG��zf�S��:��ӕ�6%�#mce��
a�O(wd@T�P�^�Qm�Vx{>�EB�e�(ˢ�nT�\������Ɍ��x�R��o]Z�U�-��jr!�^j���V�%ޏ/nb�տ�>�������� ��)A���vet?�o�q�H���6i��I:×H�2�hJus�73��M�)�̱�_��^|&��h>-��d3��@�0@�Y��ӡ���(�/Ϗ���[�x0�x�N2�
��ɘ�T=8y-�sq��Q{��9��<��O:eF��?�/�I�µNIT �0>���d��%=3���y8��s��ب���c6z� ��?�sȥi���a}%p+�ü {�k���� a�Ŷ�ԛM]r�b9���3�ӛf+hmן�y��J��=�>�/<B���M�MP|�0�ui��r*�T��'���i��c�<��F)6���łL��V�����ĉ�Ɏ���n�e��!C�ݏ���dj9a�>�6�T��B<��N	꒽:�]$r�1�bd[˩7�ߥytG�]9�1�����a=%y�k��F7z�Uv[@����G�,�E�EO���
~Sؐ����	���G��>�,R]�I���tHK�s_�ib]��kd�����Y^�¨��Ht�I�q�Զd�mT:�p��Z}4�hiw[�}��	/����#1���c�o����9-R��M�حxԥ�^�-7hk$��%�L�Q��l��߮�u	^�z���������o���6�f�#�+UdtG$�R�:�L4q`uX��qa��=���D��[�~��U�\�$��ةJRwPV�.!��">]�7(N"��t��;A#��C�D�����=��ÙT)�&��i�%��re��iu�\T�w�vp�0߅f�p���0��9���r���pU��$i	vؙX�zq��#[��rZ��I��+�B�>An�uQ��cac�-U����v؋�}��Q������On>�Kjl�b�=��<N�l����� ��&�S�������D!:���A�k0(���fw�B�}@ϔ��:���(�	��du�]����T� "��Û�#����w���)�w�����"��˕����I_eu�I0�8C�M��Y�D�fa� �#Α=�2
.]o��o�5M�����y ���}�tN	�`^s	�0;?v��~k嶻�jZ����r�K�d�����n"n��٠�=�}ˉ�Ty88l��g�_�<#\&&B�Vq��5
��|�X��u��Ε���iK"!2z���?z{DN�%)�8*8��O���^N͡��-���Ӊ���K�G�|,�a¯�K�����}k1�̟���a���0o��8b~�׈G�>�^�����8�Pl뿵���eepW��a"�y�A�k�Z/yo�|�W�*�kw�ݞj�,��0-�y��Nf��oQh���Ar�DU�>{�0��TƷd
ĕ��Z#&���e΁�8r�F������ڭޢW����k�� ���j#�M�l%��n�x<�_>)I!�֤�Jh9	#����`��F@E>t�E�9!�~̞c���k�q���muF(Ú� ��(Gv�m���ek�å�[;��I���p =R���{�_�o6�_�B� �k튴^f�:��*;�o�>��i���F#�,�n��[5:���cf�I�>"[�m������0綰��Ŝ�W�5g������$O���%�1�qҵm��\�$A�%���0�S��:���A'�����
�%�Q� c�żm@b��qsR-e�{���� �^�_3P�Z��n�a��3�'g��dUy0xT �Uq��|2Ipԩ(m��7�}��aup�F1;G����Lx��(@nYt����d��/�6���dZ}";��֧�*mh�%4��6��N1h[^��rԡ���� �S�=�H��h�9&r$h±O�}@}v��	��M�������h "z��[��ܵJ/z ��_Ly�x�{� .=˷ԓ<�/Q�fH�U p�^��sð����^g�2>p�A�4�7U���L��=�G�^����x^����ᆽN�9-�!�}I_eb)�G��~)/�/+���QMW��o=��_�f`��a�agݧ"��� 
���=�cv��ҏ�V�,'��atF��O�h �����9��J�<$~��W���z�3o�賽xH��WK���� 3��Ũ�揀;���7p��V�b)z;�J���"��L���Ӧy��&9����?�cmx1!`�t.��+=�X�QܽQ�/Y`���{��v�Ad((�� ����܂��M$P�Fi�=�--6���Eh6��`�����7��Ww�T�t��X����մ���gV��/<�JJ=}>Mdi��^[��n`�ʩ��g\xj��,S��q��|��销��;Xg$�`eVr]ί��6�*��z�Ŝ+���5o��