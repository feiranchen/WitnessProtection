��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�ƶ�biA�#��m}@�%y4*����'�  �2��e�{�E�q�L~����j~�uR��I��9P=����>?�̦h�Өs�M�|��|���<�����#�h��O:��c"K0�5uO���@�G`��jl�VM�ﵧ�]�ĕ�	�j��❦c�/$���J�! ����!�º�\�gh�4�r�̊��w潊ß�c'��ޣn]������^k�\�9�IS� ����F�΂uЬe��1W���WCl���|�!�!8�(L��١��m�[�N���>b�t�i�@wX+?ad3̌ex^����lW0��B�j�_��p7����9��R�8/MoteͲ��`>�<VԞL��NK�� �t�M`�^�+�6�P9�*A�3@Ir�~�Q�g[�Q�þK, u3��(�f�$�x��?J+#[fW��Nf{�̶e�U�*�S匝�w�&� 泧����_hA���������"�v�!�d�3M̘��t`����}�����A�}_]mF���R��
g�X�븪� �2��9��l	+ӕ>ܗQG8�K�E�}c3PUK�Q�[�#L�wo���f[G��i�|����ל�L�{�>D��z��x^�w>kx	��;�7/�6z.pE9��-�M?~��;���W�]4:Q��ї`�ഏo���H۔�/S�Mb{�n�Oq�Qc:�����j�s�?Q:�C���8�XJ�����n�~st��/�+G��)a&tN�Sv��g��c���Y=�R���l�1�C�c�,��
����h��\�)`z?�\@&��2��j�\R����Ӷf�����s����,�\'��0�f�Y|J+�)?���w���K�����'Wn���oL�L(" 2����J0}dF�**~�!�����aF�P���ߡ�;�R�o�
��+=(�<`�;-f�V�<��Q���hL��Ş��^E*�*���8����_K��H`���t�V��r[�C�Y�d��c��-_�`�3P��xJ�:�\�q}�4P���؈���%�O��U��݅ 3��+�Bhe�H�ޚ�Ø���]!�a�8@��N"F�������zf= '��e5.[�v�������nQ�Ͻh�?=��ñ�^���� Ĺ��K�Zf��N��NZ��!sS�b�d�ֵ������p#�T���m��s(�q�	��r�=BA	��t6|9�8 �U�T�u����WL��/{����G�K�����$�n��w��~L��<�k�����g 5 ��ܩ�2�C�������L_�;��b�;WQI�eTD}(d´�J��ư����3�)����&8�+��tjHz�}\:��i���O:fYM�_ﻮ��N5�ѩ��l��q/�����OT3���lfO��l���g���w����n}���4
PW���y�S� �,�P��'�Ssn��SU��)�h��u��Xu��������]��[H�M'b\�1�yLe�|ze�Eu���')V�*��8��g��r���@{)�5����U,��k�׆?��(�YxY�B<1>"מ9�%m7�*��~WV����|'�Op��]�a�TD��*�F�7�	�9u�	�t���W�Ex�)��lt.�5�
:��S��5�Eu<�scw���5	�1�b�<������Qd���HL��LT�[n�p��ÛPd���N�$ɺhz�ü����s l�����cg+��
��� $�n���� �����wZ���"4�\�����PQO����
b'5�̠~�[f���6�!��W�xL�kP�ϱ��b��
er��*@����	r��*gGCY5�/�;��_��?�-D�y�4����/�!^�{Ufń�g���q�$��o��5CW��3L6N���*��!nI֎/�#�)���&��SZ;�4���mH0.�߲.^|��[]*��[h�E��OP����*Gp��{zrx�}!1e�S=���'ȌߒJ�w�<\�_YfgG�vP
`N򖨧z��x��]S� �^����o�K�EL��aU �F ��3��	�}�����Qw��:.�C#:� i4L�`,[#0K����Qh�l�+2Ql����b�&���y^
L�����g���M�)7��su&��C�g�;*��*�x�qu�$�W�N�#tw� aiS�nV�����2�AC��Bg��`Q���=7u���pVm���h%W��(�qz�칪I];�Љh�#,��6Qh��o��U�IJ>�����ɕ�چ���>�R��m�$�?ǧK���,t���`I��P��^�)𾌉��}� p�Gv���R�w�̞u��|��F���e�]p2C~���Y=�-�r�q�c� �;.��j�Pg�#���Nf���;�]�Q�W����uvRKg2B�,�߾�S^z�¼����[?6��2^�O�4 ����@������ �@�(��4=��٩�Q�)��#7Z�d���B�χj*j�!��&+>���0������ ��> B��	�@:]���W�w�敛�U���V/�B�9�iSM(~��-�u�=7��Эh+�r�wu֍�iO;�@���	��M�_GE���*?�u=�/2����@���˲<�TO~��{ur��Q�Ӡ��$�Tį�5)0���-��j�0ber-]���(�!N�P�O�8x ��~A��Ӗ>Q�b��J�4���4Ik��Aǩ��C��<(������`�R�V6'u�	(Y%�d�0}�*"	�
�=�R���t� y۶�дT2� i]��%Ga�lwW�_׼�������+F`��Λ��WR��'��>Ѥ��z���B�5X͙9>�FČ�5,�I��R�{�).&s�7�'4�2�*3
날]0�'ꛇf٠~*b��_$_|�輙���L�PӬˏto2w��)����~��"CSl�=��,u1�
�����Kh�2�(vkL��e ���0_��_J#��TC��гu+$�Y��B��uBY�gfk�a|��"�;���0G��&b]qq����Z��	�#k�B`g��6�P�R"��ZlK�f�]{�2���%�#(r'D"��b$�C5�p,�i�i�&� �+�.;i1Pː�X'ҍl6~�f�|�=f�c�Cq]�ZD��!<���4���&tH���������w��g��$�ړLWS��c�3id�	Z5�C��{���V%O�x>
�?�%f�(�Y�	�v���=	�6�}�8>̿8� ��������XuR5�J����z�,}��\-ڛ�\�b���q�q?��A���ǜ�=��mT��yG��"V��U>@��u����^������J�MgZ�g4>7B�����z�'1:5yH��
x~�S������g��-BwC;�@R���&����r1����A���~H�Cf"���1���n���T|�4Ȓ��-'#2㷧`��	�Z�-�H)���l}?��������䪢�����Qfڐ�?	�e��R�h��Q�\<���U턚a!C'&�x6�"hg߷�?X��W��/@V@�O$�wbO��n=�xoٳ���׺��TY�fL��p��OH	�h>�7M8�ϲ?�B����Y����1�7��@r4�E�8@���� ��I��Q_��D
a@k����P�1��
�,�ѧR�Lճ>31���՚bG��1��^�i�S.^~/T����㛕:��k�쀶���3f�L��Y�0F��e�X)�(zEƻ��
5�EHp�嚑�sbƑ��
��x\:L��Ү�pn*P�oc���ת[f�azzJs�",>�"���u�4և@�(-��_�'��K�6��uK^N�E���PY���;��tx�����v>u�pZ�cz�򔢚%�%��a�ٶ��s�S��!�fB���w:�s��\)fi�K�b�X4���@���F ��"���>aoi#=�x7��Ҹ���B �!V<���Vr�|Is��sr^�o������bf��DT��P�h��Aa1������FT�ˑ�­d�Y	��$��]���-�\��gj��1-��J����bYg`#D]ЅIE5 S��4���D?8�A��=7�}
j�f6O���<��]Ӿ���r\��4��L� �c} +2��'E��#�΍5x�D�Y2���Z��#��<h�l�YRVL�=��(JOi��sX4��*勭ա�0y���[	���eX��'e~��Q3K���!�ˑ����lW/��Ϥ���l{~H4�ױ����vV�)4]9�:MP����;��;Az�׍�Rx�61y��F�<�
�����9��ߠ"�y\/�(H�\�=Vrr�t9A@S��q�+��qܠ)��&|��)�i�nL�-�"���+(�'�;O/a3�5ll��e�{��W2m8�#�j0���v���W�@� g�j���^nb�ϕlHW���=����2|�7�a�u�a�ky����<A�K>N~l�}x�΍˕���@J�<������'9�Q�WH���E�Vѳ��L���>�	��pN(3y�E��qR�k_�	d+����1��
�ɍ �A�e����'9�3�=�W�ji�P���F�ӓ7�ŭ
<����=�y3MT�.�5$��;��,��t����hՖN�۷8SW3#�pf� ܄����^����f����SH�$���2�D�Տ|�;�hNZ������̮<]}v�$�h�B ���Kz��n�!� 7��2d���K�`��#��@�����ފ�Թ0ʼ;6\���t��U�Gh�=����U�5x�jZ����x*C�?�(�u�t`�$���I�����p�=���_��2��m�&>#�ˆ�bFJ�Q[+���p�=�<�8��g0Y�����``�E��=�\n�	#�3��Nҥ��5�6�@�ڇ.������K�)Q!A�q�E�ewۯ�BK�m��"W�]<��fs���oH��q�=t�GE�b�k�rF��S�!��^^-$3��µPdˢ"�#�}�|�ЍZ+?�#�<�u��K	���\
��m���������l'~�E4��2��)��Γ��b���g?��5�L�">+�K�
��ݒ?m߰{�I�p�����4��ŵ��$�tB[�El��é~�m��fB���4O��fX�aI[���
��lH��f&�+o�E��]�.{�p@�n����Rv�HAJ�0�>� �4�lr+�ӿ�,��O%
O��@���෴?��>�;7K�1l�gCM1�8	ժ�e��քi�N��,�
hx��+X�!sN&���4�b�7���0�%'�}mW�:����A��%MKR����~�v�m���{!�����V�<������m&��'��f �);��I��(ܩ���c�i�N#�eYEPݗ��
YJ��]��I�UvwG�U���[��)����a辎��L�	������RŊn�R��e���#��tW�O�QO��=�Q\����Ө�U�?գ���I�c���S{�j�AT̵F�|s��r�X������a��S��5I�C�n�a8��4�4`j�$��#b�5�>�s��u�{�����ln��R�6��rwf� �D�wDdp����a�� �vF�N��]0��ƙ�`b[�A��Y6NY��0r��gob1�;��-u������Π��B}}�+�%������(A�����b�j�q�� N� &y�H�VeWdcwѣ	 [���3���{�]����u"N����;8��u��,�l��,جn/��u?.��zI
���L��S��k�IRI����M�%q�/�Z�q��NHU%V��	�SXGغ���	 ҷpR�I��Z9"�mvϏ�N���n{�TR�(��� 9D���zڗȰ�kg�����J��(�#�TV�$�V�Ý��/D���Y/n���(�/����轓/;t3��/�B˰��p���O�fn�R�#_��ڶ4��Vv9_u��>}�A�����~�@�BT�^x�䷻��_���h2�~m�3����i��7�=�B{��9��֏=-D�����A�U ��h��=ܔ��#�'��N�8�KUg�F�@f��Q�c��T�!~b�5��S)��A���ҭ(�"Ȅ���h��}p
z@��*�j���f�G���&�^��̸(q2�]'p�}|���� �{�^�6AP1�&3���V��+���z=���i�/�YF��,-��P��c�Y2e%�h�)x�Y//�����۔cc���ăn���; zhB��nJ��#*��	�s�7�?4[v�.��b���[�HȎZ�n޴I���l����K�gV�H�����XQ[]����_Ng�Zؔ5轿Ė)�B�L$5�u4m���)�s�v.����?P�=a��Wp�˳����
|��h9
#:�SB�l4 �;��j��40mYÂ-�+
�PG�W8i~v��'�����y�b�gyx��:�	��(�"�5At�}�~�"�"㆚�#GkC/�w��A��`1X�OQpr��fC���C��,���G��_ ��R�qo_f�?�-�L㋞mP�w�NJΩk��$��0�	�h���*~B�LE{K����Q�;6*�f�1���Ƭ2����9q^��#g�z��8� ��������c��M5��о�!?C��nriwQg�������K2�ޣ���k�4�=��uF����R���,�X�T���Y$��*�qg3�0�c�Y>�����w�齭G�k�v�&ҏ41�^�O:�y�x�'����(�.�
V��"�ŭ����p� ��q!����ڽm�Y�o��A@%fj�^aW摒����l�0���5=U+���߷+�Cb�\�z#��]�B3��������m�ɊY�e��ӡ|+�L���u2���
T�r�>)h�����a�a���h�R~EZ���Ϻұ35I�QK��L(K�gfW�&�򈸣X����KK��j�yv��x����#C�h���W�b�P�&��ő:\�IE����$��E�8XN�I�U�z�_z��m���M#����ٸbtiو3m�a%�1�pHϸr.&gօ;�"#�d�e�[��M���y��:�"o ��ಆ��R9w"�"7����@�u�F@���+N�3kM,V����@ rY]U��N� ���܆
�S�^���U0+�FSx���o|�QJ�@������Z҂S�CQ��(�TJ٤���((���7�@g/<F��%.�O��
��23la"��\	��R<NO��O�UK`be�9J$�@/�AQ��yI�	���������b�dS]��*�����:o@�mv�Mfx,V����N�2�A�4BzoO[$�zLQ��t��� ��MU��2�'"r��:��ss*�M�������;HP|�Mt���C��Wfڙ��ښ�d�E���b��p	�Ĩ]�Ȅ\Js�_M�����>i�N+QK���bډ���R* �g;��Л ����	�01�A)C�stĊa��?���d���%�>�ֺ,���9� ޽"�p�HGժ��.���:O��_	�>�M"�Z%	w���t���`�,7O.ښ��㩚/���vH�;,ϙ��4
���J�c��(Ԃ����#�;�g/kl9�!�~���k��b�7c��o����>Ђ�X�7s0�	 @a�5Õ�]�}�m�VbOA�E?��T)����9w-ߤ�5�4]a�lUX�Vx���r����#��+R���#nJ�ps��E��A�6l�u�:�Q��s)�iiz�9S�\����&��;��r�dk^4H��H�J��)(�u��U��5�8W�,�OH��T��n�,0��Bj�)}$`��am@�5���!���ܽC��Q�͉���&�lY���N�ȶR7���1	`��\� �FW�(G(��V�-�D��U�Oeq�SV�`�k�sŗ����|G.�K��Ԑ�E͜�x�挡���r^�=�M/�D�V�k��>��;�����d�l�󩺥�V������ϫ�H]C`r����(KG �6�7L�m䓌Lx)����2��1Ŭۙ�ΐë��'~_���~�cb�'HO1��ڿ���bc$M�쮊�B�hKRz�W�Q>11j9�fz4�
:Gd5����PW%����nZӹ��+�{��N���H&�Y��-���o"�x�<�=�cYcd����(���'�-�����8�Lq�?�vb�3Ն25↖X&�(X�J���'f�ZA����+�W �S��4�F�|85�>n��4���1�~�� �
e��`����f �|*�B�Gr@o>b/o�k�*/J�}�[T��JPG.�JK�l��'���r�9��v\,��o3�GL��> g�=E���ni�%�M�"Խ�!�[����1�������ؤE��ɟ���@p�ࠣ�0EB~�{���]=ٓNy��;)^>2�5y����W&��������@	��d���N�1Q !._ckÈ��UZM��ט��[�d|�>����[�I:��Î�+�{��@pz)Ac���2�	��NKg����������>�Ww6�<����+=����� b����x�rh-����-��Ac).���S�O�5ޟ��7�_��t#f��~�G�C�L�I���1(.oh� ʤ(C�f��y�d�z����Q~v����$O�#,�B��@`V�\�k�f�9�����438ڑ{�8��g�R���.�0hSϜE��|��,�N���z�j�:�<Ӂv��h�˃�� ;��lc�łs��Y��\�q��K����r�4�c��P�