��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX����q:�}��>��\������FGm PQ�?���sU�9�W�iw_۷2��g���0f�8�5���?�8�.k ���L���<���Ƨ��bͽ�I e\���M��F�=G� �ut�����I�[�a���cO�$��XN���YǇ �5�g���r,��ne8����1�g������%�ygH2���s���ſ�'h����N7��%K��PK���2c�m'�/�s7�OK������ӻ��$޾�0YT��{O0���I(1��-��ԩ�(��|a��RG�#�Б��"%�AVN���L��n*�µ�\����xr0�*�����b.�]�|�G[�4A!�>@VI~�rӁ�;9@Cݒ��F�{*�ufV�H������z%��[$�!�1o�GcY�V��m3k2M��G8/ �-��G��ڃ+�pl���"Ԩ�Ml�1����*s��N�*H�oF��#s&T���9�EY���g�ï�)�f+8�M�.>�iԓ����Cӷ�Bዥ�z�dn���=���\���i� ����L�U�"
���4�*����!���E��|�	������_\Ǝ&Ȝh�XL'RِB&�-l1��o9�J�Mc�v�-������G���K��0�ߙ:ĵ�T�����X�*�Ev�[G�.�I�6���T/��u*��~Ma�kr�$wN X~LL���V�r�$>��r4�G��ǡ�hJ��)���Ixtz���M� �*8,1�M���A����g��s��1o��B��2�ȥ�����-Hۿ����%�/�{�UR׃�=/���!:R�A)5�Ӵ���J�s%˥-�{�ln@R��C�S̝	���X�� 3ݸR�)ls��{gL3T��D����l�X���r��[]���:rK𻽰�o�e�ΐ7���KIp��f^��fLsy���?kE�D�
�Az�\Q9k/kr����+�����L[�R�I880�e͏�'x8�]�B�����8����n+�ƀ��3pY�(\�I��`�詮�
	�k�" 5Jn�OX3���nk �'�ڎ�;���rNEp�B�����h�4H�˾�Ly(cxIp].1�������[�+��h�� �I~MҌ���'�QxE�=|��z�yor�,�(Nk+��r���\U�Hu�ZI�����*�|����j)k���n�Dھ�����Z����㑵��S(F�x�<N��T.Q�v��#�gUQ"�+<�=aXB��V29K��֋E�.�ƋHFVI�E&yPE�|�\��2v�_��s>"�BKi:��3�V���(ʨ��ɰp	�Ε�4jHA+��lP'~:�;�}ˁ��o���E������d�3�@F75SQn>1ߢ��i��&�ȼ�HS��*��I8�=N���u��K���Q�8K���'�[Fȧ�h�����?�Y�H�ʸF
9BN��owQ�/�.�+;��T����[>��ȫWx�'�
��S�%��a81_z�{gn��$�g���/���I]����XE{��H��9*���k̟�a����j\l"85sW5,Ʋ��q#J�WTȺ��ҳ_��wa��\�\E�d��ptB�MB��1���� �LyX��>���z��+�x�A��W/���ź]�P*���������s�Tq	с7+�m\zx~�Xw���p���fAS�Ƅ4�/o������)�^�ݳ�+hâ�/�x��b�9uClǘP1kf�8�sĻ=K5��wV��j��CB�Sg�:�`�&u��<a:��I���x��/�/W�·�%�&��Sd�n��@%>�Z{�'J�l��Cn\#��l�U�lﱁ�[�iLx|�C�t���ldy�U��TWE�-���]?2ߒ���)���H�o�[�d��D`�eͱ1#��MV�+u�5�ҒK�m­�y�f������d<�$�D�M�#L?y�h@��`�o��F��]�ʭ#6k���Q��I�N��0'\s��Z��8��*�s�w��|�=;� @�$(CS�C5����q�a�A.����	�3jJ�h���j��v�ai֗C{DjL���{�����9����&B������]���#.%��!�v/}~Qq��:O�g��([���0�[X�ZN�M�`'����OJ��JZ��@Zq7 ��i]J���Gp��7�P��J�ɗ]%�\k����4:<�eB�9l@�ݧ�V�W�ɯ}��N�X�|���Y��A�����2 �J�Gt�Mz���BFJ�
��&�J��?�q���э���W Իc�hQ�X�d(iZ�����Yy��&�?-�g��޳����XMpcX�%M�DkُJ1���wv�U��Pn�2��(��*��u&U�VYl��Q(�I6br$����y���γ����l&}:D����쭠 ��U�=���,��e�8%
����sZ�{#�J�|>2�QjO^�v����e��u��S�P����y����/���+A��Y�;�;`��f�p�Q逳hn�_�9���/��5��< ZF͸.�TY�f��baTu�fd��$3i�}�v�
�����U��UR�%F�$���/�����'y�&v����	;�z8�� v0%g�]@@�J:��B�� �up����J�_4�l	{c�nH�v��,;b���AI��U/��2F�^17]sԻ�C�#�m���>�a���K�z�.�҈$T��b�M�ņd>��D��`m�D��v���D���=�tr%�7��-����׮ݠew(������=� i�_ԉK�c�����^ Vo��%�<X_��g�m��+o�Xt�i�Bvq�-�&��C3τ���O�+�ko@�=(w��(�[��1�B��7}\�&	_-25�`,�>7�������7��*�w&��?p�^[��cӨ�Ŋ%����S�bn��?��n��v�jWl�3�{�e@(�h�e����{�<[���'
�qhD+zfu��enhw]�_~չUNR3~A&�6�r@w	K*Y#�^��b��v��
wC�
�jP>�m?���E��Aћ�!. dJ2}���n�Τ��T2RVDx/�_U]
4=��Q��"j��}�S*��xj
�t����I���w&��y�}m*r#���ᄝ�B�u^�%@����.6쳹n�2��BqAZ=�1��{���=HX)}�	�Lf$���g��]`�h��/ Ĕ�[����.��v���(~�K_�K DD]RDBj~/&$�=�A���e�;�G�BV����G���:��²aJ�,�n�yq�����
Drٵm���a�c���R� �BƑ1'UG�i���X�Hs��]�g/����l:�ђ|+�h	�Al���@T�M�o�������%N�`+s`SqTo�����.��z�\����Y�����Bؿjg�����p�F2�ǲ����:B��O�]S�k�� �h��5�r���|?�c�]1�����,0k$u<�N�6[צ��v�&o��͑4Y��`æ��dv�ӝ�Nf������?�I��ޏ����c/>3N*%��Wbb�K�w�ʿ��JN�D6x�={c��TwER	j{�]�J
!��{R�{5pC�vP2�Hi�|nG��o��2A�V�]7K�+pk�$u����f2��Z�
V<�����;: p�Ů)Ԅ�,@�y}�"�ӹTLz|T|��P]��[�:r-r��Zʡ�%�l"�|{1�<�����v�9w�JҠU.�B,�i���G;Ϲ�ȥ�fZ�j���3x��&�Vދ���%�,��k�%���.BH�e�l�]�uʧM����Z�<��/� �3�Xd��%�$��I�s}�aG�t��<��>�\�f���P�۩�z�|`�x߇�"��Vy��N�]/1W�rK�y`Y�0�)� qwА�����(�d�,���$k��n����!�^�&��RK�Q�
B���/r���2�y�8�*�,p��>I�,�W��Kt(9�DmpFw�4�0;k6�d��?��yztg�>�{����ګ�]�=���g�Yƾ����;�!U8�a`=�@���� �b��X3qt���Uj���[x	7I�(-=�����?`U��"^n�Me�i�\l�k!� ͼp.X��;"O�5��I���"��j��2����l'ja�?�f!f��FML��(�l��$PV��x�z�L���|�4A�s��������;��l��>�cP���	h��Rk�P��ؕ�X�33�|O�����J���Y��s�m ���/��^F$��?w���5�xS9�|aSy���75�r�%�U�S����/��i$)pW�������w�}��C�6��=ٷ�dk��7�7|S��D��^ɔ�6�}����<�<!5�څ�D�3��ջl�`�Cw�����2+���YQJj&���J��ygc?�����A��g>�e	e�b���!hz����Uvk�Q��
�9O��$��A��Y�2��N,ϵ���N!#p��D��Dzb���]>�X�z�P��2�Ζ�% �\9dsuŎI^�L�Cv@>C%����t� ��1�#�׾�ӎ���Iliatud*�Fⷠy����,
2��H�O�P�˖Ǖ\[V$~�DZ@����*������8QVG�����9���9M�ּW�@�@��jQ9M����5�>��z���ۺ @�a7�$XQ�ХG�̤<}�k��W\O#�<?x)�v��Ԭ�M+��q����]���U.���P�v�Y� �5~�)9�i|i�5ӣ�]5W�H����E�u���L���?���Z7������n���\��M�lGz�v/�2����	S���1�(e�\�L��h�t��hX�N�ۄ�GQg�Kى�Nfؘ���	"��8�Ro���o�-�}�������.@�O��[�N8�f�K �1�ܖO�lM@j�>�H�p���y�R�F���ͤ"��Jv�=S����ݢ�&N�>1ó���/2�9����JSr��F�I���*yD�M���P��%ju4�+@h__ߋ��j�S$,�w�ϊK���IU�X}�KB���?�J?�*[�t�@���/�w���Ӹ�^М�}s��2�j�����d7��&U��X����"B��K�$M.��_ �M7���$�$�E[�yJ�=|��b5�I}��s�2s������禧ӝ�@���J*�5�D�d<���0���t�2 Ͼ�@x�WZg/����k�<�����#�����@'ߜTI��׿���<H�D��0�&C��*G$Ԟ�����>�������0�G��L��֘��ؖ�?nDd��ˠ3���y7�'��2ꂞ s!� `2>�dL��h��U�#�{Γ�'߲�[Ha%��� ��@n������Y?ֶ)��C��F6J3q��.nx�y`�ϑ��U �2Q���0~J�[�lV���@.bT<���єx*�B��]�-c$$��&c�9D�<L�~��K�ˣPk�3B�k�ނG�rK#LH\��G4��q�YaX�4�j�0��V�$qy�(�7���m�ް9Z�Z��X, n��h�2��L������<1�I��\1���`#�i������s1���柽����E��� �P�����D �/���;1��ro�Lvt���(�ƨ��E#G
~$�op��v]���� �;�)M�V]v_�ҏ>>�T kNX����˅�2��T�X��������X���\��J^�D�H�6�☖��r���d"����@�zM��9	��o�Ir��e�66͘�oWW�f�~��v��5<��,܉����t�O�������M���f�/Q�
d N���E�����Db^[�I�!/Ho��� �W� pǬEХ7�y.;#P]���� n�7���97l��7?LO��-�w��h#��dF�R�iV�\ ��:_�[�I��ﴳ$7;�ZZ����� �j����a�` E���0���^�p����/�m��F��(0
)KC� �5'~k]ϵ�D=���ty�zF�qtQC�6[[��j�֕_�N������r��Ym���U7BU�T�IYB-�r����T�����Ԋ��!�2���έz���
e��M�l��7�Bf�!�:�D�ja&	O�0���@��ZAj~D�<~��~F5�g�����I��ʷ�a.�:�K�D�n= H�Zc6����b�i�!��N�E��e�Y<�3�LϰǷe��*��G���	��k��O�ce	G,B�+e�|.)A 9�P�ķ>�6��[^$�2�mp���"��\��eR������n���u�r��\��ߐ ]��X��GBu4�W�P���#����̘�ğ�������d�/N�t���G�����k�� ����7�c��B710�� ��8(�Ai���4���~���Ĉ
9��*	2��3/��k�~�t<�2L��Yt����r���]Da,����R}"}��ͱ֍4#��UaJvLw;:���Č뻟��e~�Ng�Y��2���}��"���^ui��B���H�ڈ�	5P ɗb�[0�e��yI��i8Z�b����P[?�&���S D�a�g��S������JRs�V��o�5�m� Ü�KmČ�b�{���ț`���wf�x�?��@��@�$l���!�m���}�����x=���q�3b��w��h+Y�XL R�X������iߊ�T�6�֋�Cz'46��9�E~�Yp���,b`W؏��,��U�ek��k{`�1?H��Q'a��7g���
J�>Wd�t�t�E������d+^�Io�	!-�4��WV�X$�w#��8��_)N�Dޡߌ@���CJ��i�K�������p��N�6:2��x:W�ժN<'�ƙ��${�+��)���K}d��;��al���V�`e]������^J�R9��1~��-<~�<�b��d�(���Z�&�FH&���d딸�tOF
���z��<�z��I�u{Ee�*�d�HA@Ϲ$Ԛį~b���� ���:!G�)V�z���b!|��^�K���l�<�&��-�C� >U4�
��0���#^�R�t3y�k ���T෵�4P����M.i�4�I�TX�3�=#�BJ�T�����s�豉��4�Z��	����ia?ߜ��m��;�(qv	Z2ujc�2&�=�j�X
=M}�*A�Y��Ti��ke�mqk�E�	 w��]N(&EM~�k��'ՎX=?���1������3���΁��~��l�/�QϘ˶� �M���{����uO�@Q#e��y���1���zE��{`z�9��^p��y'a�;8+@�K�;���@[Bxs5�*��P�Z3\|�m˾_�.��w���ꪮ�p�E-8/�cķ�ݜ˼��8�b_��V�"�[{��+�sh�L�!ZA��*861C�B碆� �3D�]��U-sCu�ܒ�xC�s4���"9��ow~��mCg���<x���C���A���̀�G���$���ԕi��ҹ��ڹ�B�@%����,�T�����u�R�B?@mÆ�7*�6 ��[I��O(YFywG�� ~"r,/�yV���E�գGQ��i�x�$r��O|���I?{��~69��;b�}��J���%��0������$���BX�>.B@���		i�	]��$́����"*##.��6)b��,ӕ���.q�u(���H��1�,����N��7�rg����j�<FF�������8}�6+9	��C��O_��ζ�'�}�{BHC�����P�8T@�8�e(1�A������l��7خ��]xߝc}R��=�k'���:�����Z�sG��/\��x��V�x�����_)ۀ��"���5�����HG�nS��uE��:��a���D��*�?f����,_��3����b���[�r��PV����P��5,�`,S�^��|��n� ����[/��ܧ�)D#+��~��n9猗6kt؉]�F��IL���eԘ��aA���ڡ���;NI�dr�~�'�~=0�F��DPZ��&	0�=x�}J,]�k�WX�ijMz�B���Ā}��-�$��w����W��lJ���Ɣ�㛒����M'�����V��Wݹ�Zs[	�Xzטǧ>�*uǀ䃕���Q����h��ظ:��Y�=ul��U�u{9�Y�ZH�d�9R����8Sw���;2>�d@ĐS������	�{{�Q+����a�mD�`��Đub���]���X��H��E���L��4t79,�kFnb� $b��LeW�ؚ��N�rw���D�Z U����`<�#K�oD�.k��+�>������!\����|&~ߪIVA߱e �۱�%��n�^#1������	"aސ��1XL4���𑑊�;��Ȕ�"��mRsC�-�X�z��_������:��*!6�yU�`hBV�_�|�!�֋�N��%��p~�9逹���T��R��?��2]����z��(0棈����FJ��b�-2��{q�g���҃J����(��� �A]d��í�Eϯ�R,p!y��Q�o��nDSQ5�3����S�캶w>�%Y��͜����O�ơm�_!�/��A�7�O�Q��PS:��ErM�!�:��:>�(��&���Wa���ֽ#�0�0���<�Z��""���z�x��i���#̺̼W��B���J5�n�Ͻ�S����2�H���}`,���:x,�B�(*!N���ԠB|V_&�T8�yR_ܭ���}$wY��á5��}]+�+�[SԙI��OyR֐Y��؋���ю�D窒���1-�v�嫢#��d�xU4�-����o�%~]��s�f�P��/��Jx�ܘ`��v	F�r&�C���(@���ҹ�7b����#K/��!�a��71�N�8�����s���S��p�s��aw�",��4;����1T��,\�Hc���P1G��>�Can��y�O}�Yч�`��*´�G����$��]0Fa�=�֭�K����J&��!Z�����@��q��ǡ:��
fU��Ú1h��ș��o�s� {�A����ͧ�K��Լ~"''�=-��f���[oF1�@u��#����y����)�#U���"�W(���S/�q�h�?n�?D��s��e�Q�OR����y���؊{l�-B�+7R)�����W	����t�#k��O��^�"Vc;l_]#��V�5��'���� jc��X���K���6������o�"�]ıK��EN�f�}=����;qPL�K7ǁ�7�[az�Ý*��r�����u�����^)�ٸ�3%����3�
q�n�0���{l_���ݭ�С$���Q5#i�H�\�G
p��n#g�-Y\�힏����2�g�՗�F7� �U��+pK+A����
�E��՛���Ը��y
v�Nh�=�bܡ�bݴ�m�o�Q��C�c��`bq�p������G�z�J8����-��	1�	�	m�k���MWA��׊�o��^ُ�|�$i��s~�j�k�ņDƯF��͜Q�7BqO���hl<�y�{?M([-��7���&��!'�\2�$<�F�'���n�P�g?L�vk�r>�Q�k���{aO��$P!�b(B�Q`�N�&�1�N�2�6�[?V%�{�eѺ��e
2i�S�%�*=�W���:O/�#��M��56A�R�b��DL��`mM̩�V����Vx�=1��>cT�O���2el��k-��c!�ӌ�X�sm��,��r٠3�_�I#qhR�;1y3���0g�SL�s���������|ۿ����&/�,N<�f܌X;⃉2�"���H�M���td�]����dW�oL��JP��{�M[��"�Yn��H!6+3�Ƭ�`�d���0׽���/�-�~���@�8@��o,��u�S��|��r���YBU������Ĥ�D�W�_�<�FS�7<mT��hb�ј�wyL9�����/(m�Š��3�M���rW%@��{��߆���hx�s���N�s�����;�`�:ӓ, /������'���)����*�� +���J�H#�V�J��*�&4��Tǃ&�7؇�������A|��p$Y�\,�3�d/�s���)�|.��ڪ^���8M�ύ8��rW�3�Q�|E݄o�#�Ym����`���h_�C��~Gkaf�O����_t�dz�n��6�����NXh�����6_y�9&_������5����r��a�@&��*J��kDaNK��"؟�t�w�� ]��۷YHYU�/u�ћ���ܒ�J���,F�hU9ޕ@^��!6"�vpz��vLf��."�����~��@�%�[@�Y6tZ�J�&&)��.X��C[Kb��~�:Z��9sOyGl�
,�)'z�~I������. Gm�Cm�ܛp���J�J�������c���Faִ��l��I��I���a@*�pD�����zM+���=����<��{���3w�~-�h<�����!P��~z�
9	��R���y�Q�+���P�k(r��X��}af<�z���Ris�ڈcJW,�����:@b�n�?��� ��ڻ᱀dܷ9)�Y�\:T�Md�����:l.3��(Ni���c���'�k�ߥ�q?����]8[28Ҋ�z �䙘�ʫ�YbZ��ѷG�����!�~R
!&�[=C��=��8Yf+k���.J�#.�b�z�sH�'H{q�V��@戣�U�Ū�ɧW�7i{�r^�׳8N2`�TB����)����\����֮']7m�ir��Å�U���`P�QJ�^y�)��7�H��Ipe���V�6��}$��}F+�iIn��O�OZ�dUI�Bk�I'�h����&�C��K�gX?|k�;s�,'żNMS�4CPh7ܭ�:�򢻥�xxlm�D�?�]��t���A+s	j���f*�Aq�1���'�U�Z�2�����S�M߀�X,4f�wpL�ͫ��p<�Lq����f~6�;�ս���N�V�'�1��JlS�(�,�#_eѯ�u��LΔ{� ղ�R��ԫ�L�V��׭����!}$el�h@�i�ݩ=�]1tB�X!l>�Ӕ�ވ��k�f�wp%e��G�b�Sti�w�C���^�� �:j.</���n�{��3=�s�f*�����:�=Y���d���I=�6~�D�����~�}[�w�@mP7lD�d�O��zg.�L���6��s�â�\���Lp�����+`aϛ��ܴ�Q�aC_W�#o�w�g���t��:�[�[�ѪP�/��U ��o����Z��[o���
L����<z�� &_z�l>w���Tߨ��F�3�s/EyeJ��Bƈ�*{�Q�O�(�gI6�ç��_����;=T��.��ۙѸ���nܒ��U�ƫ1z�8c�n����!���:��~a�嘑� ^�T\�]K���;O�U�4`o��δ�A��Oc���]������M[A��������k�d�*��3�[Ջ>DY�V�����ڷz��	�:��6��y�q`�_���+\
ӼPd�y�k��v�{���bZ�_�sR�pO�0l�����q-��ࡥ�>��7}7m�1��Td_��4%䅤��(�H�"y��n�j��2d{t��LCt���(��r� o�2ֱ��6Z���٣.0��ʨ�zڝ��m��jk⸈x%��?�)#g	��?S�y�>�{���������K������^����tfw��l�+)����#�=_�#�|�F4
7���X�O��8)f*oR� 0s����}�>*ꉡ�u��@����yOآN
	[�eJ��N��9j��d�"�I��6(�n����&���v$�8a��qX��~A(�O��wd�G�?�g���Rp��\��6��բx�����t�x'��**i�a+Ò�^���*g󩂾��o�f���$ʿ>b��E8���b*�"�]qV��A��jp�937�����Zr�c��2��o肎&�΋nMۮY����Y!���a~ۮ<1J?�����ۏ����
9�|�.��%��k�{
+�$�oEɔ!�z��_~�u��ih\�տ-�u��b�o���Q"�TT�w�w\����O�3��52OJ��:��e�����ml>=l�`B.>�$���� ݆���W����V��v��r<M�����bLf��EJϑ�� N˒��P�$�(,�64w�*�$M��5/�� ����K���a�{.��F ���Ik�vG���8]��ѶU.����7�I�$�p�ޢ���	����9�~�c�M���+a��cI�䕵Ǿ��i�"�[[�(]_���W��Wv�$�1���{D�{=���Qv�Y��/o`u��Y��ؗ��v�s"��Z�Y|2k��a$�:hh6}�g���8�ػl��^eQ�A!�eI(��?�)�EE3=2�w�aOvi�c_&o��r�V �N�5��uL�7�c=���Ts9�W减�:~M'�^[�c�����I���j��L=��� ���ے�A"}I�&�Y�x������e�+ʩɥ谣��w����������b��9Eu�V},Z��}��KN��z�.�\�8��J��p��-� �lJ×@����Z8f�5��u��F���T778j��@��m|��X�%]HI|�`.hu<v�V{8d�L����HRdyN��y�C$y�1�4��w�	(�"�5\���>���֋��u5�**�� W�����s����8��U��a��s��U��1N���@=����,�^Iwݳ����ǒ��蚦��f��4���W� �{&*`Ee�o��	�ޭ��M��;�4�ͥۅ�^H�i��̛w%�g� �DG|��Ҏ߲�|���+�F�;V��"N3�񑔷�n���!��� :�00>R��ޘ�֜ݟ}�`Gہ��W�k�>R�6Ȓaڽ0d��w�C;�F���v�#��Y༚�����>��`Ԣ2"i@{�թ�5?{��"���Q�]]g��.��ET����P�3����@HZ�ݓ��۽(��x��~�.���6P���5|x�.d��)"�;[]׍���[ ��z���p/m0�ˢS�BR��tw������y�[�3�� �m�i��϶"�Ç�$�Hd�_lZ������dT8x5m)H�@�2��"�x�g���R�����N��A7���#�	go�P���8b;��ͦV�Jd��(u��床�`�og��6*���U��J�!�Vf�^����3|�/$;�́I��Z��--*�zf���G��ߋ\�YK~�gG�P� �l�6�"�v�dOꊷ�>
g�r��y%�Z)f{ҭu�ޤ�[fw�~�'F���I*?�i�0�mn�h�}��A���U��+��S��̈�[�yf�>���],}*͝��-��J��2')�O|�<�as�
D��YP}�3[D@�ŖR8�gj����KD���?��D����H�����s�7	}+��@�^�I��#����� 8#!l���\P�#M��-���6��r"9Z��	�	��W��2�Ȧ���R�
G��}�=�_�#�&�A�@O~�`��ؽ�M�B|�f�a���h�13�ߚ��Ē�^��/�,UA5)��d�q�+�Y�H�` w��k�Oa�h�]*b�}�t��N�F����Bfm���"���7�B�����p U�0]�m���l굦0Q�'����E���d�Ѓ��O���W���_e���)6�f_��ڳr���A�vg�l�����)D߶�u��K�!3�r��jk���\��qmR��nUO }��,��-�饠#C0O��lh@ ���N��&.��U�qI�d�Hpu�D�V����P�N_��5�p͒7��>=����X �}���\}�(N���	/�z��!�~b �7낟f�<�Y+$�JI����1Qj���m��n�z%�����u|�v����W���MoC�2=;�&7��Z2�|4g8�զ����O��l�,�$hR����). ���5!��7��h;_������Q.�-��Y���j>�����
�ʴ�_+�WCrKP8��;�U:l1V��U��GH��s1���k�&y����=�$�bc�?�H:ګ'?;'�ٵf�<�/�%����t�$�W��g�a��&�XUT��18�v�c�%r��q�T��dA��R�y�	C����%.��ݯ�ʗC���L^�
�(b�^]�M@�{ĵ`�V?B7�2��{������1"+t���u�p�۩�8'��	tl�ɘy~�|P\�%L��L�	ed=��l���>.+m'{�����ڰ��r1w[Sƃ��:o,�^y��{�������A�+�ӱf^����*�#��p��F)l�xYas�9L�4'mm̶���ѧ[�4��̸sa�[�!Ԭ}dٷB�	J�ҜP����"ā�
�������>F:,1��{/Ni!l�H�>a����&�gc��u+��7�(1�o>_2ReP��X����s���h��pW�Ƞ�2�Hl)h�1��t�5|��?�V3 W���v�	�,�ZIV��.�`�Bv�����(��}0	�H��^]f����L������ǟ}���4��Ajw��%�J��1B	��֖�e8�O�79�5�i�H�U���`.(6�����O��F�%y�g0��vP���B_�e��z**��>�E��<�2G�M)��\0]�,oGH�j'N������Z#���΁�:�hX� �b���T%�NN��6��p�n8*)=]�aI��^%,�a'ؐc�>j�U���tǑ_��i��?=r�J����HY]B~-8�)���i�hH�p�ee���1���

V��|�hR�3���0sX�{�����,��I
�w�b����-/ɬ�D���%�]�O5��]_;�L�m�.����#������ԏ%?u��J�������j�GˈKݰENL����->X_;h�&B�Z��	�{MhSRֻ2��j�R�ͥq����9����49�����_�=��ޗ	��o�S���a�0��&=��ގ8�j��G�B��\k���,����΢�� ��J�y��Mkpj8q3�,�~��4��e�hhԒ��dm-\��4��vFS֑��H���$#��t��M`�.Y��q�i�h�u��T�Q6+�ZUs�D��4W�p=��/����2[�q���6�]� jo?a,;�N�.�o����Wf��s��a`<���N%Y��	�ik���z�����e��ؤ#e5E��O�����U`�����<2��努�-�k�3t�]q\Wp*\{9c`�S�cx[����^�	�]4��⁶?�`�Z��:��P���\��)�����꫇t8�j�ǿ=g�_�����$�qڗĥq���t�(�fs������i�R�Q��
�'�.����&<?�k`�x�ƢlVC6���zP&gix�<+�N����o[7�_���R��&$�AQzH��-xz���o���ZwI�e��2����ǉr�_�2s�G�Uʚ9�C>o�b���Ƅ��:���U�j ��*��Zn�Y
J�?`��O��8��m�:{@�Wݮo�8]v�%��je�����Y̐��f��2�3�<0�M���;����z�g}�ҳŹ�=�������f����#Z|��8�����w0����Q8�,˅m¤2���S;UT��(�6`�V
�a����_���>��v���|4F��p��f�����p�I2F�^��$�P�li'�Lj ��R��Q�ų���}<~�y�:���˟��m��t����>+����*�4zAɮzg���A;����8%\Iʻ֓+K�]�C%��}�a;��H~��"#�H��4���G�������{�6"�Dv���:2s�^�d<�"��h椲7�5��Y��)��E�KG�k�a�D^���J��!e�H��`K�s�ep�ZX��H��ς��ZR�A�x<�eȼ�U�-��Q�^��wj.l?��������>je�	^n�l@�7t��z�4<]��@Dz.S�?nA������˽��uCTad����2A��B{[.�Ð�*'�e�(D@c�\.������d�� �ɶ�Q��?�B�0�f�/95�žꚤ����;����;�z���2r|k�\ț�MQ��*�P�MM��W�c���S�K��6��ţ~9^�L��-Q�!Oh�Њ	�g��w6�q�K	��}�)&�P���)�f�������Sp�0�8�2+P�ɦ�o�Ql�&y8���8�/13ߋk���������:tcӷ[��2b�E�=�F��u$p?(�kk4��:�<;`�%&��BdoI��4�M31[� 2�׃c�%O�E�|��X=/��[�ܟ�j���7���fs-=ht��:�=V&G�������Z�c
�_H�Ǭ��YR�Μ��A�g͍"3���Ӟ�-zo�,�3�ؾ���Na�k�8X�&̯�v�{��He���U��߃�j��$��q`!�}���X՞U!2���tDVL���P#����y8Q�Ö'"}�b��D�y�r8��u��)�����qKI��G���}V�Ѯ�é�V� ͺ�+��(˩la�,x�Zg��~�����
�nι|$#w�q?ձa^c`�Gr[₿ˀ��1�ψ��M�9t̩���ġ5W�<�C��B�-�cD��4f�"|�x��JW{��$h���_�5�������Q��P#���6�L|m�L�k��E���+x���`!v��t�Jfc�4�繹U0P�/FY��Ȗ ��5�( ����1�a3�y�'�����;�"���'Ψ��
mF-��k��ŷ�c|���;��fT_;m�����	�P��F������Jt�p���R�w��ٚK�5��p�I�('��	��M���<Jw���@��s�gN=Ǯ��|y�}0Z����
�v�*Kv��?P�kA[Ϩ�Sk�-ЇڕR	�l��{A�26��J���~3��k>�k@7п_�z.*܆m7:|eԂ�=���Lɱ� $��.I��xxb~k,�zXX�[�.�S7�d��D�uaZO�܀#M;ƃQֿv1�,���Ȏ�m4�D~n�;�5�p@�'H�K��i����܊����fH#����w�Q���w�YL�[xWC�e���U��v֑]_UG��������6HF��E��2��ɰ;vYb��\�6�=޽��@��C�~n�+�i�a�]`���	TK���_��X+������^3�w�Յ������F��f�:­� F��X�\|I��5�K��sdƔ�QgÕͥ�׹YW=n3<�:AT�zU��S�Nۺr��=fn����i�M��K���B<������1��S�3��I��9]�\9�2RhȆ�s�p�9�`,k#:ԫ
S�����!�Pt�B�@�X���{���jD��.9۵�~g��4�\M8��\({��xI�8ڝ��@�)�ޞ8\2���u����l��%�~R"�}�D�"܍����h`�#�������.K�.|�a)%�i��)=��# &&��Wo`��@G9Zg�1 �9lt�XFg&78.�;�� 0�����U��{HMAZ����"r�k�9����ے�j�p���
lg_!���2�KP�C�={��H1��I�ksa���
�f��ν�*s�b��{\C�g�<�dų^2��Z�a,X8�.GCb�~;	�H�׾B#��#��V����/���1O��:A*\I�ܒ[Me��$�m/�2d�����`��e�܏l���	��i;��g���o�#���jf���]Q>u$G�?1�g3�H�)��0n�C�&�e��e2VM���H@��.���xG����v�������kG�)��)��3�P���V>�fE�����Ћ��d�$��<��q��^�]3n�zO���>�PK�h���5I���;�=U��dQ��%�Е?L�����6]��p��f�d�&sL����TP!. o��\�PKZ�����U�1N2����b��������{���Z��H�)�9�ҩ{���ڣm��*)�	��x��(��\r����~೗��$�0�=����t����vYȲ����8ʆ7ȣ��Zr��ab�#�
��q&�c6$3��TPc�{�(=(�VlP�n#ػ�9n!U`C�����5�8� E��Vu�