��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����F��':�ޜ�2̼ߵ2D�c�k	�?��lK���ګ�6�6K���}^��xF�u��hkp;���j�n���WVܫ� ����c������jɭ�L�5}��>��<L�=l{��	�Q�D�\V�d�s�囏���Qz��
2W6�ol��hX�| �/�������`����g%���9���/Y�ځD��uy��bPInb� �Zq����a��!���!����[3Z��{��0B�}���K9o�T�p��Zl�$r���^P�Uh���6��[�k(�3�~����NR)1���Nj*�:N>���y�5��-w��z��4�j�*HmĪ���/T��4��{.��*٘S"@'��A�4�Fa;hn��߸ň�Z�榧�m8d-�5ѻ�M�aSR4�����B�wOX*�2$��v'�T��V�C%�	���c�=��`a�0�f'�� �]�r�fb-]���Q���*y�i࿲l�=m�����R-�ĲXB���<0��\��KT��jEKL����D��4;�9
��}��n�L�2�C�o��B��LO CE�C}�gq�.��5�d�J�1��.���0�s�3<\���d%�/^� 2���o� ��M���������i��ﺶ�Fp����+�-0�q�0Yp�߀Fny����$1~>�)����m9^�sqѕ�ɽ��I�e\�g�I{����NoBS}�HX�e\��0]�X�yw$�~�<|m͐�����F��H�M|�_�!���/��*n�m��c�);��G9D?%(�4��e=�ޑX�Ra =��F�jA�S �Y����.fr$#��.�����C�d��Z'yV2��>��'u�Ρ)EM��"����bn3�B���{y�wZۄ�5���Q��{$�E�5�Ё6~���o�&�bY���|)˩}�YJ�6CX�����a*�w��#�`D9�R=���j�o\:���YB��1� Z�xČ��jMƕ��-;���*/%mL�Ե�9A6�¿E_Ub���)�H�}��M[��?�-�l:Z��%�t���&�o ͌��[�����b���G��6�:�7��k�%7�a��� m�t+c�Ԓ0������L���`O��8Կ�P]��- �~:,�A+F�ќE� =m)$�9"���n���!�0 4�	����Ǯ����3Tx��zG�Kv͑Eí�v14�%cI�¤�����D�ps��.}2�d"I�QoBHsj�z�5�*�tIV����ʁ�g�1�)"{���1�؅�ǭ؅�{�1�x��p��TM;�g�z�5{��زY�+�k�CA*�A��4��@��.�U��r�G����Ĕ�
�i�G����k#��JҤޗL����wH���yJ|�t�yџ���~�a��%���9Jė���Ekm���00<�ڦ��2�w{�k&n��P�}�MR�j5�tJ˄'	ʊEq��"AS���_f��u/��pg��ؓ�Δ�r[�"�a�.A	�Q�~���U��7<�+3�M2�
[��{-n��Pd���h�5�x�8 (W���b�U�61 ˁ���{!��|QRZ�9f-��[�����*@�J�*�/#�����>CA�w�%������W�ae��Hޡ����V���H�5F!�k3��?����)�a�`��ZP�������R��1�ހt�Cz���I�ܐ[;�0��0w�޲L�m}��b乎��+��[��J6��
�4�s=���-Z��S ��0��X�������uɃ��� �,�<��ȳ����ʤ�w1�����2R��&�щ��ĳL5��~�W�R[d�$�9���)�  ���e���\6�9� [�)��q%�"�6�lP�y�I�G�ZL/#�4���)�(/:u/��S!3������nȇc�T���ڐ��x՜��'zi�긔[��M�U�Y\x���F������>(���F��V4�[�Tpa���L�+]ڑ�hj6}V��{M�^��X��f�C���BW4���26�is�;�6�+Ht�Yc��_^-�O��@MS9��`U1�M�<���E�2	qv����U��<��
���${�� ˨���b��^r�pվE%�c�;�C��ƅ�O%JIw����.pr�p�I���"�򮄂��[�!�w(Q���ϣq��l:T=۵�е�P��7�1~7v��k�.�o�LmBɼ����A��&RrK��[�ɛ/�����zYŎ���T���.����h��t��ّXdYd�ݧ{3K�`G�.��f��`.�j������������O���>���E[\AE^D����j��U�ݝ���6�>��Y'`NO�Z�5e1�Z~�u�'Z�g|)��c������F�0T��C��Zp�$}޶�>�b=.fy�XE:�hD��.8,\`�B�%��5s\��_�:R�zy���Ԙ�I��`t!|f6̕6ǀ�Tӽެ=�6���RU�<���<�}���N���ES�a0+���`�δ�!�'����o�̷bW]�1��w��g:��gQ=<��/�&C�����A>��uJ]J�����$(��B�c6������v��4G+J��H�Ȯ�P�Ӆ���F�Gycy�&�J���^weZD!B�0��A� �t�=�:�Ǜ�?��#��'�jj�.�RS�j�ێ���Z��K"��x������\��(ҖZİ���o�	�GyC�z�&�%.^�$����8�v���"peW�P�9{:��S�q���ui�빘�9��u��@xl��>H�VYv���{[��$F�Z�����2��k��%ny�lm�ZT� ���]ay����B�)�����]BR��Y���s��jn�J�������#�m^��yM9�o�'�k�2Y[QL�rُI�浬��Jh��XwC�w-b��n�FZ ㏴ ���)Q�yC�+\���ķs�^�4��L�HE���Q^����m�̖+���;�y&�,�~M��e�q�,ʝ��J(J}\\��Cq�G��#-~k�[�;3o^�w�_@���H"xEk)SW�,���5Sīp/D�.c����f��\��=A�hڪ�
ĺ����9��Xz�9�5�{���V���g��x�\����{���r���M��0:VݪM4P�3��,�@u�bm�r�Ol�(4�L�`AK}o�з`�:xO+���g8���e��=Tl�6?(�=�sS�+p��(��'��h�a���䐽P� 2
�O+����<�@c�_�Q�=
%^
;���]6?��c�J_���ND�fr��9���۵�� �<�*���oYdLz�~,��ְ
b�+��d�]1lL}t4|ޞ�`?��w��7�u��w����L��ѓƵ1�x�����ߓF����-&�ֈ���g���q�]U'�SO��r5&�^�`���_����_؃�,�u�)�mO�3�b��8q��Bdf�*Q'޸�7��΂�vq�,���l��t���5K�,��L����È�����̩�S)��^��n ݹ(.�X�֒�|�1-:@��k���	�Da4��(�c�q�GZ_uS����	+�6�U�;����~A��3l�C��.�x�;lC��ARG�.<���($iˎ�'M�R�U�[�\��������8L��8wX1��}��\]��}��ԣDě�%�[�V����_�nԬ��!-n�O����𚙼�`���x���X*��<Lzˠal�z9�fU���;����b[G��YK�� hG��G�:*d�)ۊ�]S~P��eI��SNs���n���w5�}O�J���N*� 7�V��v4����d����'Fi���d��5�}�Ŕ�`��W_դZ�Ӽ����He���-�̙Ao�����B�;8*�\/�����u��*_D^���λ��sS��D7�Yo
w�R�ʬg>܃7g�S�ď��~�~U��R�ik�\��F	�[��VD�a�kP�ZE`o%���v�S�p�GG�_*�nʹ� ����Ζ���z��}"�����:7��$pۨM����}�sv�����#Z����[��wԈA%�"?
[Y�� XO�aK�j��S���Z��e�j��ӟ�l��+���&j^s�yE�9�E��w�O�]�MD�ն�`A��]������$��Mк��F���Q
��E��y�Ӑ��Hҋ�C��f9��_G���_�8ں���@��"tg<�J��r�c��-e�� �_��E}�u��u^��}4L_$˺��\-(*��@Se����I�vІ�H�6m�z8��
Mw��2+�*�@������Tj�����)�!ߚ:tL.��W��񻯈�%W�=�����F���v��MӺ�����ؙr��%��f������������p9^a�����W2,rf#��P���=�&$f)N�m�F�y�v�@i2v��n��.�����B��������v<��	Fx�J��B=�б�D��vs���'�n����i�
g�Dh�G{�]�x�Q���kS3�(�_G<��?h~)�/�F�r�m�E�P ��]��4��g�,ו���Щm(S�==�A+hC��Cgv�i�_[��U�G�Į��j������p��\���?q�>���t�����~}Ox�P����x~���G��.0�������g�H�)T�E@�\����~$bh���T�;���C��q��C���(I��q�ӷh�M�}�X-<�W�o�Q��J�ձ����Ww\�7O?��M�ۙn�U[C	P<r���7>�zG������^_��gU���'��c|X2'G�hܡ����;���iy'�.vÚ��l�T��S���.��]kP��Y����E���8G��=�cB��t�R1S�aO�WB1�a���W:+�/C"�ՠ��>��TB�y�FE��$�x�g<��n�'���mu0D#�%�h���I���O E�:������Ѷ��7`�KB���W(�wʏX�M�� �M�b1" ��������RPq ��_)������/y��Ȫ�PIM�گ��p>*c��L�l2Dr�m5%�zcC�TR/_�]��ݲ��m�"�9d�χ8;��S�+Æy�N�%�i����G@�5�/�D���絃�F04'ieq�l����'7�G�gi�J��MŹk([?a����_�&P����x�
�����!���T��S٠P�^������'*L�(�"�5|md�����'�����h�/��מ�'�`A�z�&[wi~�y��K�gwlE�s���[1f4�B�����//KD}�T�?�K�r����9W�ƕ�\�F�D4lw<��}���	y�r��?3�u�d)T�]tE��z�̺����s������\��?F���7���ڸ^�E�^Sq]�����Nǟ���TZ����^>�{����kg�����|���H�k�!29����)��e�}!+�%������ᢽJ�H_'���ݨڌ��\�_��خRb�&.4�'�kY*�+��'e��ۍ�#���2h�o�S��3����gA��&��(�;���oug�=���Ziy�`�,o�5�K�^���OŐ ׀�@.Z��6�)D�Qi�Yf�Cg�td���a��V�����zX���9p�B'�e�r(�M���(o޸J�!H�oxCw"���_�$]�I�O��C��$�D��#5�]O��A�p��zК�j�=ޖ����c�Nd���������(�nڼ<�t~)	�|O��[$��OT�M9����ڗC�cW��ە�ŇIJ�y�8D&Ia�O
/��,�N�H�b��V`���}�liE�1���)��������;f�HCy��Be��a�T�1�A:$W6���yɶ��ϊ�r�\��2s����M1���\��+6��'�;H���/�
+�$���o�8E��h!���/l��7��Z;��)����3��$з!�xa��w���!�|�t��&�óH௼���0&��$+�ۭ�Q{�X�~%,$�D����2��Z�m��ބ�e�.��D`Oz��AC�K�z'�G���X�U*E�$ߪ`�ry�.�z�7���иζ��`Q+���)-8�s��W݁�g੼z"/_��a���*�ۃeV��bI=_LV�8�G�t +�`?i��o�XwL@z�IfNp�Â��5���i�*k�a�nً̕�҅�-	�|�1е�JYou]/�C���`u8��8u����˅Q�h���d�� &�qN��c��Ɲ�A�D�@���);��&i����8.�*�y��Pv�ؘ�(�&k�G����|H�!&?5�!'~zxQg���B�\����3��(�E��A�Wŕ��Cw��K�c��\������>4�G�v��*�`��D��_BdP}y����H���*�0 �f���QN_�F%E$�C�vb�`bz����Jxs�+����� ��7�>�3P��}�)5�j�{2p��(C�W��D�-�.�w��B���C�D#���|�m��}��C}p��y�T����:���A�&�����}����zKȣ�v�ل�U+K�bԝ��Ϟ-��Zײ��ָl������f����|e�j9.K$��>��-\ݏΎ2;DE"� �z�rr�
�h��}�]������em��j=���"���Y�C���w�y�nA��eo�K�����;�|m��d9u�6sc�"$�[�M��d�x��ȲC��-G�����j����&>^�w6�d&���)�`}+�36����ւ�a�i���2{�q�>�9�ѧ�_�5��'�8�A$h���N��k�G��32=>su�R2����:�Z5��a�*�Ha�|�tYtX��@qNݲ�W��6��X��V�yF�#t`�&���+򪺎�b�[�Cq�M��\w(z��t�} G]��h���Io�i�R8�����р�����[{��ɝdq�l���Bs,��}a��u"` �;�G?�. �ҹ�"�-�="���ވrC�3.���?u#&2AP� \l��))�O=tS/�!�aƷ��0��7
����WK���1w�kS?��̞����&A�?���z8,�d�j48w�� d`�&O����Tp����$�z�����!3>��{k�u��]��kk�X�4���+�-�O@����E<G����y��ǯ��0��g�*Djv ����9�k�xsXԩA*>��P��?�?���+�hn�`3��?�r�s�W_�f�@$i��(vj�(ec$��,(�p qR�f�C�_�(8Nu݀P�d��a�hV&>�Ϭ�xV�A�	x���M��7�-Я�	f�����Jr��:�]A�p�ʡX��) �\�Cp���hŞ��b�U�8�.�Wl;H-�W���u.�kp��I��[7b�|(_az���y/Uz���u��ah�[�S�,]�Q�/��%އ������m_�}߲:��
|"�N�?�y������9X��Y`:��V��2>h��2��
,+�^t9R��Ŕ&=�cA�����^�\w���O���cy��9꣕#�O4?���`�;pwF�M�d�wC�1Ji���c��\��I���,l��Y�l��7�]2Q�)��<�	)�=�҉Cdm~!����]9!�9��#'p�A}�s����e�U���J��+LW�bEAk 4䔽�V�8ʡg�k&���T��/�����`�-nH$�^�|�)�`�(�M;]��Ft&Z:2=��k#�0%�;�\ݘ!���=�%[&�.�|�!��l.�?�"<���P�h������fG�$�/������s�o�E�	�[!���!p��}�����W\���g�uo8����1��&`[Ȱ��⥀_$�t�q�:�����o�7*���@�Y2>���	�M�X�Qk)2'�����F�W���Z��vBM��	�}��(�`#۾ӯ2a@6:��<wց�9M���N��A�kiFj�_Cf�P��\䇈�i��ڜ�!��Jn��N2�&gD���nR�9�sn޾��M?��Ǳ��{]�������n�ev����,U��g�v�f|#w��^�u�	VW�	L�nj�("3�$�)�`���91T�O�4P��F��>+Oy��V{[�����Ļ�<N��͛:�V:7N]Vh�e�[��)�b^(;~4Ѵ9~��r��3��8Ce�ҷ��#QH�X�:�AD�������TkGG�lu�"�l���4�]����PeS�P��#�~��؜	Io1+(aR���=�q�r���+���>��ݒ�r��ߥ��O
�U�V�X�r�N����F��Ǆ �Z�u�Ik'$nw;����Stc+m�<+��hy^�D���:H@KY�esc|��P���l0�=���\K��tbCQ�ɖ}��v� ���W;�N�/S2�^�#MY���汼,�
�Tɩ:W�r2:���_��c�kY�I����3�h�0�:y�L����2A��b��[��1�w�?�ś���*ˈ\8����3�*6$��ӱ�!�|�75�o�B1�L�ޜ|A�u�ON ��ݩ��> � ��uh?Ur�[�1Na�T��i��ȳ$�X�oV���q���~��8��i�_xM�M�\�������ɗ�U�A��Gv��`�=k��&ImJ����ֽ��K�fy0+\�]pE�|�E��)��7mN��s\@�Do�~��H>����i�B��Pb���=�B��:_����Ws!�#H
C2���+�w����ǒ��<	ɹco�|N�m[�����Ϳ撊9J25G�@I�{�Y5�6��R�M�7c��3�<�h� ,)ڪ�8u2��P[�;D��0��A���xI�pS2��#��%3<)�ڴ���oG<S�mN����H~1�`�-_�
h�8�ԋ`�<�;�h���tW�R�w?Zn�	p"e���:M�FcsL�@N��?A�V@R0z0}!&>���"�!`8�/����O�8����#���v�����bfӕ�ݤe�W(��B5�z�ױo�v��D�ti�n����I�*i��F���z֬��'����C���.�ɺa����g=��cSZ� ^�������r��/E-͹�;"�W�g�lX�޼��vꪇ�DG�`</B���e�jP��6�N�uB�nw��x�>,p*w��v�,��f����w!PvUt2dGy���,�9t&�g!cc�����!���YGF{Q�X�^���ߜ�s�3IG�28Z(uUג�9#Q�/l>�)pMH��s�{�����
��x�DkO����o����Fc���W����+�p��U���J��(�r���45D``�~���G]���J�:�L��KU�^����j�>T\��f�q�\��z���+�I�V��:_0#��Zn�2��#�'TC9��T�+�/i�`��X�a�X$3O�|;�r�"о��2�7�5�M�+i����j�u*	#8�|y��@���ŪLB��d-B�Y7&7����(�gw���_ų�^���m�B�sz[%ƭ�U���
*�e�V!��g���MK����N�l]�٭eCv�6|�:�;�1t�������F9ٝ<�Ϥ�X.��@Ax.l�X*z�];���'��1�#����*��["ȟvo�6[���aŮm](z�X&���>x��O����+���k�5�uV�	؟������J����?�Hr�3̗sL��:E�N�u�������I��|��G�)U���MyB� ���g���|lҹޏ�	��etu�#x8�·K�W~�ّ�]\�\2Yil�:�1�W1��������MGZ�VS0[�S��L�á�v��g�9xg%�ϳS2����ܣ�G�dM�v���y�^�n�$.�N�5�gv/�54Kǚ�6Sx�6�
�pd�J���Y���@�����1���F�e��:m��_��:�U���hH8��bD*|fb�θ��ؘ�"�b�Bk'���9����+3��.[_{�u9�B���Z$83i��� ����N���*2�O�9Nme�Ќ�Sz��_�6D?)RO-(�fՂڳ{���m�\x��d4�|�2<3ۆ|7�~%2���ձoe�Y���>F���xi{ǩĹd}�<刐b}y�lx_>a�`���ꬊ�|�"E�C�i��Ug�hW��.�Qo�%�+n'�e�s���7�4�hHi-]\�D�q�Z�Z+~�J'��쭜�F9){7&����!�t�Z�˰?Y�I����T9
J�D��
�?���'���D��#�4��P�LA8}4���'�5�aH�Hv�ܿ��tddR�N�	=u-d���S�5�˩��Gː)�7N����gD�+�S�_��IPht6��8EV�i)��%��&�h��16����k�u�i�w���Qx�����¤8ۣ�I��]��c-S�{��{�ř}���9��6ƶg�(v�뷦,�-�_M���+etiCfM}'�����dę62��[��0i�%�/g[¬K��FY�����i ę��{�`�V�a;͈�)1�K���#}�d5�8-E�[sp0f�� �*�y��tT=���B�H�����i�z�9F��b-��.�og��LOFζ��X3Ĕ!U��D�c�+#K�L��q�������V��/�|Ȓ�vĞ�xQ�����|dp��Y�9Rc���J�L�Eq��Qe)��}; �U��hL���H͏e䎾�������ulw�/i)��jL1���-�a��'V�k�}��:�(C˗����
.�%6���]D�Ѽ5��7�'v�n���|���( ?���IM%ޡZ��2�^�Z�%H%�D�m|eH1�K+��>����Qa��k"�Q�����[�o̼���?��V78p� ������|N+=�b�2��D�6����n�_9~��H�Hp8��������Q���X:���{cqPm���$�z�}�6�r�S8�R��?�578N�ЀNJ�a�pΏ�$5��̥�[����q�L���u����qz0;��c�p	�Q]�ƃS�NΑ��(j�]h��]��]�Z��'_�
Ⱦ��L��ғ�5W��.]>��ƀ���ɯ;��n�\���Ե�Gf� �˱1���42pst�޹�W-���!�0�Ph���&�
G�3Ua׍�}�u��+lt���?��t\�r��2d�ڻ+,)@�ߺr f-y���q9�	��B@��Y,�(ig��ܳI��a�Tp
��nŃ������I���������X���9�:o�;������j|v����ƾ�C��C��%0�|t���<�JK�R�=���C%2{�9� �f�\̦c���@�+d(x�3� �p�b�Q*����Ò �x=F�X�I�N&!J�1�/XK�M�7�i|���j��ϛ�WWI<��"[ڍ�+���GV��xR�C��C���,�[8��O�����EFrx\pL��d=)�i��%�R�G=�k)���R�;�S�ɉ6�Cb֣��c+���P�6J�h������t���ˈ�@a]��#q���^��zMĵ��쨢R-`NU�
6����APL�����@bO��>j��@Y��
�����B��y��ܧa����]���M�^u�!0^*��k��`�e��{)�b�����i5���D�
-a�]�>�8DUu�ذ��N9��Ouk8#�k��ԢlI�N�KxWefc��
�p����tCSz{#l~��E�ȥ�`���Z,3��H�{��86��v��1ҽ�"6��^�d��~���V���[[x ����>T���w��}��21z�:'���S�(|�2�� 2-]���7>=�ߺ���c��X�����{K�M��xҜv��$%k���2u��&u�ױg��޺�g��1*2��)��E��{�D6��!��ŋEN�̺
�D�CR:s��M�vh��p=:��W��c���%(�Ѵ�HE�3�p��]�����c[͟�8L�͵Qn1c�\w�:eh�%{fml�q��f`7�
n?D����k쁕�*�4�xO/Gc��l��E�\�ú���3B?P�?��/O׊zE�)v��t���W��~���3�W����Cۭ_�ŧ�aS4~S%�E��mԕ��V<��=�
T6�?�2%��Ü�B���}���{�.ː�@#�<p����g0h�Tmʍ�a�V�"䇷j�LoQ?�*$���?=�����Ø�<����0�0�H}�Ƴ� k���4A����X!�W��2N��_�µh�^"��d���C�;�Z�����c����y���n�^���S]������֗�d�n�*K����t��-{�/9Wo4a�_p��֙���jW��8�="gT:S������g=t��63|��J�&��&�3EV���!�2:9�|S��2iF��>\�%� ��R��'m;��R	S9���lM���ԧ����Nq+��-ݣw�P\彖��6�����c6I������S�Ju/�l���	�d�/�uJ�0��Aһ�]�?w��1e�^�"��p�ʚ[Xl��(��!�9ߛŒ�s�(d;'m�K�s*��;Z"]Hm��:�	�GPh\ľ��a�[�r9qG3����Gyr+�U+��&�����W���O��ǽ��l��6Z58��g'�U�Z�b�p���m]9=wW =��gk�H`��@i�9�9��M�ۀR��,7�/4��ɍ%SM�&�5���~ۄ$��Yg��2ׅE}�]��Q��W�<�U�'���/{*b6=lN�kjN��*L�`�y��8C�O�����_``����"�JH
��cp�x-����zp �b������:�px##��!�y�TQ�r�Af|�^�1���V����1�Ls G��Ս]����ֺ`��n�g��C��s�Y@+��h�Ǆ(��I�鵟��'K��~�4��Ov&�o� ��O�T�t��[�?t�[�?3�)�'���%,�u�`Kn_�D��d��K6����n��8�.%P��;Y������+Y�h�����κ�R�펿"�((�����V�-|�\?n3Ρç�d
ٳ����ı}����i%Z7ܔ��!�����~�Ri���i%�����4�B� �](��u\>*����%�&wl�G��P޷�D�|2}�W��IAGI����2 y%�}MW�������uK6Tb�n�����Ե��A�ʮ��:�'0���v���kU@�O��79��ߜb�6��濏7ʍg�R{d��j���A��1a=a)9���]��]�$�܌��M"`;/�gE���m�{��Z�J�Zp`���MeA~�m��[����+��SW�w�5���4d��`Ћ��� sF�kd��s{��<v�����ezi���#,�=��.���<�|�g7�����ٰ�tegM�;���g�}E�61�?&�I�殡g*���U�j�zbJ���;6ª�H�dm����ZƍA��q�c,.a�ME)~�6�� +���s�Mc�����|�C|��!%__���[)ʿ]�'r��������bhj;�[��W��2���D��Q��s�j�q�>�5v0OJ��x6�����K~��1�
�*�rMgR~�@Y���z��l���&��6�-��wN�������y���r�P;�ŌLECv+m��v��a��,DL�;A���^��z�t5bB
2�*r3҉$�a�*��Y�ꡉg���X�}~2�h�k��*���QFO�٥y���G�R�0	0�&U�qM�@ZP.M/4�O��O��v����RgR���y-�ߎ�sd~������ 2��VhO��i�w	a#��7j\�i�Ř}�4ǶmuOl*�<`���f��`6�S��'IL.�"�|�kcJx\Uĭ�w��A6*�}��%��oir.;J����N,C�$Ng:`8��>�g˺]����ܕRc�	�(l	�0������?��`���`�@y��a �T�� i *E��� �z��Nt����vG��@j=<MZ`[;��5Nq!��ٚ[�B�8il�i5U=b��-{�q!]��q"��b߶0|-'F,f-��6|��(֭n�g4	=��D�I�tL�̒��W�9.t:�o�?v����鴼i&�Y[�1�aBr����G�DȒ�
(g��$�P�d����f��W�t6E�n�U�����`��捍�\	�8�Xb&�V%ݔ�ڒ���%$~� [k���YTT��O;����H旋��s1^lG��gD��9��߲fm~�w\��ұ~���)X���	���@���^^��p)����rż#�<Cb0�ө�����l��&�Xz���ɒohx><�.���h"�C����u�D��Uy��jO�ȜO�n�2�c-5yc~����R����JA�>��٘���(��χC��������؛��/�h�x���M�q^9�]Δ�K�r�/�Հh�ُ�[s�������ۨ��>�pe��Ⱦ�Ǯ�c:#�ʵ)9�܋���3���q����n3�@�є������8��,��B��y�=w`ʶ}��pI܄,��L���@���[Ǵڇ4��:L�~_��o|�.t�֨�y7��v���}e᝱6U��7��N^���� �]{IA{�����,�n�� H��e��g/Ĕ�  ].�ʯ͝&?s�i����B9�������,J�v_������T���M��܄P�y� ՛ M{�%.˖=^�N̺XՍ���Th޵����o��>����;��{���U$3Xv�9����=]���ؠM���d���L�$lyZ�5 �r��[>�gOzU��Y� hi�SL�X���7��a��e_]��%+��K5�*�So�Xw}�a
�	{J�T���m�V�~J- +�5�O���:EҘ��Ł�y��_�D�_����Aў�P���H�p���v���B��O�fD3�8ɢznx����U�Rt��U`׈)_'R����Hj�[U4q�WȜc�v��:Q���K�Q��W,"���?��k�}������9��Rk��k�'Eq߷�}" �;9[����{���p�5� Z�p���݇?Zn@��=�.	<U�oOK�` )�QI���C[��7WS��2J������M���O���Ǔ(�t�e����v�����R?{���lՑ���焃t��h�/��P~�H��ъ�7�WB-�a�]��0K��`�%�͗׿�b$���{8����9E��ݠ{��ŋc|'��y-���2���q����T�(�>D�V}�_x�=�{�q��q8����!Z+�Ѕ�|ʒC^��R��<� V��Fc�6+�;z��I��\�D��z�9�\��X��t)Y(z�Y5�*�`��KuD�AL{7q�gsm�S\�G���:j��X�-p6������T�QQR�c ���7�Ђ�e�c�6FU�7������{�W������pD�$7����5�����&̏h���[�.�q�&��>��!��?�+�o��Ԥ�����&G��jωR��/`q�w"��[��To,�v��ad�)Կv�qŐL����z�$H�|��x^���c��K��� �T�E�W%c3�C�-�2��:}��#��9�^���s�H��1�8� \�!����=�F�`�z�b�W�� �^s8Q�^咙�a���N}�ـ� o�G�̺&�����N��8�.��z8�na�i<��A�֜����]�aH]�x#h��L}���s�L��Pnߜ\����n�S sp����!?��%Y&�ؚ��[�&������|t?�F.;�X�e��JX<��N�S�d-��^ ���W "�+�  U�����̆�4j��f�R��Cq���S��`(�]�iR�������Iz��*��?�9�89�D��q͡3�`7�:�I�;�$�24�@U� K�wbCH�P��?::f�5�?{s+eN���h��dwc��rm�ٳ�uDG�|��<�{�[5�@�F.�K5(������s)|W��s��^��b�挴�0�B�몭�_BKd
�k������NQ��o'-�.��Β�'=���k9\5GR�'�fƅg+�D��������@t,=�jb��'4�ɪ-�Y&�i{&�±,vbQڬ=u�e�tʲ��I�*�9nTW��O�Qڢ@L��U���P҂� R,8~b�/qʏ��E'��(��]F^VFd�YE�Yk�0{3�"� �@�a�&f,O��FrA���0?�(S}�|X�"��<+ф����A�tTGtU}i:�S�����)9�IԆ�`���B{8	��ko�/(9[���kS3ʌ;	�.4xN~�4��EHl�yA�p��iK�ኍ�'d�����ޮLj�-�G�Or��͗0@@�_ ����hK	\G5K.�@^.~j���m�J"̽��e�FK\�@��l��0�ַ���L���*�P�(�\ R����ʛZIE��rsت/Z�2o����ٹϜ�#�	�1EPs�Iq)����ɶ�Ч�y�I����١��B�QFԶ�����2�: �N�2�|��P�*�{�tۊ�B�����xw� Ɨ݅ƀJ�|!��%Tt�b�{I!�������,�i��P$�otmun���7SxD'@�dؘܲo\ǀ�'=�эF�}
����84�h��wqW:�c��Z ����.C����K��2F���h,-�b{ԉ`����V1�Iy0�\<�,8�*N4.z���NBd;�`E1�~��pи����6�c�ȶ�N��Y�[ߕQg�f[姐�p���4�_i9��}JAA�E�!?�#C8h�.���`�:�u�@1]�K2]�w��P}���6NjG/%>�S鍾<C�0��*Mnc�r��W��*<NƹW�lL�G_mh�x�y��s��1HK�"
�=h�h�S�� �/���r���:�.H��9�nqߔ��b�7t�U��r��[%��o�zs��݋H�7�-8�-�i�G7\������̈��e8 <{���dy-,�Y�J���c{���s<hM�T=�3
�E�б�.D7Esl�R���|�h�̴�<k<$��mh&ZKY\�$���TBⶭSx��|c�g�<5����?4Q�,����_��|#%��ъ�e2@Qb�6��}�=g��$�������oF}y��u��`Yۓ9�K`�>r�Z�� D{e-��ɾ-^�g�����<�x��`:�K�S<C�����U���K�w�|/-m2�3FL	��'0h�#T�ތ���=�!��2� �e��h���E���'���ec�pF&�����?8ؠT��xi�1�-L��:�%V�a!�zӻ���NL�Ys�W8%*&� ���Xm.�Tz�Y�Qg��,.��GA��ϻ@�'�t����I�4s�;]۹��F4���h".V��d��דJz�Ir͜Z\gV�)��$��Y���S� �%%ʽkp�����t�
EA	��q8w9�*]�e+g恚7V�r_�t�J``����VU�'犁 'nO��^{����<l�Eq$(n�x��F�ÛN5��zP�������1o�!�	�Qde&��E/t��'M|Fq����(�քK�%��Q�=�T�Jfj�K��� aC?�O:�]N���yGde^9�}�3�b�%j����IG5)h�6'�Gr=l��B��U�VF�cw���l�Mq"�ƾ7ea 
�6�b7+g"�"�u%�ԁ�U��`�����*hc�]�&@/���^����4h����4�Z�G�<����،<#�s�:$�� �LM�[֞���������~(�T�%>���iG^'LR��Ȳ�>���5MR�F��?X��rL8��$�HYaZN����~gcUv�B�JE^�K������nA��9�R;y^-Oj4�/1�92��g|�_ ��]����15�QN/E)�az�?�i�Tzn���.1�Y�|B�,��~)�fN�CߠM-��<� ��S�����^�h����}�Z�s=�\=�[oXz�G�z6�3[�P���g�zI����f{��=��q�&��<K���E�]�N�p�v�-*"�@/\�p�5���Q��O;q����V7�}[�2�����oA�.EcP���T�̥A�"�G�����-5	T_��@���
��C���Iom>8�?L�kzT��@gm���&Ep��b2��DK�{x/�V�1M�l�h^��QE �1-tN��9}gr�h�I�,����-<X�`\�� �Ё�1�ࣷ��P࿆�����/��2`�PӁT�fy��O�O��.�W�=�d�rH!�ҿ�"�񹌯��D��h�RG��MٷH�e���C�N�cu�j�����noXI�J\�3�w�
�*�u�T5됅�x��3���-7>�����e��jb��ӟCdxgR�,ݹi �?�%��k����DA�g�/',��_��C�\�V��8nq����D0�A�V\Ob������� q�0�R�Fat��˩�>��OCЏ4�F�X����|0A���k'�D]�}��N6c�ИiU�f��un�K��Vڐz������_Ҍ�L��K����>tl+�ƪ�)�rJ�)�2�4#u�m�F+֣�!g��7�F�>��̊�90�h1尿�b:�륧�Ģژc��I�ʮ<�">Ktљ[v�DGo��	�xQ��c���
�"!
��_j7Q��x�'/uz���~�ҸjlkV��k�kI�p��_��v���Y�`�j�Ur��j]�q9�M�Kw)�	л�n����ؔ2V(�=���R���V�t�\��t�[���ߜ��,¦���E�ۄ&h��h��翩?�v���J˕B6y�lZ��99�x$�e�n%�E�'b,�u��'��x�)��MLX�.99�۸��E�V �S>��Z+�o�Ȉ���C���-��$)��2k��6�S��9$I�{^����9�>e�_O��_�����G�]��`U�P�n�F/>�}Ї�԰�1pC�����VU�U+���yg�3m��3��Gu�[r�{Yn�f?�q�A�|AQ����{�3W���X E��Իdm��Y��Ĳ��������>Co�Cv����2�,Fr�̢kb��G
��<>��J*W\D~1!L���`a4�\��q�:1�6y���֦9<�@=H���B��d�5v}B,1�>��ƙ��[�4���}�w�&aT�c/KKW:�u'0$S����7��:��Ѷ%�gF��ONϢ/P��o�)�E0�vE�E	􉂛��s	�Ô{��4��<Bw7�-�f�"G�x,l�V|h]���>�gs('���	�J�e�_��`Т��m����]�Ű�������EЊ�Y����Ǹ�^�b��7�P}�'?�#��X�@��ad��N�n���%���48S��yt��۟x��0��E*B�(o��Y_R�ݒ�����R�:j��|7-qsr�����1U��K��$���g��`[w���s]��~��A�GK�|�F��=��D���2}�u
�	DRh`-��0��1�9�){���Y��ᅃ�y��w�Tu�Ĳ߰����]��[e���l0 C;�C?�)b�ʛ��I��g���d��,�H���D����"m��v��p�R,3�Q���t���3QE�uЖ� �%��2�Y3L>��S�x��>ݡ�A������N�"�䎔&���+��(r����Ĺ�3eJ���GDq�lqTO�,U�#�D�kR�l�(��Q��b慆�4I���E��TQˤ���!z�G���2��6���|��р��A#�3n6樹*�p0|D���#��ݢx�;�]$���s��S��^�ʘ�E��'��'�b"�(�
�mb6�i}ZQ�pH�'�s�'��0�d�e���X��G��Wn�7X8�7���sأgY���y(u���#�r�;�NУ�j_�R�!-ţ%M���֞�c�3jm��G��Jf�}����f3���k6�>��/p����膖I���s��W��Vp�E�%`�tzz�b)���n6�&����Q)j{`�ׯ�]ƹ9%�U�� E����=�j�K��-
�:�^�Б�":�A���T