��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�o��ȃ|s�Pq��T
��xG�{�a���<	
%�yyȈ%��!ݓ�������9�#$������a�p���8��dޅ�Ki"q�0�	|�t�6_���єR����d1�k2��k*0�8�fS�M�|=O�Ņ9k>��A9�.���2i��f5�;WcTƋ�oo�dbe�R��"�<��	{ڏ4�$З����X/�Ū���`�[�ѱVQ�,ʙy����)CřY��Cf
�6C�8s�ľ�.�E(]0�Yu���ѿXF.�5��6��a1��o��7�݊��9�Q��dx3��/+K�٨���k{`ڴ4@�+��]�d�4�G.5$�Di'�x>�[�L��/z6�cν�e����W��z��V�U5��x�ra?���Ŕh�IE��ϋ�)_T�n�J�����ގ�0U�h����>�eOERb0���?t$���tG�k[�v��1�p��NߥI�U騁ޠck[�����oq���ͺ0@�~���b`�LU�p�~A��׮� �{��+��8�����|� ?s�u�5��)�&.}�<΁ފ�����Q}����������G�<�e[Yfg��.w�V4nIYМv�Ƿ�Z7F�O�� $>���{��3HwXO�P��Ƞv�,x�k�0�|��P#��h��0�-��ET1k,�ŷ7V����E�u�ե<�5��CVͩi(ؤ�h`x��)�xFB��Sa��Mq��wg�rI��Zs�0���--�R��\��
'� #�O��4���tYFN�.̘L�����[����~�k<��Ƨ��y�<��D�#��E,U�y��m�֝�`
�3Nh���y�z��T�D��6���PO{�+�c�N����]�S�j=x�*��q�(�d��3�g*Be��D�d�l�Bs+�H���4=Q������`/ݯ�0�v�w� A��HD����0�]������.�dWnOL� +<2�P��Pu�O�(9���Z2@�Q�W7�;�1����S���_�r�7��YE`��k;̝+KQKSN-�n�kb�DO^�P�I�֐N"٣5_W�u��ȷ��	�ƌ����N9]E��>���e)ݫг7	0�j4~z�(��I	�o�I�A�|ҿ��!�i���ʑ%5����ݓ�g�=y�2�5
9�J�,���8��i���Uʨ�h�O�p'��ś~�$�@�=�q[�v����o�B�i��Q��G�Y��;m521 �樿m�(yr�לn�z���:L�f�<Ʌ�_��1���$\8�+a$�8D�L
���M�g�Fv벒�i���!cSr���w�0�9���>Q�UZ��	2�a�:-�1T"ŭ	*����-�/5�W��4!Ƚc�;��|3�e�����������@鉯�
2��y�`���;6��)n�l	|�%��'�ˬq��T�<�b����C��ÃcƩ(`�jv�]As�����囝9Q�E!*W��:�\SX��Vz���T��^�jl�s�>uၞp�3�oë���h�S�7����#�6��cR��'�e�������ۀTF3f�7���I�Ż�Ť��:T_����{�p#�ŷT�T��j]�N�]7�R%��x0Qh�G~G���ꈶA�~0�%�����X����T�/u�b�T��l�N��b_�����h�J�%���V�r�p�Yӽ�g���A���e(�	�ꩅ'Bs�o�����X7����_v�*�	��|�arHc}} Y&�P_�B|'u����͆�%���F�>\ɇ���$&�24Vi�ҙ��,�wV)��I���6Z!T��J�����%���>�,K��@!��a��:�;��ѧ]~/Ab�������ֵ�*����D�10j���;Ū	�}�s�Kf�G��7�Kj�_�Q��Y�z�.�L�Ǘ�>&i��:����R|�~{��JE=e�9�jPc��f�I�� ܌�����Q���L@�#�[�=����['�����L���%Iv~�JԚ��As/�:5p��0�{[�r�$���M7��xQ����/饱M��56�#�`F&���N�=��Z�@��]��#ȬO�w���S,���j#y�ukA��)nE�[�A�z5Y���5�a���%P���������wV��2z&�ňe�Ψנ<mi�R]Q����P����>	|1�>����Ϸ��y`S�/G�=�4$C�7V>��O��>��N���eT��$ ��y��2��I��@�+q6��/zZ���97�B��n����6�LQB��=K��+�z��Q��A?����/�.����b���l�)EqR�f�i��)䷫4+�P�A���N�*w�Nz�Vci0/|"c%g�(9� ������ ]Y����Ȑ��K~i`E�K�^a<
�C���[^�|9��	(����A�ޫ���Tز�cM?I��~�r7+�H���Q��rh*Җ�.R������U�9��Ꝕ�=Z߄�z������`+��\��$T��j����Sg�'�C��)y�͗s�E4%ג��j��oj�<p%"t�/��`F0i�+Ab�7��Ү���)xk6�� Y�5�&Z|,��F�И*Tс5	�a��=*NE���/><v`��8TQ��û��&tmd�P:V?64��F����Tf��8ѥ)���5r���g*w�Ԡ�g�a:��)���ܧ*�
��=?&g��c���=��}��q��V�����-�����4kl�Ɖ���x'������_�����z_D�D*Eo�J�*�*����GH� yn�av��MM\)����}t*�Z�Ӓ0N�-��ݱ*�5�͗��T���֍��m�Z(�Kg�nn~0_"�|I�,|4���U��f_ L�E
�?e�,A�q�l�%�71���eѼWޮ2wJ|�@]�K���w�IL6\�d�|���Ǵɸ�s�f�O�`������������=�f	��|	��B\WI*0jA7���4�'8fs>塴N_6����Q��]��3��Ԟ��ҢSo�88Tl}�Qd*!�
eM�1��=Ƈ��Q�Ů�X1Q#4^�M\^�/�R�	=ݒ�ͩ��x����b���c��{���@�;R�pGuw�j��v9a��`�o�3��rK���3�!e"/:��X��y�cӷ���{�0�[�l4�^���|Bq��c	�GL�L�S�gRk+�e���u4��ytwԾ���J����@��skAi�o��z�]�k�1Zp�p�T� ���98]���S�D�˹i��۱����Qu唝��t��6I�`��Oe��Bل����Q#�}C���4W�0cX��p�]l��]��d��a����\��7��C2*��3�1'j�v��š�a������������ϱ��o	��@��w����L�DF ?��g��}մ2�z}P& �c7����P}��	��6Am;�͇a\R9�dl��v%�n�\y-���c
Q��.Bt����9��x� �[\m�}�0�.M?�k	�|�>���㯂3g�$�B��ݯ�eㅢ����\������Eg����|��X3�[��P����7��)�4���������+�_�6��esb���>TزkF�t��Eē���^X����d!�!%fa�.ވ���Y�%mNx��S�3�B��ʍ=�^@��EPH��:��z�?�Ds�?T��Y�@�ȵ����k����z��G�Ǌ�w6:C��κ,�J\��Xq|0�!�4�f�*�Z����r�"��Pߒ��:�\�r�v�1V�1����S�"��~�Is��0��{=r��n	
�/����H5��z�Y��t#�������[1�a�d0H���_m����B�΢�O� R "H젃` ��P�+� z�B[����� ��j�2�v?<N��Bx�õR�r/���Y ��ha�,�4��ݭX�T�|���kZز�����ω2���GZT���v��5ү:���D��l)oh�u�DVw�
R�\�)@	&n�S��RI����HQT�h@�$zG����*�=s�������3�r�m!X��I�\�1�G�t]�KEt�i"Cdd�Z�}籠
:�Ej���m�i�ѭ����(c�:�2�vBɟ��i����6��,��b"�;�ڳG��Z<k��)�Z�5FEj8���i�Xl��x�4#tI�@�9�ѐLw�fQ�������/��}?f����_
�����Ix��|��6/���0��02��������������:ku��I[��'�j�w� c#��O�cb�7*0r�4�_-o�8 ���?/�����2���Fp<�]�����l>�J�g�eĞO	|p�����e�<��Z@Î�X�Y;���F�\fxy5��⫝̸f��'��62�W�ފͲ����԰�6؊n(݁�v�3e^���]�4�ٗDj��0Y"��T+�8��I���`��}���	z$��D�5�BxQ�0/D�.��Rd��C��;2U'>e�/H�z�.��OA�[%�ͧf�43B��ޘN������l�\.�<�'����]K
p{	���."X:U�=�Z�Gm�M�φ���ع\��>�3��]�T�JԊ~�Qy�h|��9	)����0Qml����=ϧ$gcZy�tR3j��s3��W8/4�;!����jc���*nA����]�A��-ikb������2F�Ӿs�3�