��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��x���y���F4˰xQx�O�u�x��rQ���%�5��,�!�*���Ə֜#��<@�'��/�=�Q��Z)����y�MG��/��V=w�2ۈ���]��ٱ���$�5��E䰤��f��/�-E���D�;�����:1�t��L(�;4�Lp�X}@���8N��*���rZ�g&��r�9�Iװ�:���1�������nn��#��;4�79z����o���g<2������Z�+=�f�p;n��:p���æe�M��H���]�/*w��3���BoA�[����s�f�hP���
��;-&:�e0�!�<�6���� �g �x��l��u�0��3���$�-�a�P�ֹ<)t���S[���J�._���9{�������I�W���=Ơ=��.\�e���ړ�(����U��6F~�U�� �\Bud}���m������%��5o��U��U�y��_���H
��Adq)�V]�i����/,�����u|7��ŧ\�l�)���M��J�5��a�<SYr����>)�{kD���ы��ﵬ	=l&j������X?��ln��]vGA e��|9|�V*�?I�{1�,v'�v�+�Z�7�{�]����Kb�cp0�2N�7����[@a1+Sbo��:-�d�4ϪFk\=狅�5���9�u�`,J}�O��<��
U��!�a��C�m��y2JKu�P��D�5�x|uF�vcB}'/(y�v�j?��8�O#e�����գ��<�`�>��nr-���)�>�k�GmY�+fD�*�3�3x
�biV�#��"�����6Ͷ��UvwMR�5��Aܔ����.��
�I�V��W�z�k�K�m����N�u�W콳{Eϡf΋5lf�a���W9��!����LO�������e������3Z�M��%���)�=�(Ńv�q4�׿�!�h+k[���-!�-�c�;�}�8�2��m/M^%�h��JX���+T�w��l�;d��{��3;�B;D$��I����F"z�b�(C��0+�#���	l�fc�Q�zZt �k@p������7��oy)M��x�W�'#l��.x�"�C_9|mve�-�I>(a�)��S�`�1K�eN*nJ'�N��Y��&��#Ϙ�Kuf2��-zII��!�(���|x:�[�����Q��Ʊѯ�E������w2Try��y̾��8�����wi��z<��B.7ﳚ����&^���N�]hy��MM6B�D@%�`|g�3P;}�k>��7���v�vkrO����W�=����'S�Ӳ-���ݢ)���眜�6� ��}��͆s<	��Z�m��讆��U�	�6,�+E�;J5�"l��E���O>��4��'���ϔ��q�L\녬;o":�c�"���S�Ik��ZL�b�ї�����ǲ�"���˛H�u��C�	����<������"�)��d�h�.(՛ɔ����&P��i��q�۽f���T&G���[Cn1�Jڍ���n�ao$�)Ż�F��[���i�1/~���1�>i%f3����|�܂�R�`!�� ~I�`��ʨ�o�"�jK.�A�%h5���é���-�Ua��@ 2���tl��I�!�YJ3���L�K
��Euq�����%�f��$l�Aڣ�6/X�{�i�����i:��6�K/�n3�RFx�"��5�ю妋]=����>�2�bB ��%[�ȩĨ)�-%�b��z�Sr�ߤ-�둮�U[ٕT�0k7aI���0��#!`\���O�=��Jh�V�z��j M������� �����O�,�X��OAn����V�4�L���M��p���#"�tc�&�Ȉ�hh�*�����eW&���<v.�ZL�d�:�w�������
c�?