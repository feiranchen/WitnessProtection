��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f���*�x����W���jY2��'k�c���x?�i����$QbT"`�Ȋo(��2�a�s�q��S[Y~ ��O8�0Z1(�K�U4x���H����S���?�<Nm�s��S��w]�ޢ�L/D{"vf��rq�>Y0s��u��Z�l~D��oJ��o�;wZ i��I�ڐ�Q]��=��!��5��ng �E���>GCqܾ�֞�L�I�j,�:�ǌ�=_�7j�W�s�tϼ}�d*��m�����AJ=98��%"���_H����߀{��躴@�j�\��o��Ы���[�W�R�L�yDh~�?�+�P DA�b�ԓ���d����Bd�t]�E������&�J��.�E9���[a20+�f �L�����z�� ˣRBJg�`�i����8���ܱ`�H�z�����0+lk�Emp��9�ʝ��V�g�ߚ�6Г�x��%�����K5q��dU���w���&�J.dcX���ĵhS9�T�e��[�#�U�=HCw��4�1�,[���˨�x����Tʣ�v=TU+cO	{������`��DSവ�z�5���<�4���o�q���Π�+9�~�,}���ޒkA�lǷ�O4ՠq7+7�?n�cD������t����X��_9&��PQ3�E�M�H��+
��G\%s���Gh܀$�x� ��7��ueh��'���u���3���=��..�ͅ��8w�-YGr.�[�MZ�J��Xqi��f�_�j�юW��mGX�����d���	]���P6!���F��˩,gh�AY��~X����y��O�����yO}��{���~��
Z�`�ŀ� ��i��K��K��Y�$_�<3�p�O���Ju��|c�lu<F�'�^�Sw&�y»�=�I�FS�,��jP�a\>���S����_*Gә�����~w��ǥ��� g�O��Ȗ���B~:����cT]8PRYE'��Q~���1�(k�( }�+)!B<37!�kQ��w"s2��������k���� �g��Mt�s������lq5����z"�x���F=7B��HεS������{;$/r
�̈�b��$k-�ۛ)��CdH�g�C��&𣁼hF�_-`��rIG{/�=*m7da�I�j��LJѫ�Ua�v����Z�ۉ4�r�f;���-�e �q.s��)X
�r�"�����WQj�K�eK���=E�DH/�7C͑w�7{�=$��P�퉋��7�L����E��kv9�C�?��ŗ�R��j���Oa4��rz����	[�-m�	{�4���S����$@�<zO!>�]�����hQ����[�q������#hW��0|�$� �X��� ��՟�~��(䳊Iv���++����ʆ�b������f��]���l;~�"\���&����Jg������ة�m]=|��F`C@�&���@��g��L���b��9�78��Ͽl`�'݈,�L0U!V�B�3i�ەa�h�Ln�4�8�?�ۂL�JSA��rd���/p�1�lM_�-c���`�� >v��8�l�EQ�r�i����v��E.8�#��L:��X�����M[D��L։]T��'�&�1�Ǌ8p�'ܨ�E�보����w����hi�2�|���>�^��[���:'�g��bv�b���o#�j�nd"!�8�����Z\��L{@x7s�~�v|+���̎���m�6Q����3عûT{������a!�˚�k�-دD��42��/�R?��4o�����F��N�f;U��*.$�����9��cNBǡs,���HW�����W���g��W�[/|��J����V�\�S��/��tp�{o��ƈ�A��H���IX�Hgv�}�yi�Sh~����������k�8��t:_�?����k�G�Z�LE3�$�����<v�a�w��}*g	���r"�N�%�wւ�@���0R`.]�"�=5���u]W����]e���P�G�g�g�A7=��d��n�Q݌�h`��-K�|����R|s�y��*�W�lbBg���F�n � ��SF��]�� �f��G2IMs1f86�[K?�p�eh��1�d-v��Lh�ߵJP�G���Xx�RQ��]��ݔm#�,%nk������v�Q��P�� ��B��r�r�����VFhk{�ȣc���A�NL�����(���r�! i^��K��4 ����}����dDV_��n���nj��B�v9��)�m�n7d#��S�I}���wԖ 2>S����=9���?;���ǹ�J^�{�w4g���c���+����j��IٽG����7�J�� >B��8����V��` t�T���g���V;��k)b������4V����6_oǼl���-1	�b������}���K5G;
����Za���
*vȼ���-�h����<�2��N�W�^����!7� nH9��nFg�pmCG�D�J���H�1y0�»���n��]t��kP�4��j|o�0�}��^5z��v����Q!����B8ja�����%ֈ䉻���:�]+Z�c�SV�~���_m�R[��tZj$�lG�ķho�y&e�UW�sV�z�w���o$jJK��G�lh��
C�9�1L��	��P�4��bxn��
l(��jk��|C�U��ڡ���&����໷=����{g�I�ПO(�=>�����H�.͝���E����+!�B����7D���YQZ�&�7�J���,R��@+��j�J4 8,>!���w��F���kq5\	��R�;Q�+��T��T[JB'��K��jB!�y=�A�D��뚊-+��)�/v�	\
S�i��V��I��/cȌ�ܼ*>I���i�������z�P�НW���y~H�"DLTM�����GU��&�Ι:��R,v��H2'���j'�ј��4����!jZ�#J:t�öF�gCȊ����������9�w��=��xj�����\�5X��U�<��T�kj���\�m���#N�޺���Q"���%���)���Mx �.�K<Y���M�[���c�^�]ۚ3qky���;��v���C	YθQ�YM�b;|�{}3��
�ѧ�̕G�P/�{_J���fZ�K�޳6|R�T�&b����HLH֝ĸ��A>��t�!j+gypI�*��O���!�ܞ��H�\�ɲALc~V�}�NI�-�jZ�B����$��:%�kV�'�p���s;�^�Z{×�"P��5Wt;T��П��}
���c%��s�ӕ�-f�3�W\�p���:nt��3S*��n��6N�����A=�[DnN8���
���t�jf�-����
Ʋi�������d�*�b��~L,���1�){{s���Y^Y��m����
0h]ڧ�d֥1S3U�_bt?�|��,�� �^��1#%�?tYňP�h��qg=Bn��z�QL[�m���K���c�n�e����9!D���
w�p8l�)-"�J������
� ��kq���g&	5�w�@Qeս����ٯ;c�K��,$�Z]ߣ�w,��{���:�$�%��g��߾�%."cA�1��|�3$znׁ/v�B�����/�WB�F��*���E_^t�~�6N�{*���aΗ6�5�G͋�\��"h��H5yb�u�>��{HC43�'vɼ����9�n�/���Ϡ�!�Wq��X6�Ռ�RTHd�,	�ոq�k�W�Z����J__@��bo��u�@AP{������{�����5�KLc��Bv�u�Ee�&.|�8�j�Z-�W��Y�5�J��ea�X7QF��j63�*B+pMO��y��޼���Z~�സI��b j���(��dpa&���k��z=Z����Yߓ��53ɬ��y�]�%_���RY�:�����)ۉ�U\x=�u�(`#�$�k{<�*�N��t?g���;Ϙ1��{���)?���e�s�p����n��E�CS]�+g����������2|���Kl"�+m�����+�j��Ew:£W8S���;2Q� ��<8-�S� ��%PI9��9*�X�f��#Mh8FI�	/��w�@T�Ž��	�� ��BOڶT�.����tB�d�2�`�BtF���ܽ�qZsL���#ӵ�Е@b�BUyh"8u9��Ke% ���I�c�*	b���m��$'�^qf�;�{��UG�3鑄| F�>��\˕��F�L^�se	C�_�� ��S�]6<�4��ykJ���5�0$�.+��2I��5����m���=��˝��`b��,�TVU�Z*e%�*��<�޷�7$A~�!�r�9���w	�hYcN�.��H=�F����b�>��w�7�5;Ϥ;ԡ�AB�����Q�%�E��n����k���&�Vt�*�eo���V!�dx<[��N��٠���p��[R�A��!W�(�����}c�����c5 �!*�Qj��F8�	��鮋������8+B ��,�$�Y�h��l%�/Ҙ�M����� v"���K}����o{Tud�7�PԳ��Ķ�q(��Oϼ����9Ks� �|lv��OS����<8<N��f𖏸���(|(kf��|���d��T��ۈ]��A�q�����s�{�Rl�#Xn�f�'vNuuv��O�-y�U���{yT>�/�gK@��97��{']��¸�rY��5�nu��p� W�?d�vۢ��5�\<� �1�.6��-���I�=���:E��o�M��²�E��� ��z���"��as0�YĞ:��#%^�Q�b�w)
q�r�i����9!���?l��hzmUf��D�mMLMF%�-�0^��N2��oq(Ep�1�k���k��6̷_�� :���(r�Y}�sW�޸����(��-btN>H���A�ڠ|�.܉��MYL<�J�A-oz	�\���H����w�29�h�t;�)'����$j���X�b!���sh���ϣ���������JެZ�~����p��O�w�����l�J����R|+���I0q�Jr��֠u6��o�+4}]�*BQwJ����	!�a�|DTp!��7i�|���^,��x:����W�$p-�X���\9�+�N'����w�����q.��HTA�g�J��� :Oe]�g^�ɓ�x��5��#��W�p=0`�yk��i��`,�.�\�y�-��߱����ݮ+�%�ƋI~m'aS�:��gּ�K{>Z�e�z��i�}咜k�ax�1#�C����I�N��ͧ�mPG�G�4m���r|\���IB�^M�i�2b� gO�bׁlv-x�;�J��,��fQt���:y�흺O�lM�㏧�c�.�F�+'՜��M����y���gмw�~����!��	�\�m43d1|E߯�+%n�	���R���L����fÄ'��t�!rm%}��0��1Y�s(H����#uްQʍ��$���<)�}����gJ�)�a$@�}Mڑ:�����G�n�����U¥V�`� ��w@���$<C���M�f�r�vM���0:�����J�� �����g����/[�o!�ҕ�?�N�r��&4����_7c�Z
��@��cT<@/�!-�1٧[������*�?P}�%�!X���o'��g�՜r�{ş���<��z�5��WuEvl]2�Ѩ�`u�3���#F�]�y"�[�o`h=�Ԏ�M�%�Z%��a#��7�n�d����a;M��PT/�N��5����'(�a�S` +/ů�8�6O������%斪|3B]5j�q����Y6&Ċ����
r��
�ˢ��.<� �Y��t O��D>�WN�����~��NYp@�zԿCֈ�Ϩ�G&�tŨ4|�wm��q&�7�d�.�&�Y�ym�n�zA�?V�9��"���&bBw.��`8�7k��~�jʢ��n[��:]@��U�3ft^v�ks)���F}pt؇�V�8V�1�(S����|��a
nC�0� ���}BU�iݵ�=o<�b�ʽv�V*� ~����:��H���D������aSĢ{G��)�*͏=5^�f���q�yM[��b��t�0��{l5�����B�^����Uȩ�N6����[7� ]8,�������!Y���mx�[���/+t��9#Z_3`"��$l��#\�"���`oi�d.�W��Jq���'Z�������|�l�+�P?�4ǽ�;�L�O�h��:5,���ט(�b^��P���p�^}L�	����'�0I�x��n|,�����tX�һX1�͓�k��ܞ�t,�9�N6���:��Q���/`Dwjgī���7)0�[D��O�_I{�AexQ6w�F�q�����TMh��H���7�at3\HV��yy�CM��X�}���ZDw�8Nk���1X'�Yz,@��ae��[̐����jX(SU�s%S�8t�o.Ly}��u
hs]>��$}y������R˒&W�A{��leO��w�[��<B���b�����|ҔH���Y�l�O�9�q��?�Հ�up��O=���?|���JU��ft�;F�E@K��槫<W�K�Vk�/w�V�ڝϚ�xM�H40�g�00������0$�<�U"�Jp@`���vIx �ҷ��:��$�kW��鐂�P�-�|:�@�nD/�AGܦ�}B�����J����uR
�1F�2���틻�)�l��z)���D��+c��~&g�{�(!�Ro"��-�t�Ӱ�MP8n���`Rԗ�'-���LO�恝&�����h�+��sQ�8�Xep�(��C���L�.�Ғ������a�G��'o�R��lO�J��-v ���N�٬9vg��W�?�nE�E�����5wkH,�T/�$z|�`n�b.��������T���zS|V}l�u_G�4:w�r����Q�����hn��7v��U�D>5�����q���e	 qv�W�Zg��L~�:��)T��X���ؤ�tAJ�Ξ�a)�p[��(��Zq��J���40���Ԑ�u�
��4�;l�����R�`����)���Ed��b`(���=�A�*�,_~�"sí+Um�����vL�%<��h1;�4&��eXv���~v���WWh<�J�|v0�����H٬��\5�#T�ū*zU?����]�Җi6��`S[�h>"�?p7./��%~1����n$z&���'*��l�A�eČ�:#����VV�Di]��k˸\Z������[@�e�J[gB��r��	�H�]G��q���w�9��9�P6�\��~o]�jd����o�7�C
��0X�@i����BGڄ5`A(5k��/��E�a��ϤjtO<^��i�(�Y_����_
�*��;:wk�Q�uBڧv}Uf���C弯����J��e�ډ����{�b��;��P�y^��oI�O���"������N���ʣc6n��_k�2�Dc���B���+�auQ������u�$,o�석\��,�n�5֭M�Z��fm��?���!e��9���#{��+�ok���^�b��J����cZb5,���M�դ2;�آ��붯=�W(��V1�Ec��[�$C*:���I�1�:I![����mh�ϫ�O�e�Z�.�}q1c�:e���ǣɎ������H��~���uO�»Jh��� C��Qf�֕�[�?����@�X��M�J|M�}��u��Go-�I���.y�lFW|n%�1�$n�&2�dj�V7� �����?B^I��DZJ��X4�x$���ULB��m�:�j/<��/l��������_�h�G��kʥ����",�wS�}:=%���3l@�t׬	���H�
 ���,A�h�
U�R%��Gm�\��ѳ��4'�q���G<,Y�pQ��ߢ
^2q�@�zG�?v`�M���V��7'����!�E	��o�.��[��ir�
�Gr�!#˥l�W��Q�le�� �U�ݷA��
����	�U��5��3Ֆ<-{:
�7%�W�U{V�o���샋G�BS[��]���:A+yU���4�����zQb`Ĥu<���oƘkݫh�]�6�M|7 �1!��ǰ0���Dx:YO{g&6='������lk���4��?�n�}&�i����8�*�}��u�	���w+<;��u���ҶF�μc�+���/��msk ����e��
9�)O�����!�0��Lznh6�XB숞��!L�B�>�L!����P���������Q�w9�Z���������Q�e�;m �O��� nD t��Zq������g�����M����\Y�u��U�4��m���`'7�$�~{Y��/F*���Ka�*J!�v@*�����5ۋ�I4�w�D����Ÿ�%B�/x�=+��kAا�Ӥ!c]uJY�YzE_��i!/f%"VN(C�˃Pb�0��=|�{�r�j��A��^"�g?�r�+1m�O���&&�rZ� .�\���2�o��Oc*�Q���n��\�!��B���z���
����@�5Rꚷ0s.��[�%>��<�O[-��t?���wej?�����]o�"�ןv�҅=�_��9���������LY��<'=B������+ILX� �4�y��A� fqSD���,��q9��M�l��`��	a2�����M�dN�r�8�a|]�䔆�\�{����X����I2c��`�y�% X;}os�_����-[�������6Zx���{�|l�d@�G,�BF��	����m����i�؄6�����]k���kTX��H�{ C(R�aȁ�BW�I�w��_U�)�d�{�W�|P|�ȷKU��m]hr���69s��	~z=�D��>4_���&��+W4���9�^�J,�/"'����q�ܹw�p�$�/<"g!Q*���RTݦ�P��)�Y�}�3U��f�`cs�Y���r��+0-�����,�j��R�Yˋ� p���a���n�mҭC ��OE/'��]��
�U�����j�N�q��L9?v|-	+pf㡉ԛmyX��AI��)��#�t�(b�Tw�S�;?ڲ̲)1M��~"�Lq�%�Z_����e6�*�X��5�`�'�<��OnL����L��@R%���� �*h=�%`X�rij���gf�N}�K?��W{�"�{߲�w��sf�9�u@P���cԾ<抶�
'� �� �{��W(m0J9D�ƍS(��h��9b�=�.��Ҁ�O�����]�� !O�'bP ?:}--�T��&���ncl���1݅JZ�Om�%�uM򮾬��%m�kJB��x⦆lB�|��ݿ=� ð�dZI0��xUlV�15E�6��H������G����R;�bC���я��ιǜNԬ�Y�1�K�����r,z����?@O���qF�-��%��FJ.��lb�P�8��P��ế���ܚ%އ�ұp�:JbX�\�:^�uZ;c�s��?�Z���P6��>�UU��}� �t4���J��[Ѫ �K�+j .��Έ��uCd�"IYV�<�Y�y��<��^h���Uںi�0>��\���n����M ?���A�X6����g��
�pU���~�I��G�t����9c�\�a��b������5��*�F��5��
A��H���1��,x���t�n�&����r�fB?�A�h ��*! h.爍vU>q��]�B�$�OI$S>�q�ph��V�;�IQ�'PP4r->��<�F�Q��Mު��'b�Ϋ�j�!�B��QK�0a;�+^�WW�pvd 7Rf�Q���B3���o�Ii[?0�45)�zŧJ��n pE�荷�JO�����C����ϤHj�ԜMѕ��ȴ�<�wT����*o����5"E))�Q�i�ӓ��@y���м]:��wߞ%�?���<���X	Ӿ�#7�u5�qd��)E�>X
ȧ�n�rd�#
�j�Ƭ�p�i��5��3zI��D��i\��z)�B�q|xP�#�T���o�������i�a-I�0$�������E��|�ʸ���8���-TQ����J$�y�gw��aΒ�� "�٢�3�X���j�et�6�=͸���3��>-f�����O�RS�I��wH�
���s�xGT�b:u��S�-6ƞ}-���l�ֶbJԊJ%!�J�0�����G�ϙ2,Y����!e��{b�2b���[s�^�8E�y��"��Ua�3L��v��
��0�@�����2��d����	<�#�`<��0���i 7���ES�x�ETT��'�,�:͙�J�'U�Ǵ�����Ҋ��~p[� ����;��ey���u�fs�#۟{&�H�8W	E�������L�v�s��ٻ,�#"˸����@�Ĉu�Ep� �x}����f�i��>�A�{�_d�.R	Ybi{�:Q(b̥��
6�<�NP���q�z^_�n8��vD��!*]�}22~Qg5'�:DѶ�*f���z��ҥ����lpɇ�@�3�]7'+ �:�n��c����Ҫ�|��Y�X*�2��E0�0*^��*-}p�')[G:��d�/!��c_��~�l��hf�b
���<�휒U�嶣�����ܧjr��Y;e]F=�[,�=��A.�-!�^��N�z��iU�������G�����>3���/�h��F��8Y��T� Sg��0s:s��u���x&'�T �s�7�Y����B�X���J�t�{���{o0�ިt����;\!qk�����{ɨ�}ֵ���D�6�� �f��!������^�83z{8`��x앏��ǵ��q���BEt`^���^gw�됦(�uc������W2WO}&���s�@&���@���6���:p���T#��d?��04�L�Ba���Ui�V"�A^��/����0 y������f���4'B�1&��+�*(�7<�B�N�/�����d�
W�g_im�+`���W*S��![�K�.���hD����f��w(
T��ٌ �����xm;%uҏ�G��<�����Fr�����s36�|��}Ū�M�j�����Ĥ�bM���n���Rr�n������ۛ�/�CZ�8�>��;/��5�<
��4�Bԓ�o���܆��ya.�O�ܕ)�O��᧝�l�w2�O�Дʜ�Z?p�T+T�S{�!֋'``Z#���h��������T,���T�ϕ<cf�z �/˘V��v��>�Č?t~~F��U�8����F(� c���ς�a�LP��=6�ёHԤ�E�ˤ�mb��aCJ�\s�f2��q,��Z��n�/|ob�����\/���e�sH�M�������&ah6�����Aq[6jS(�5Tt�l�"!���!&�#qSM#��p�;�.آ�c��C�����<�f�0l1f����6�#�$��ޚ9���_4V���$"E��_L��hs�'��9�#��!W��BC����%���Ϩ�їcW���ˏN��_6J�FW���q���O\52L�D��/  &|P<��,qgq7LP�?n<ݘ�.�[}�h����$�rY���XL�W)��z�?i���e��/�}�������=lۦ/���،3=ܑ	$���F�=��Q�!�uځ����`]Nlh�b�c�?�T#<�����,m���-	J�����5�`D1<9j=�B�\t��8q��C��9IBX`_$i�!yl��/d4�@�a��A�Q�#LJ�k�G�*���vBpKp]��	i��>���H��ty:��p5�h@������f�s���R��\j��$Oi�!GY�������O��:�EwB�W��4� 2O��H�ys���PJ�8�ZĖ�@��G;}�~�7������Zw3�`7����&Ҿ=�.?����e)�!=��I �Jс�C#��i8�nT�DA��ZQ�D:Y#=䓁�� }���@|�em�m�_���>� t3�,��? ���M�N���c�����m
���
�U�h��H�{����SM�J��|�͓ȏ(�2��J���M���`�P'���1��ųɘ^��`���)l:W�N%�4R�z�n&s#��9���|86!����I:}Wb��@l?bs3��!��*�g���L-�g`���6l^�|�~<´����@-�4v���@� x��s�@G�Lƒ�&�a6�!��l/���D�/Rj[A͝����ʷ|��ir5�Vz�y�k2}:�
�h	���i�����g��-V�'�u;
]aG��λ�$����:�����~ i��Ϣ(-����za\��a��<�4�q�A���Rbwp�����˶cx
��g���B�hd� �՚��K�� �"�T���	�\9���uiRDC�ԾF�F^��������C��n�)|��=���Az�����H�\7ݪH:��q�[�c.gU6�]���0C@h�Ve��DigV�y�~7eiހ$/`Ԇ?B��;L�{8��q��7�[`�j.H��V!�=��D;�%�z�s�����37o���0Qa���N��7�
�i�\�+�s�vU�2_m4��\����x�A�xY���W�S�7$hv�7p�9L�G@v5�wx�ֳbD���"�H�m���s�h/�Y䙁H����k��B������3<҅���'Q������&����� 6�U�iG�ŚI��F���ŔF6*ڑx�㰐W���ei�ys�M���Y"�b��RR��mg"��{���0U�μ��)�+����_��<�������mƖ�i��x�vv�p񕜸uт!٭��:ل�	mro�.`�����zyчz������yJZ�{���������?z&�M���I�7�����Kמ�,�P#��Hzk~�+�a4#�+��A�"{� &B�@�*��w�E��_k��><#�������.�L�[D[z�z�]���օ��g��̴�H�'�Wm�o�(��X�	�!���'pi	W���Y�U�����$����/ǂ&v�mK���nUK�r��m_0#dͨ��:燕(���{ �B�I-�ϫ�ƩbLI�$d,��=�/p� �t4��u)?챭�w�XI���@6�[�	�E�S�6�\B��eU��J���hjC1� +{�6��<K,[
"HE�5a�6^8%u<���?��c]&4�i�l�����.�}$��cS�a����?���g��݉^$�j>N�O��!���2tD?2D�ĕx�N���J�va!���u�j�8%���,�B0<Z�w8G-����y,��cK3Đ������p8�B,;�0�<�8�Ng���nB��j+��s'P���=]��N�,�;��d2W���؛J�[� ��U�>��H�N�����Z���3�	C�s��hK�f!A�a�*��lI�������L`3����2��#�r�z�n���R�:���!�n�Х@l�:�%o�斀��D?�i�$�x�6�Wq��Z���z��nM����b�v���8��h�Nyꭙ#y�����u&w��]:�qbc;C��^i1��G�H�n���&�z�۰�- 4�x" �V��k,��I��N8$����~<��uN�uf?��8X�HV��"���7X�|�4�k�Z^t�2Y�b��s��e��ѯr�� �[��s��'UB ^�s�)���^%~���a(Q���@��VN���%\���:�>[�gX,qF7�L@)�yR��py�LI�,F�a*�Iv��
� �&5ش��LMH�f��e�4Bq��7����Z������>C�Q<c��S�`"ݙqsbk� �K�89���\�ނ�p�e��X
�fN��n5���!Q�Wչ��y�d���S���f܇!N4�C0���'R5�z8=�ܿ� �(�Z[_)��H��6Q�IK����nA�ա��F8אF~�����vA/�! �2$jP��p���x񞼁���S���X��ǝKߘ�����O�5&G�40R9���S-���܁��HiO7~�Y���c~���?��'r|`�1[j{;�	xR)��P�����(����y��O)�䖤�!��7G�߿!1��NE=���2��pbNoX�^�Uq�rg��m<��,�	�c7�ό��[^��.����5QK���	�(Oxmv����_���_������?x�g�0����?r)�H�����0�"'��K��� 䘜ܚEnv��U�O=�-':9�����T{@m�8t[ ��j�1��A����L�c��r�᎓�vr�Jh�a��5�d�C� �$�D�%C�����Z<#�g}wEV�d��J�Y�T���Z8	E.fl�I�᫾P8z޸�m��a���eV�c2��p�:~��ny���M��W�aH����ɲUV�ۖZ	�$��^�!
��6�ϝ�a��A���Vw���!�c~�oC���5F؃�םa�x��C�a��v�~����/�F�|���8�p:��~.]P��a�F�L @Y�<cw,T�H]�� Mե\�9�6�'gt|��屋�4��(��΂6؟!�jo~�T����ԓ�wQ/_\�}�k��y�m����j�{fz�F�*%|Dչ8��I[���sur���h�ږ&��Yz˟׵vg����P�d�3Nd&��@����}��u��h�#���
2��w��#Ma֙����V�L2��V���� �4�+0��$a���l�j<�n�7�2��+�L2WT5[��\9j�����!���m5���3m �M��ǠY:mK��/�qx��
�cwF�*F5��	uHH�[�?��K�\|Q`Z؀���٭��E �����g��z؇���K<�Q���3O�2K���ŗ)T$np�+�Y�4::6ĳu@Z��u��Si�Y���G�hf�BB��$(��G����O�^�'���9�Z��wEz�7���1�O>o�Ѕ߳�3��a����b�v��V��z���V�U��v�Je�'�
�E�wx��o����f��%��o�
����ڦ�����MkU�����`�R�+i�`Dn�Дve��
z�&"{��|3w�i.���D*�G��p��Ip8f�C��,��YwP�OT������b����:F�G��xs5��%1IG�.Y�E�r�
6|w>��z=�;�H�	]J�}�Q�������t�^ ��b�	��WUv��W���m��(O�H-gFx��K����ܘ�']��A<�^q�ؽ�?0|ڮ	���������
��<�;�R��1����iY�Lݚ�:_s��O��wI�:��߅��������*`p��ʠ(^�md;�[bETq� ��;���ϓl~9�h�,6��b�=��H���<�(Li�;"�������fI���;���+0'iw]��I����ֹ7���r�.�L���{K���I���Uh���3�����KB����V�8'���L�x��!�͂��-u�>ݯ���V&p)Pt�"���J��WcY"=�u��V_#��b�xFu#�2�p#Q�
6�>����i�;]�������-RX-�8Ȼ����*�/�#f���C��F�4�"c&\��T�
~�J��	X������M����DgPp�U���C�9)sA*���M�P��oto��:�ƣ�г���x#�a�`ȼ޺6{¾=���5�J�D=482im_�q��[Ie���O��#O��+LrM�W��n%�Nr�ĉ:.J1w"��o�����܄����0��S?�A%��Rs8�`Te觵��|���\m��0�0��æ�0�,[P�V-���̘5���3iB����z$b��&Ӂ5�+�	�l
��w�*�]2�������YBN��K�X�����;ы���k�r{ZP�`r��7;c�»�T�<��Xv\+���(����!�z=s!�
�#T�Ty�ſ��
(��
���y�z?�Qt�Y���죡�R���ޔ5��M�W����0H������l�)��Q��nc�"̍��_���My,ڭ���H����bϢ �e��l�
�����4���2k�iO(uqK	�tD���Bq���i��Ȱ�EX�t�F)y!3��SBYU/�&�u�b��<c~�tVQ��0��+#:=�4�+����P��!��.�5����(6"��<�҈"dN��N7ܮ���:[������1,p��
�y��Ԙ�4iK=
�Z���k��Aߒ=�0C�)#�h�PG�H�p�@Ѡt&�U�K}+�<4�)B�W�(	�T
�,���{��O��e�t>�����7d��|�d2(!�����A3,�QQ=��W^�S�gt��v���l]7�zW��ŕ/#��i�ԭ�2����7��Ӎ3��� sn]�]4�����5^/V���(-�w��O�R���w��1#,�\�~-~:��pSj�r��臫 ���;p�0 ���_�����Z� d	�9�
�|�#"��;a�|���yђ���t<]PN�y��ְW���r_�-���Z��#�աIw�r5�見Z��N���4�}O�}`N`�*n��uH��ѡ�ը����m �`�q����/�=,A
7�*�[]����M��V�ğgߓ6	$��0f�MT9R�sdRs2���W	��ݯ%a�nT�Ł�}�|��7b������~�0;�YܞW�G���OT�qB�=zu���'ϱ/#�@�\h����߸Ci�^�H"��o�1���N.	=���C������;c�lؖ�c���פ@
�HXc�3��6�Ǩs�"�>	n�u�N8x [=m�02�������\������?�T�K�Z�S�*�wd �7�500�q� �+�m�",��>'�=g6$	H����j��6��4����Ś���n��'�)�|����?��PE*&���z4���jc�0rPU`/O�/x\+�+U&;��e�� �4P�%W���J\"�`d#Eqz:Dx�a��K�<�#� /e�9�ʥ��L'MW&A@��ˢ/���%�P;�$�$!>��ޯ^��/�}F&���;�S�O4���]�T����%��@�@�vкYa��JQނ��7���s"���MLѴlj���	c�Ү���F�� ���l��%KT~�tX�M��������q��Ĕ'��t�4A�gF4���^~�Ʉ���ԁ4��6%6f2����PT�˦���goO�l!�^Š�ޮ�z#��"^�<���s�N�ǫ",#[����G:�I`�SW=I���뒚�j����$�s�5�:\l&h���U��f
��;�iM��Q�����wi~N� "�$͗�l�V��*TH]#�_��m�˼g+�	�Kv<ٗ���L����"�%'異��Q����J�%@6��,��k��0Ύ��FH�JU�GR'm�|��VeKN�rʳuѣ^�$D�`֢~[�C%�2�j2�М���jt!�=8���3��#��N�>���y�|������%g�*ŉ����EAΛ�7�m�l��A91k�o���| �V��1g)=��X����H�d��H,����pm�6�FW��Q�����J����>X����N�ϭ+�5Xq*Rk��*�d\1v��Lf6#L���sDC#Ё=��ʣ{ p}ԂQ��I�F}�6nrkW�#/�ke���X�pV�z�����z$�{�~���p���a]�$�5+�H��ȣ�4qӕ��aW:M�����:u~:F��b\�N I���'���U�~�=u��2���85�<U̱�hѸ���"!����v0
8=)m��J�sNA�e�*��e�B������\��mH�4)y��2���Y��%T)�;S�÷���feK8�W"4,/�S���.?�C�s��콀I]e;��3�'%�tV�+6SVBk����-3��኶#|6�w2��8��t���Sc |�I��FRжQ��N�йl�6=)�U����瑖��D��Z�z�G�9��K��1s�Z���֜�&�=}�S2\� �m��<��S9�%�>�(�0��us���f�7E�;M�Q��wQ���B^�@a �d����*�=.����a�q�@W!�=���]��H��砎� Kyb"]+*<��'�����*q��:㔞��27�7l��D|7��SD�,��P?�TY�֙��3�+jY�#_�3�ef�g0WXn��0���k��%��_�����=�
���l�o����ÃbS#�5F��4�40a�e�U��0ft�UW�/K?q�(����q�+&�=��$A# �J�"�8Uòe�˲���N]�y5��7Ӫ�܀t2�p��܉++��9��b���h�j�~�d�2��p��_�dT(�9���]�I!7u8� �|Ep6�jЊ��pB�1 [�)���nh��O����񊘜�RW�H�I-��t!p�i�uӭK�nM��tI{/��� ���d٢�$����j�]�Rj��&�#�ۍn�%bW�u�I)����Aa�4_
��]�熬��@µ��U���:�YЁ?��/�����J��8���D���V{;jhF�Z���2b�׈�>W�/���z�	��#[$C��gF�����&��t�2ş���*�?%xf��!Z�=5qYS�)ǣ�zMXew�c|�0h�q������7k��mfYִP�üsʋ�X�����z�EH�%#��: �R���_�Iڎ<�'���P�|��T�& �З��dXrѫ�m�������P�g���0���f�O�zy@��w�XY��J��H'Ϳz�
;��4����m؆)�+k�<�|4����xp��>����E���޷e�$>C�V�0pw�üK��/�h��� :}U	������&3��k��'.3�O���u�Pͽ��)ZBE3���Z1Vc�`3��:��p(���/`4�J��	o��|!Fn�b�s�Y���?W)ɶ��8�t��ӊ�gY6-?���.q�