��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX����q:�}��>��\�D_/�ܠ1p�n����Ro�*Di��&"��g��D��7I��f- �hE	�9M�P�褆���^Pv�{���P��'����c�p���(_Jb�jiq��k"�r-i-�9u:D�ia�1�9�?�����A�!M���1	���}]i/�h�{)-��!�)�Àq��2Y���1�1튯8���5�YV��uh~�0uZ���m~��ċ�_SK��u��(o#ƨ���&+B�%��`�^ę�H��_�ӮُD����q�U8X�(s���=�#\-��=U��r�1�=�f���^.S��\"�E ق��'o�jA��k�4\���o
�y���fE$�^؉�aVd�pj�7T����T#s������	�|�Y�g�}.Rh/�G^L���ٰj�:hH
��DV�4ʅ�ru�� ����O墪�g�L(��K�11����3p����f�.��&oq���ez0�]ۣ�"%r�%U���脊�Sh�L��YC�{w���@y�����V� �e��Q�*���jf	K�fc�q1�N�m,�A�&��TP#���괮�R�;��yR�J;��.�q)e��{���<x����,g�Tw�	~�!8�e3{������5U��u��� A�6���.E�o�l!�5l�i�|T�SS�M��'���n'B�L�����#o���VhS_�RM��� ���F+3���ØX�������8�������X.P��+Y?��}P�Z�h�!�^{t�s ��<P� zʣ5�IȲ:<�m��4����R��<˅�_�e��YEE+Ɂ��$,�L��B�E���"n9$�k���bc�U�Iui4���(.��WTF���ۘ��]i ���;���#�#���/_܍i�M�o�:g˸�XUo:Td_�9`d�Bp�(��@b��@�,��,��3{ט�KA�z(��&�&q�vtrOp��)�N�lrE��e�2�?�����<�v�9�g��@���uW���m� �K?��*�gʘ�(y�\tī<[��-g)��w�f@�m�����lk'��?���#��V�ȉ��"֗�Yf�I�C��B�ģ�%�T�m� �s:.9�P��n���o�?Eܠp�%/I���$���V�?Z��|sOZgx���:rՕ�,�U '�wN��^*�k�H3siy�7C�M@��TB^�]�'�Jۘ���/��J��Zl�U�
0ly��3GV,�`6��+ݢjZhR�1#و�H����'[�N=�Ja�l�����]�Ω	�����q�n��z�cAd0&���[������)�O���P)�7B*�����E-z[�Z����j��|�	� ���H��Ӎq�T������{#���C�M��r�4*��
����P����� �)TZǹth�g�31�ڂO�ɵC��O�6&���R��p��w���4�t�&k�y����{m�$|�T�ԋ�'��F���͂��ID��\R3�@j��%�܌&P���s�Ƙ��j���t�F��<���["�C)����q����gn��Y�Tez
}+���RL�l���yx��{�� GFZ��И-Gt�w�5L�1l��A�w���f�W$-����%a)K@����mC,��Fg�/Y�n��V{m[RP���"Ά(�hU���	�e�6���U��@q�)Í��&�UJu��پ皎��'�6|0���jǭHja�V��'�[�y�RP3�H9>�(��" ��Y����^`r�#B����C�=o�I�������{�}�BȫJ�Ӆ]���c�o���6�Y��Q�ړ\{(P6��%ˋ�ץ�Dk�"w�h�p�J�؂CXgp��C.q�l�U�P�T�P��\N���F�b~2�Id��j"Cgr��LEʝ��M�M���ko 0&U�N˿�/Gi��rS�Κ]��jK�ou�7!��B̠�Зo<3��0!#�s$�ʟKI 2��F�Z�%qGy��p�h#���Qj�B���K+�珩�Dr�ğ��(wbۚc�zVԋW��B�Aް���pb�˴�[��s�H��r`�%�C!��;�/�} �9�Pr�o�8I#��m�{J��_7�d_�)-sǟ�Hn�Q��#i���52;�*��&��`,�,t/�C� �F�d'΢÷?��������G����Ĳ�W�@�AnP㖾vW�a����e��3��ؠ�JL|���8,���j��f[�͑�~�����D�St�*F:%r#�,6?SC[YYߛq�҂�P��7�I�<��}�2�R��*';�D7)[m�(J��f���s;�z���T�v��3���:�lg��I��Z����*qu�#=v��nS/_��>�mK�у�%~���)���gW�P��}M�P���9��?�("��[!&AzKG�8�j|'����xo�P��L;47�z><����n��M{�t�~Z���4s��S�|���Z�Қ�+�Cyǟ�ś��m�T6(ϛ\M��y����9k-�d��h�f�5.yJ�Q��߯z�J%W9���̔�Ym�E�_z��JA�0-��J1wP�e
��R���'IW�pF��&U���ڢ��V��4��Q1Ww%�QC3.��'�+����]ľ��qa���N|��	��W*%X^w���!����{ɷ1����i`:"(����9����O�_f�6U�OC.��ģ��$q��c�կ1t��j���(f�D&��b���D��u�zLn���M�n�e�r�o�%<9!�Q{�ڽx�s�
E\�X��Y�P~���q⡊h���F����+&+Bs*S�~M5�Y���f��͒��U?�}�3�Bl�{���Ҥ�Ā�[�B����qߧ&LW��!���
:
Pt���`
�4*~*o5듑�x�r�����@��	^86u��dq��X��!�P/�ƺn�˱��\j�� �{�H����8G_��-H����;�Jq�}����$w�+!��nj��HB���r�VfU�5�����2�¦����؆�Pi%�h)}8�y��T��;�f�b�v���G���ޘ�D��>cL~�-;�;U�N܇c��u4�ڵ���(�w3@Bf�����'�5�zR��mk�Ǽ3I��H���:�e���i�g/$,�'u��q�E����'�_�Ghm-��ҵ�2.��8��d���şw����%Ŋ�GW"��~�R�n"oi��#��%�593i��ɰܖh�
�/V��V�J�	��!�Q��S�,I0��8�[�{��M�KϿ<`�v0�B�ga��5Z(����ݐ�����w�6�xY߉J�P�;w�(�=z� �B�:��ȥ��d���{�F�z�9 }U��;ƈƴ�,��������F�b_V��H_S�>�����Íq)��,�{��M�I]K�ɹΏh�̳'�O��&�br��������TJ�|�i>����x��
1S�x���k�ɯ%`�g� ��-��,�9���*����?U�t��ٔ�>�M��>QH�!��,��"[�s-N)�(׬_��/���AjP1.�ז��&L����J,@⭤$�b��\p+R�ذ�R�۴1qv�*S��'�[,#\���NF`����Q�i�["֏SGcL��~�3ܨ�T|��~�#����N�)6	��������2��s�Cx�8B�B��s�
I���'0Ğ�V!E5y�Y�;�$U��1Rd��z��������F���J�	�f�d|H�P�������N4pw��Uf�����q���V�^�G����p��l �:���EQ#��|X����a�p�;���a�L�֠�T�a��U\"��lJ��Li���0��n�����d���%%�9ץZq������t�!Z�MwͷZ�.���_Ѻ��65��um_�p;32��o��QN�S��e6�;;����y��s�5g\42;Y4�GK��p+�5�����We"X_ylL�K�j���)bqyZo{��y?�x����"�ok��V��&��O��p$�q�,�S˧��č�C��Z51�gq�^���W�lձGH���n�Xk��z:�z��_Z�. �b�%�ƹ���s�i�֣��2��X�J8.�Ȓu\(���B�,GM�����T1wߞh��-��p����g��R���S��$W9�G��߆_�� ;ҁ�B�P�Ϡ]�E2̞�ma�dq��7L�)���Zj�oaΏ���W��<��k��		�6�����Q�H�q+�{��C+�x��)��:�Hqk���kUlm!y�J���(�Ój&����2��Pw��[�yhS�H���X>�s八��(j�5���~5:������vY��gº���FX}��A���%�7o y�;���A�~�xw�q*�L�#}$���L<b5#�*����� l�����=���y]����O�E��T�Z�#%�ؖ�U���As��s0:��� ��xUL3�;;�#}�l�sV��-$%���rI,�7�`�-�S��{�$�"9���W����j.2¬��L�<��Z�_BK!��-z�;�"<M8�9���갠�$�f��q2��Hw�!��7��W���ق��O�&>߄�G�	����¿�y��<�P�˷4�����2����	���t��׺�C\5u��&l�M���k;B�Dqq2g]R~���لL�Q�*oW�BQI?�K'[�̶�������Hʺ:P)�[���h�,�|5n����m�G�4(gq-���=�|�7��V������(�I`�t��:�0��\�Ru��^���Bo����Eb�T��Q�89W�c���C�"����F��)G��9��0� 7#�h�|�e���R�i��|P&�n�gw������웫�j�x��#M�����4#W�7�(��\Q��L�T��;^��L��҅	аN�G��V?@)eL�<�oCd�hM\���@����[�c��F�-mqk(ҁl��M�����'���6�d=��쎓�#�ݹ.d�q�PI�В{���ڮ1w�ԯ��P��i��b'�ij�����+0��d�E�q�i�|6�wnk*r1�#��~|��^qh�	)+9�2q��v��{���?P��I<�(�V�����r��/���l0m:�s���s�m'Kt�OלV� ��.� lar�/٭�n��pJ��S͉!hAx�L�5i���Æ��iQns���s��B�.?q��^N�]�7�Ar��P��R�@N\�[���ߟ��Uz�[��������*n�V��+E����j������p�"�Dj��P�����z�bXY��I����#w�W<#��w��X ��eԉ�r��_��������Q˨#�C1���t�:0$h] � �������s���Y�MPs�������L��9�mW{
�I��o[d��(���=�|���~�:��9.	�

���	H��ٙy~���]v�R���99��aT���j�H�ߍ�}�z.2� �q�a�"�Q�,6N��߸1���VuHEZn�R]�G
�a��Ҕt���:�����,��e4'��Q�;�	���н�Eim.�cOL�݋N�f�n f�V]G� T�����*Qe:���;��e�i��\��bd�~�Jkz�S/k�%~?�{/�M�k�:$9�M�6�o�T���[�v\,`���D�K�٠4❕�3��)�_3��c���4ʲ-t�,N#����T4��PǛ���^�v�6	�[lݸ�}�2��Y^�,"ǅ��z�%\���'��Xw5t��M(
EY9��<,ƘJn-��Ҭ�kG�/�eTT7zc�If���8��˞��n�p��e��Y��/7��;QK�d�@��Gͳo��UN�X|i�?Y�a�������aJg�[��P�@&�*õ�5GG����r�;���:Q)J���7`�8C)�����g^����tZ�Đ�����LqLg��.��͑��U/xA�̱��[�_�1Ta�^��N���\�ڙ��>���6yy���8]�_1���q��Z�@!�)���O+j]�,���t���/�$��i��7l�P��n12y댯B�9B�3�uR�CW�V�xp�-�嫲�Z����YdZD���"�ZSc��?y�ԑl�Er��ع�v�$]]O�,�-r��%(=��/DGk�eo7g�)瞍gs��vU�.&|�ۿ��\�9�P4��O,�Ԑ�^Sww�JI�C�p����3X��,չfON������B�O;�U4p��6�pB,�m7�'�oH��NN�Xn�*��y̢��?�%sQ���'�{yU�X���Ƹ���V�"�F�'z��}a͞����{��p�`��;#��6=�ߟgH�T%��0	�2�Aoo�=O���D٩�P�c�p�r��1f��R͞�. �;�ݏ��uuh91��a џ
K�n�a$!��f] �f�����NvR��W������R���K���7W��K�9��I��%������z�a�v�K�x�W�ҼN)Zw���~�R�Fu���?�6�X�i�p��9� ��aZ�ɵ|���al�ղ��ziռS��vo��a�>X;r�5Da��̓;�ۜt��W���w��l�⪶�L�+1���'	d���nr�c܂e�4�6������u�)�wvwh<��w�#���J�74���/`�kS���9/\R��Đ2� νNz���c~�Ȟ� �=�l�W��q�V�]9�g��Ac�e��e��[�M�|��-�ܲ��2��j�A��0�
��8P��kJ��XGL�|r!I�TͤA��U���
�`S���{\b��p,6���H�,���K��)��}4=%}�?������������/W�
i/�pDY�G��9���7o�Z|�g,�!��]C]/·ʅ�v��⠱4�r���(�3��7����g�m��Br!E�ץ��DO�$�5�t���OB�Ȏmժ�i�C�_�2Ie�5��7�����˪��x�V����9݊������	"�=�B�%���?��Y7?�!��)c�鍙�?PiMC�e���6�����*d��h�����K���BN:�C� ȹ|��(�!��=�G}m!n�bz��&<�/��izc����!3��VF�cߔ_��VU1g?lk����6���0]�g��\�+vqӥ���:"H�z����KNF�F �$R`����|�G"1���򚗀pq0=�S����}Ґ)�	��X�l�9��ɽýC̡��(u�b��9.�$ ��(�W��3?�=�@*�T�qo����	�"��jÕW�'J9�������IY	g��O��v]`�����:�Ts���������V���n*��ڬ����>W��j�Ljv��ք%F���#A���ȍiT�W�6�(�����6�|������D'P;.�}o�P��M^�yJC��M��5��N�o�mF�Y�ϐek�Q�<&�Q{�H����r���͊g����/��R�����RgJ��(W�gL<�߇k��P�R��N�I)�X/��K�_�g"��3�;����B?��{UD�Y
��J����Dje���.���eHl�hv��3��p*4�:�9ʝ��P����:�tO!�7��p~)eV�x���I��&+2@,���	h����CDe6�g7s����L0z�[$�e�i�6�>����E�P鹀r+���U�A��W�a��u^�j��5��$ͱХ�W�r�����rɎ+T��,~m�F�m�x�\������1-I
0?�6�n��q,)���kZ_f��I�0PƨOš\>�2�Ƒ�������-�;��$�no�r�3�4	��H[�') nmZh���F���+�P ��+83rփ�ِ�/lH�����C"(vo��s<^����R��9mk��3���3�&�����G���Г���MET��Szd1�(���1���q�|��w'F��)�p|�I�T���M�X�RNf1�m��w+-�J��K��_��C1�'��i�����xrI���R��b�ƪ�c[k]q$��C&MY�e����_���鸁��x��%�$���x��C��뼆��~�	x�]�+��<x�s#�BOjY;���^����F��
�d�O>����&���`��]���֔H|�)c�� d�U�����e�IS�	e�[f�Yx5]t#ng���wս��d����x �1X>�8�=��E�o�s�Bv����G�K��a�.W!��5�n�BI��5�;�#����C����l6e0�U[��z�� ��!��G��O�Tk�EԎWy��,!�?U�p�'��9��K�L:�c
��I`������du8�<���L�C���j�ζ��u06�m{Day��v�i�H�ď$]���1X���Ms����$�m�D�	sV1�1.�MaD X ifL
�E��
P��^��͍��������ڔ<\f�����=��=�c���e�Ԏh�P<�~OV�ү1��[�E4�Z���� �^�|m��j�mUj�ln�nqv��Nї�'A씽��Q?3�Bm��Ooݔ� �r��-=�L�j�o�^�f$݈�����kv��ik8��(�&
u��g��+�zk3�����OG������Hj���3Q��~3ۉ��iu	�R�L
��h�L�h
��Ȗ�x��䙊<��%V�g�m��V�s#d�����`W�m�{��}�����J�W�/��R{,��"��b6I�&����}Ho�r>�J�����oU���,;�����D��;�n_,���z���
W���4��ߎ�³oc��Sn��蔅xcr$!�x��M�v���ո�*��E�R��,S�3Ŷ�R�3�4+�W�4��U�������e�x�%��r�BI.��#/V�j]K'.��c+�	b���]���(j�����$��,�q�w����ju�h�S�����S��j���K�B��9�xӅ��$��*���S��t�mo�L�Q�2 ��M�8�
T|�?��~d�+*�Oה�1q�+eV80��"�ڢ�f_�=�)Tb?S�<��M���L]7wr-��W �\K^�N�_�Ok芒��>g�����_�����E=2�/PsN�Ǟ��%In�Ħ�/ln$X�;�7�.H�W����6s�gI�|�����\pEBy�J�+�Mw_�;����U)���'���<7t��LՖ�����j���>�=�W�m7JP��6���EȰE0�v��Ej�(�m��࢓o�s�������U�)�D�+m�T��ok�f�&{�Έ����Ge}��꫶�s���!��<��Ҽ��Ʊ���7��|���P���w^h{���j%�	_��U�焪O����n�� j�h��_jV��-�o5-W(�w�i)���>����F|)��1R;�������b�JF���������'��`���Q '�N>t�� -#=��pD����Q̯�ujZ`(�/��X6h��ɗ��{�ͧP�=�3�y�5���P?Dx#���Q˶��5Sj�����$��˾i5���6#��d���O]�ۤ4���z����H�e0Q>�����"~���]��1D����6d*4_x��e�Y�o�;KRz�n� d(PR����f��1�O��}�ȶ�WC��Q��Ԓ��_?����[&ѭ���sQ?���ԯ�-ro��/.�yya�0Zf��W�k���W�2[�h��r�����'Q�t61�+�h˕������k��V'��VwEō~��%�]�� %������l
�s��ۤ�Iͅ�16	��4�}!��9q �; )0�kP]Joj�ltc�4z���!V���\��[㞬~��n�!u&2Up�|j|����GQ�G�.9�U����q���j��)Fka�$}����IhJ�(�X�A�O����� Aŧ������A�m�Z���(���`�
P�������d8ϸn��[���ӄr|x^h�g���R��'n�D����&����/o�yS�aQ(%u�
z�$1A����85���Q�8��"}m��Ö�i�Ն�q=3kt�J�Q��ݒ%��A�v�+���" 4e2��&+F$�\W�Pai�yX3��	'>��b�T�_ew��!QҸ���}:��F�9�ξf{u�}�\u���f�Xn�+��9ݣ�,�`�����h�eRB|��i�A�QU�C{�:b� �����j1u���c�d_@Qű�2��
>�_+��;�Ob�=U�-��t#g��k}���3�Ơ@@���k�C�t.P�Z���Y��3g�I���]bQ�/F�f�XT�Gg�[��T�s~V����	BvB}z=��p��UE�[=C�V4�Hp]Bv}��p�+�t�?��I�c�*p�6�.��m1��@uF��>�q�tZ%�\�"	[���9�9D��V� �ժ̽,��̘W�R�LmӰ.c6���i�����\ӥ�xW*
,�zO@Đ��Ɍ}�@:��F�eep^{�4bGq঴�������/u2���{6[�
w�F�JW���S>H��3�I?í�F4A���Z�\l��m*4`�ŚR�G���QlhX9�^^#Wq�:4�!d5���U�i�{\�'%-B�����^��l:G�;x�?���R~k��a��f�\!h���RE(��s�z`���j�NL�eS��.��	�J7�p��"/�y1JԠ�'� y� �a~���>?
�BC=;xv��ȼ@�]�ױ�����Ρ�g��ґGie����F��q�����4�s
\c�\�?>������[Ģ|�/��r�����Q���B��"C����6e}�N�yϯtj�t ������1}DB�����Gr�C�`]X!��(X�9G��=#7���j����sU�	ܠ��)(��f�F��V�-[�;��DFJ�苅�블����gވ�Th)Z�b d�]�:��Z�͵mhw��?�7��}`��Jh�򄈉D��$2*��$��Q_V�A��r�!_t�P��"�$ʦ�V�<�25��<�e��6�ElMh�ķj�U��|