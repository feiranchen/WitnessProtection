��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �	U>��h@��
}c&���`=����nB�&��=��3�&����C�e�4��U�Q3��\�*|��;y���#�՞@4/�6!��	w�A7�).l֬���32#EPڰ}��oS\� �����l{����l��,3���M*�X>`��z*�j,�z����?,i{���W1�	z�X&eY}ZMMt�V�ۃZݪ$ M���֞fZ�cE吕����Yٸޢ�uƬkFbfk�WϙY���\Nt��6��5L>yKVs6��ߥKw��oJ��`�<دӬ� 0w�b���۸8�&��<���g�J���&А�����~���t��ܜ�1iȖT=��k�:/�k`Q��:l��f^F��dZ��kO4�R��%6u|�\�}��IM�<���_���ǀ�*uh�7�R�;�����1���s3�a�z �F//��P��
�5�s'H�zï�q����55���#�-{�V�X�(_��_�w7��y*sO��0h�_W�w�(�2i����]��9��}:=�k����߉�/ �e��r=|h��Ոg���q�g��4M���Ctr��"�54'g��_:��	�N�7K��!5������4E�rc�t�7�8.S���|P=�s̓ߚr�|�R��(�Z������{���4��"�Z���;��	&��s��ѵ�ZV@࿜���^��q�H�p����<�/��j���*pip�S\�����CM8��<;%��Y���i*]�jg���&9@�A�������8三U��T�>�=�e�J��6�5q$�b���(w�W�^ׅ�S�*��������Yk��Z���V�|�h_��"�x�B{�7J\����?����|��r� ^�T���;����.c�K�w���l��;�}E�=Y0��x�'�z�5y�-$6�zr9V���L���ַ��Ҡ��+%ըe�-/m�ʱR~qW�|�#<7rt��{�ՙ�r2�Rj���C�8�?�.V6Q�F���>rܦ��ʁ���g��8�2�}�X4x	ά��Kn=}ϯ��q�j�R�?�£�x����I�
��k=ו	:|�V����#��t��H�`�����[c�׮YX��{5nf&b%f!��I�6G�Ӹ+�u�8�DG�g{�TCɏ((wT=Z�JPy})z��(y��s�	�Vɰ�cɨ��>�����xϴǶ��w����|5f�5�N�9*�$���k�ATo��,���#i��嵝��)n ���)�� 7Y���O��Q�8BK�g��h��U��	+W�[�AǄ����Z�\	��'3䁚BɃذ�'��+��p��T�D�w��l�C�]��c�=7�23�G'L�Ӵ�*M/>9X�=���L��@��:X���HF�k��C�_��eUB����� ��|�<\)e���f��;pz΂nv�8�B�L>��҇�cӢ�e�8n�LہU��6�,��4)�˄��4o��
�O=#�	aKm�Is�ɻ������[F1�����U3^[�Y�(�������E����<�:"ܻ��ƒ;��*�y��~�����[�Bw9�v��3��� �M�/�f�X�@���H������_d��H6�;�F������[U6��۪f�E���'�|����b,�w謟b��9Ռ,p2������ڒ�����G��D���)n�� [:��{�J;��S�ѫ���A8��ytC3WS|�.��"�0L���]�!����*�� ���Hp�=P��42�/vڄE����
wɅ.�eѬk2+s�]����I�DJ��쯒�k��L\ -?�����?5�Ƽf�2^�����QՏ�|IƩ���X��Py�	[&+ٯ<��p�}������b�B��V2�j�YP8�����{�_u���a/�[�kઝ��&�]����JM��+��.�)ܙV?|��E$ֽ�8��qj���7�o��ol�P�s6����e?�bM8��9�;�R�#^ޝ���b���_�ոoHxp�@�~6�[Bo�=��Y�Y�  �Z#�e���YP�B@:����č�,Nb�]SW8���H#�y�ť�"m����ą�� d�����f�8D,�1}��G�]����I�˓]G���|́�GWX8�>�G}�	]���l��Q&�<�6W,�Y��9¶�m:�gl7�R�i2�-�IsOf/2'�Q�?.O�6�M� #� B��t�5�`�$o#��#���5,�Cڑ�%ò1�'!O�M�90m����칓Cp�{�݂E���Ѫ]D�/�a׮��es�t�"�^HB#�PV��(
�!��0� 5g�B�~�ME\&��Z�u|-7Rw�кj�C7���>��t����v��V5(qf�KX�G�S��\�O��a��<�&|:8��'��q�^��z��Hތ�plImJ�*���=�������0c�ġ1�6Ȏ&j�I/�ΐ���JI���+[�j��k��U�ҊA)r�В5̱�6� �������R��-M���P��r�Fع��2N�	��'6�(�wA_���Kq[�fFP�9�!7��4>I[��z��ge˙�F�:�C>���s@�|n��Ŋ(��%�d���~x�B��I�C�?j����W����@X�'�Co��XB���7��R)�5e�D � \3?=إ�fw2���5D�d$@@L�]���xr�r���bB��*��Q�	��l�努}��E�0�h�w������&������U�@��>�`�B'Q)8�<1���k��o�����ߴ���mL;�t��k�<f���gg:>����ܱ�{�X��
\e�����n��R���1���'��Ek��[-��Hg]�S��b/�k��t/����h�-��P��.g�j|�7��.2���1p!\Ϥ�seȻ3�TG�]��b���F}��Kx��L��Ԃ�|����1��O�{e6E})DH����.ly�~�AP�%�3������_$��V�I�="m$�UWѝuL3��a�E�x)�b4=��HR&�Ix�s(��w0H�ax��q7=pcאZ�?��MQ?(,��������G>l���ｴz����^��Q����I�Z���]�V'�����"�R�?.pH=|��;՘4���,N��k,�e;a��ub/d��pU 7���d�iǥ��X'�8tǄo9qf�n�Q�������S��9,l6����mDZo�R����z��h|(fڴJ}��9�~F�p��P��['�yz�ާ���W*��Dw�������{�ȕ�.�93����"Q(�+:�eg���$D߆�����+L)��N�uYĽ�Vi�!�Г^�C}k��2n�3B`ը`�y��`&
���Q�60�����)��r
���p�����ɻ�k��9,�	?���٤�5�Ə�g�o�9��YO�"! �ji�E�`�oAp$=����K�y�x�1�+r��Nhhm�N���* sf~�?i JW��o%;����]v����
��Pr����ٻy��]��0������dѧf���-m5���5����@?��LF�ĩ�����tnP"6׬��fj�����e��#d�����O�m@l���p�I��(K ��H2�W�I@B�qA� (��)=�n0!���~�J����n�	hqj8����Ȋf4h�4��;�O��B"���{ZZ��:J&��?Ε���1��䳔~Cf�`���	Z:P�PtQ7�N�2M�-8��ܤ��(#�_GB�z2�U������]�"#^�v��F�(�G��U�"聁��1�2=�wxC1���ao����߅�t��CJ @��8b	�Tz�'�x��{�wk[��Ty�H3�����믍�	��J�&RۅJ�H��Zd ߕܥŠ�w����lxWM�9��?ܧ瀴{�x��?�\g�B��P/!�3���?8��4mG�E����s�kosѳ�*����O@�z.��}�<���{��?�"�h�����w̦�;��K۫��Z!j�P�M��
̱)��~9�i��8�:c��U6��LW!��w&W�8g(���rb[M;�a�Ec������f�c��۴����v��|S��Ķ��JkԌxggkH����*%��&<�\ׇ��A�u�U��M+�S�Z���l0���_O��V{��  R�x��LN^k��1zh�c��}����C˂�I����ph��X�h��-2��f"�&=I�VX(9MP�:ћ���+v����Hr8�ƻ%�Pa	�g#:O��P�򪓙ȅ%��e�ǁ��감�]�<B��JT��fv���s��}1��e+�_��A&ٷGd{�}kʛ,�0a�\R*c�y6���u	
˿@��\��/��4��h�5(�hab���s �PF<ĉ��P�|7:�e�F���1��}f`��x���X��\V�C��R����H@��n�pK��J�x�3İs^���.�u�Q���vCF���V��*�y{gi�"����cfG]6��A�r���.ɬ0�|x'q���AS�Q$�2���������ʶF��ʸֶ}p��:+���Ĵ�<�NKU�=���D�8ڱ���ʜ	fPH�WXj�M�� `��-@"�Y:ߗ�"�D�c�#�	��_������A�5��Bm���cl� +�6������#�c�3��kX4z_�?�:�;߲�"����^���9�N�T��+v��fWzQ��8-C���y1�TϠ+�WUD�&���D��l�'ٴG!r&��
��7��ǂ�?׋��䨌����Tc3 ~z8�a�k�n&=ށ������v�i���T}.������i�+�K֙HoT��Jm�[otm��Ȉ����f!�塨����lP�&oA��*�Y���Vnr�:�KO�':w&/9�|S����ЈYަ���UX���S��}�F<)���� �������3M�h"������mūNX��&I{�b���_%�Ůk����=������؍Mr��[T�<;�H]c�/���0]�? 牋жr�:6v�[��>�/bd�s���&4QV]�D�5H;,�J7��LQc ���8�]凶��_a$B�ӻ^��t�8�L�Df�f�չk��иYo�L���$L24�ߦ���b����K)Q�����s"�(d����lh�t	�Kal!"p�]s^2�_��_ivˀRߏU/�'C-�����	�9�v��9�qi9U?�	�؀l��ɭ15i�Â�H�	Ǆ�p�(C�����CEn��ʬ�wt�3մ[e�Kƫ�=Z��'����k�8�����\��l��m��ui/7(�a����ՅH_o�Ƒ���Ѽ��=Ƅ%)E�=����&T��X}.ȡ��T������}Pru�w�p�y��ފ�m��Tof�Z�[P����Z����-}+�G1�����o�6��}����z�4d^�\���ȵ��sy�j�f>�_S1?M�Z���QV�-��Z��4_��ԭ�WV���A�h�qu��[��q��ͅ+�v�F�a���ťA��0�nE���<���CwH/X߸$J�X��ý�E��͍Q7���.*�����I�d�x:'f8�	�I�@Y���v?ƠX��XfZ��'#DH_�4�\�+ L�&r?��4zP�HBǮ���W��&bW� ��A,"}�\R��#�N-�X~�(�\�6�N��!
�6�}f�A|IR�a�ߋq�6��:D~�����&u{�؃i��F���	լ��b>��QOg�DW���>×MP�H'w����	�-I(�P�9������Q�_ ?U�_��!�۵Im�ڠ�7�q�}!e���n�>�Cb�{';��/4�ԫ��śܭ%!�c l����(��'��_��'z��3�l0Y�$Hz[��Z���fE�����	,����^W��:��w�AA��X�	���O��c���Jg)M:�k�{���.�" �_&?�]0c,�l����Z�����6&FD�n! �i�I���0`�;�4���,,ke=�J���$F�
���9�;�u|����	�wW��9ˋ�}@�3z5WڬU3�ӭ�����AMg���A+�I�Lsa��7�Zb;�|χ_��j5>�n��$f� y̔Ҹ�rg��n_��{_�ؘ�FܺM׫��*��b6����N���^uÌm�bt�q\��V�<���&��F<$�`ʶ��ْ7�./ڮKQ^��lPi�q�rh-e�r;�\�Z~�uT1?%%�P�u�x�z7ma�$o/잌�by�_Դ�w�����`���.���-	[��K����,�D���}���⃳ <q%cHN�aWPT��;� o �7`1��4���8%UK؛�U�{�l��J�d_�#Pk+O�J"�Ƹ��:�x7kb*	����q?��ټ� ���HZ�Z�f�,��?�2��Y�B�.�$g�D��1V!<=�<�J�xH�Sܧ���F�K���6J�@�~��i�Lr��xZw�,fiE��ܤ(�3�b_l�,sT9#7~>���Yנ��������>�밁�,�u�U!O��-�N�o��;�3z(_��w�k��ls��z��M�^��Q6q,��n��;��V�i����E>2�T.��^c��)�a%!��/�+f,�zhS�v�zW����@R��ޠ��x���zc; {�y'�������e�h��X�ж��sM�)rs�����-ZٔX�:��{�@Y�����=�s[ZNs���>+���(��w)}��D��8r|œ�TkץsV���
��?XA);�{$W##�=L#l���tD|�:�{��7�eC]s�\���{�e�c���i�ۄa,��BiIgS>,%-������(�gw�����qE�n��`� ��R��p*`�R�[���3�za��F�nV�V<�U ��h,��&g~ˆ\���wk�>t��ƀ ��6+�z��=��Pwi(��̘���y|�)���Mbx8	�J�[�S�����4y^�k����_�2�"}�B��wp���D�y1U8=p��Y�r
��ol�}m��M�L,��ח�b�G�GsT��������r喳�q����T���l�Q�a3�pKXA%�:�?Vg2�
G��P�Zؙ�1�m�:���7-'E2�
3�(�$W:x��?��R���}:��8�vV�s �@p���!v�z�"������۶�R����B ���a����b��d��9f"�74�P�
g��-�z��b�.�p}���qQ�����fӛ����f�ץ�������V��4�*���=�h��+Ěz��Eկ�Z�gܓ�����x���9�V�B��c�}�I|J�z���vJ֋ݛ<�:g{?l�}.`��Eڇ3��\3	&g������㡒�QΤ��1ϧC3�0(( br!�Ցp깐��������T���2 �x�ODi���O��+k ��:������{�H�G�ȓ��IYسQf�$:�x���z$��I���7J�gHʅ_9��4��-*T����D�s�x 6���_nD��O�����ek]ܞz%���?5?&]�V��=�eI ����,��HZ��܌���(a�͑&��M���2��*~፴On���ꟾ8���.���&��'w�J�Y��%�Ԯ���8��\�돟sյ;(�t���-�|�.5̩�.p�<xc�op��x%��oa�Q��驈l��ˢ�Ġ���
%��4���J��;U�;,i+g�)���<��y���eFQ��e&u	p�����]�$�
oI_��PN���&���<"���\{�d�%s�n�/�bᬻ���
2��-�mu�,LŶT�-���*�KgF�� ���*N�]��l#5vqV^̨���{L��ob#� *��:�̛V���㔁�S�L�c/�`P�������e�(�OKb��ыu��w$�(D�p֜65y�a�'i%��+@c� <1���[v��s���rSS=m��u�,Ņo3^'
Ŝ�0&��cY�p��r���o�"�2�	�a(����Ox�Ih�E<9m8/�g�����9�D}�$D�h:b0`Z����p9>�f8��d�����4��֧O�P��UVw\�5^�
���݉�m>.a��|��5夬���A��m3��kK�K���R����5x��ʮZ=���D)@%`�gey��P���8 ���Y�?�Q�f�"H��96�i�T��&�fME��[�E�'�I^��ҫD"Iʴl\#�}>��#�\��:d[�����QO����u�Dҹ����X�y�$;�r^U����v�zhT�:cs%g\�|^���c"�PI٩jq��,E���X���2Hbyq7?��~��k���u��Y�j�eⶖ,�N��z�ļ���n��;�Qq��b�����+%��{��1���g��Ne�A���96ICH��k���{�n��:~��(x��H�|)a'N�z�їsg�36GD��l������;Q�.���a�g���{�i��,�L�mj[,�<�[�8����F2BZ���G������Q+v��'P�$����C:z!և@����aVѶ����F���|-̂V[[��bVC�m9�����8[�"�����z�wZ��ZRVv��-$�ȴ2���b	�'�k��W����>�ɽ�l�v9r�\h�4�W5��D��A:�n3���sVl���pc��BT��"�����gW��ۤ�Z)�Dv��;]��ۑ�p���Kgq��
����lW�W����tI���� �s@�#��Q5�����[-��A�$^_�4Z[���V�m�/�w�o��xp�mZ1���%$bcg�/��"�˺���&��ɽ�C��M����aQs�~�%�K]6(D �C�1�� ~���Ϩ���]�٬hO_�a�'R���&n����pn�]w��M!>�]f	`�V˄��x�!FW�nɠ=�_I�0�X>!�!F �r�z�ù�Q �A=�CV�����R��xbkg��9�B�#�10�0�R.f->:j�n5��7J8_�j�+���o>���.G�pn��kʼr1���v�o�'�:C�=��3����	$iW��+��28�j�!�]԰$n��}䔮�#ʆ�?���ɠ{D��(׸Qg�MFP����y9�D�� �E���g[���qZ���oN�	o���uIĤ.i�kj�=ɺ6����c���R&1@M��1��͸W���V�8��-J	�N�8JA��띑�Fw.\����2�p�BE]��(�A���>P6^��P|��l���%1>��d�h�n����^��	���J��j��z�P�[���9@�3پ���	3k�y;�p�V�����=�Y������X]�^8Dz�Ԩ�DT}�?��O���bH��/_�qk ߰�g����v\�X�?0o��	�;J�:�a/�!��x����s>=T*����O܀Nq[$��C�_�����g�,��*V� +� Ѯ�&��3��3�XӢ�����( �6eWn�4q7�nS��3�C��CXmX�N�W;g+	#�~/J󉙫~	� ��Uc�-1:���0I�TQ�KZ��P2;�[�K/s4��2nC����n9l�W��\�c1���W�F'�ϧRY��'�T�*e�����9�k:�M`��J�� ��|91�Fc�k���@#II��v�9�\ڱ�E��ԛ��o�'�p�3L���;#�;�#���+R��i{���k7�豞o �drv�	qM�(����[��y?�"S��N���8���%�nU�3���:�a=�|�����J��ݼ8�X�9rϓ�K����v\��x�H�i�=k6�}�����u�Y�5����Z�=g27��A0Q��܆j�t�g��	ij�LGJ9�B>��$��P�=vpr�$��EU%�)�e�
�r~3������}����]�3Rp�[�HU�����qѽ�2q��8�����[]�!�7���<`a�䒱zHo�>�+��.��>
}D 3=�����5�S���ʟ��N�R+��`)�3��36N�Y�,t!*��I��3@�5Ԩ�[��(���yj�p����b�'gp���,!��b����QÝ13�?Y�i���2�iU��i�ԿT4Y ��;"W ��ԠW2������)b�\B���F�";�v���WK5�!#��3�=�W��e��PhfY�TmWH��q�i���CS>�J���Lt7ɼ�������Zy�F�Я��){�R�o����E����tAB���n	"��rr��k��x74���R]���?��a�5��?"�O�b������j>}^'���A,K��y9��s�g�\Pk�c�t��x+˝�����ﵴ�{�mfs�*O�Lݗ=�t��גQxI�����A$���t]I�����6��ß��D>@gF>�W�5��B~���*���I��/�� Q�Y7�T�[����i���>P�R�;/k�P"X)È�����������*~ٿr��zJ�� M)V���t#r9�O��7½S5r#�z�, D�bKg:c�@d�]�8�ka9x0D���Ǣ��w�~'BB-�uR�������҈c¦�V[e9�ct�浵�����^�P"gϼ��6:|7��!�K�bp%��0�@������):��V�}m(an��^�� �K�B�%�C�`�t2@\ U]�m�s�|�$�����@�4�YN��O+�e~_�>�z*���N�)3]����w{�߾&D_�����4M��;�V5�M����6P�ޞ��?+t�^�&��)��~|�GBG����7��NRx4Pv��pXX���	N\~K�"A)w(�0Ԍ=r���o�<msPz���������r��0���↚�� C�*�{�bQy�8v��F��{��]ڥ</4rh'),A5c��!CdP�(W�X	�E�p������F�/�Gs��N(�0��v}".<@Y����8�I;��Lw�A8T0  S�3Q���m�D��L�5w[��bIkZ��Y�����;�
���~#¤<_��sj{+�$˙��9ep���l�>#�&{.[PP�����YV#� ��Y@�3&j�[�n��l`�8�<t�Ԉ�H=������5!�'Pk�]y
���A;���c�9���X 1a{�5k_�����:)� �G���[�Y�c�ow��u�f�� �R�T�����$�yÅ��V@b�v_��AeJ]wr�>�dQ�E����S�Y��]i�U!���s�`z@�A�P�������N%EsJ�6��S�)����:+��^J%���Z��R�!���iC����;���@�g�*��+ �mQ��A�\H1��G�pvD�v����s��)5d��jjR�Z"���oz;м8�!��\"Q����i+=��]ߠ���
L���L+
�;_�M|D�F1��d�5���=(�Vh�
� .}\I�6��0Z.�/�X��ZR�-9�����Ě6�r�E;�m������"��u��ű���/;<��EJ�Ta@�p�.�H���JQ5��ll���i�v�,��<$�1pjwû��Ea��L���qڮ�PD����F�� ��*��?$rm"S�͘f����/j��:t�g�� ���
D�X�J�'��:���3N�;-�be�y+�a�p2r������(�0-��Fz���)r|&��;����H"�>��R�J[���c��u��H�f�Ec&K���mHZb�|[u�2�Q0��L{ã�0����8�Zd�<�>��Ϩ���S+��
rGA���aF���e�.����P;\��<��\n�,���'=�*('�� Z�y�n���g��E�(���k�K�	{�ᣰ�����HN:�0_�>N��1!)�g�$Y�G��#�]�{ƹ���gʴ<��w�\���X�o�4X��ތO���>@Hp]�Z���Z����no[:�E���b|~��ρ�������Eٔ��7d���zU��0T�ſ���m��0"5>���N�>�~��d�`�3	/�գg��,1Ö��X'��U�E�1�	QD��}gt�Vl�o��K�-^*���Ȁq��c��h�<��c^},�Eۖ0U#سEl%<{����Bj��ͼ���j}&� ��P/�����k�ǡ��t���o?[���6���&m�2���)]��A>����[+o���8���n�P#?��uK���4���,��`���$��W<���q˧:����i�S~vS;)����!wMw=՞Y���[ϻ9������m{*ĹV�`�^�nFt�K�_7�h����h��q�L������%��/s�s}T!��w`�}��ș��p��s��f���2�C\���ä�vf���,^G�Η���լ�"L�����BX{I8�M�ʽ��6{̡�c�Y!��>͂w�P1Y'Ql�[102������ߐ��Zc�؟ޛ�+��������*x�_�����H+�%|�t�Ȇ /�~�AG�	�Ń�~�o�G>je8�Z����L�Y�n���W�`�ꚺ3�)&-r*��g=Kb>:����Op��morq�?��ˁD��O���gDZ�����o����*��]qKk�لa}��L���B�����Dx4����g�+1U���ЂB�_�&��6����M]3h}�x�Q�AfY|�lN���*F�A��+N��n�D���پO��ъ���?�T�|�J	s���E���@A�r��]SW��;M��>�Q.��<�H�oʽaa �S~��˄�+0J1Wx��DI�}Y�ϓ�d¥�(�����̀�:�A�ӵD�<�=��w�_������|j��n:������Y�� j�����O�oD@֓� ��D��k�7T��6 � |�s�I����/���:(1���f�]�&83��l?���;Vx<����k�FF�)j��aA�%L�]�EXio#��H{}R��GI͘�
[���ڂ�A?����pQ�������Q�@@ ��x���)Sj���2.@��	?fћ�I�4��R��5}+�l�Tȑ�� ���O���������3�u�E7L�_#^�{������ߕ)qNO
-�n�0�"��/ �N�zy0�/�����L�h|�����(ٖ��E���������{<�zT��4���9	�[i��%c:�`^�����L�����0�����E�'�+Z~[�tZM��܃k�����0b���֦��9����H���-1<n.�W̔UPե�Zzj�IS�����~��08T+��i�(���Nȑ�G5������c�`*�,�W�;�>f�ˏ���� ּ ��E���������T^�<��C-�\���w�VL��^�rfN	x⋃���Ħ%RKK����}��d�(p��8h�k�����( �����;{e��D
��3�aP�8<�u�6�*���п���� ȼ�a��&�{Ɋ݂�3ҁ�l��q�ܶ\�8�������5�<�V��bz�{�J�w�g�6%��׉q��A�ve�'p�f������5걲�=ӱ�OIE��� ͏�۲"�ӽ����w��, !+�7K���,�Q�@�E�S޽���yR��~���l���6�PӷlC�1?0J���[��G��N��c rr�ݪ;��L #?{�jx��	�s�4P�P��U��!72��sx*y2�����`]�d�&ei�)� [H�}Cg6���^�Y��v/����
����ux�Ҏo"buD�·���(���	�m+V�������jt;�TG��"�U�iƈ��Ya	������Q�I��{�w����N]ߊ����H�9vm�2�Ά7��4W��X����s,��t��Oy�^�����X����NoԸ ��KclH�1��Pm�Mn����1r?�c�W�FK�Ij���_	>Z�!��~��i����O��Bt)���
0q)�Ov�H��|W��̱$�5���R�Eԝ��YݦtU�A4��|�hjD���;��?��w��*3�Y�G�҇�S�M4�I6�B^*�}���PP�~jd���`�l	�^��5"GT\7�c��OO�{�F0rhh�.�Xs5�	�h�
q���']�!�~E@���7M�m ֻV�;�;Z��ZؙX��-���t0/ns��j��x����[����_��(#
�8����/� { Hki)d.��m7sp����m�G�^eka��UE��Rgf:&�`8���c��$�������à��`�v�J-��L���S�58Hv�󑙥W��Q|����y�q3M��Ҙ�h O�Y�����{�8���U෩�z�&ٙ*x��#6o������A��\�*�]��H6s�ѯ�@sA���hPV.���O)S �1��*	T{�ͣƉ��B��՛�\�z�V��Ҷ�6F|2�+��X�UTM�eBsk�CHu�:����]��]���?�5ZB9�l;���Q����>)p'g�LqO�@�L��R,@�6gؿhU�F�J)�Q^��>�&�V`Q��+������SF����;�W1�G/��B񄟅&�e���ƙ|�Z,f�֗�\+���U`R�4Ȧ�|���]�\@-e�z"H��Jv�_�_��bl_ޮ�E�����;Jd`�ٞ���6$��f��{�����1pM�gj-�����z*k�������� �B����L���x]�� �Ɵ։���j��|����: �R����2M;�(��hÔ�Ȓ�O?���!��e2�f�������]���H�7���z��6Yस��.$���P�����|k���n��\Qc��F�Y[�Y{���+��7�K�'L�'�#��ʵ%������ǡ��bh�E]��R�dD6¦�R���u���&h��s�1���Ye��8����#c�i
y8�Q�b�� ���Q�~�IO�b�#vg����ɜ�@V�����K\{=�Wu��_0w	ɥG^���o��c��y'J�����K}���%1���&2����$=�㺚�����0�h�؊5�q+��P�K����bՐl)���u�.Ū��{W�=�9�~X/2�m}��ˀ�Ϛ2�W��	�6}=��S��
�:�D.��}�9S�M@�7'��CBP��]�	�Q�(�E��r�璱w�1.q�Q�N蜗�#m�K�/?�G	u�W��&�)��q_��ͅ�`�&��(c�l	�#WǮB{�8~�F�x��	�sS���>M���ɠ&:X���ytRQӓހ��!Y�%]�s��ۻ�O4M��|��*=jS#���q	W��f��b�+��;b��Aŕ���ղ{��&fh�U��?W
��z��ִ\J9�ϋsUC(8�^;�'�43��|���wۮ�����sT���|G��{�+���s=�n37T��s���8D�Q��j�r�1�"U^s��b�n�,L�p�=��D�՟?�/�c�\��(�Ex�ꃌ��y���u�� [!7M�b��k�S�d�R�X�ҹj���T�=��>��$R�ע>� �
�c7lz;������X%0@hA�����{|�85��cS:U����ߥu�4�{�:�D�	�Yq9!˄q�v��%�5�O���I���==^���O�-��ͮ�&��]�P��&ǧן$�f�PT0�D9�D�E;�s^����!�P�TB����6���	��M�i�^���E�{���W�<�N�.�΂�=��rG�`��=�4��.�է��B^N@N�0㗲�k�Hi��_�{Ú}Ǻ|��ˌզ��U�0,*��]��BVP^�Z��ެ+��:�9��(,�N�Q|*��h�Fb��]-˭2��{�[tq���n�f*pz���F�+������>?�&X1�`��6T�.�M��պ�4���g���I|��4Uf��7�r��"�C��aȭ�L	br�����+4�3���r��w�BaxK��n��zu�/d���++�Ic{S�f���1�o/�Ub&9	޾�5�����/ҍ���y��M,�ɴ?64�qV����;���R8������2	)����%X�ıQ�N��o��`L���J���V��d�< ����*|*�Q�8��Ō�0{�h���p����}�?��?�8�K�,�
Ѱ٠w���r�,w�uz��φ۩@db�F�W%'J�k�)�E[�6�[, ���O���JW�������e$�=9�ʔ�l�}E����\�$nZ�S�Ҋ�
�çL��c���"[N����a�鄧"��=�s�^��XO!�uY+��>�j�q���#	7��-�?Xxd59�o"-�I�?�������R;Z7�=�'a��W�R���a�߈G��I �d�my��~J.�89��6G��v��HX�7J1|<�C"X��=e}������ ���faI�e��\��s�9B�:��H���y�/?���l�o�ɏ�:��ɬ�@ޚ�[f��1+���Է�&�Vj"� ��&��Q�H`�W>jZY~�����_�%�Q�M�h}x�A5�
HJT w
��O4�~�ް`�K�HQ��,M�I����ή���>�piˀD��H����4Ұ:��˖vM8�>�� ���d<���抔Ǝ����-9W�:�� ��)v��>���{ޛ���hh�
0<F�z>��mTD!���8PO>��;Z���>��	��d@�����B��PPv��S�^{r?'w��T��e[=r{!���{|T��9(l�mc��Ð��^����>/o
]���ɨ���l��jB4�ܟ-GE<v-�6�w\��ɯ����+(�n���'_�~��;�}WG��8N�&�j��*�Ζ�HJ������j0�tLNMA�zu�������FE4�4����2�>O�EGj�zyL���CJ�˪oI`r���(���o�E�&����(L2+�/�({Fm�e���e�`̵�j��âC�D%�p]:��c�'���拷"����EX�������+������YY��P�E��}���ELDk6P�g�z�$�+L��l踰�q�q߹��ۚwz ����D���%7j��t�	+��ݼymE������Y��G�p���m!����'k��}��05�e�|Ń95�o*�a�꾄4UwP.B�/΋=</R�k��*�H��6�����xuV|׋���`6��>��m�ʏ�Mb~ń�O����q�A����Pl��4~������6��iȗ�\?�&�����/P2�q6f����ԑ��'�$�ԇ���qBh���rꁢs�In�p �Ejb�/����_�F�᪊Cm|	C�Ji�:�c���ފ�;b���=!�R��ܾ� `��̓!��u�'P�bz�==�A`�VhJk�S
f��{�Ͷ�]M��'����~���Yаt�e*<��*=��x.v�sB��[��Ɨ�x�:X6E�.{�	�~���`퐵�D�ɉ�ì�]+ݕ?1j��_��m��w2 F�m�X�B0H�da�}m�Hٟ
,}�p����Qɨ��x#)D��,�T` nF���*
���-a~EH�:IB�����}�W�X�qX_8ԍdY5��\H��Ei�u6;^���5�mD��D/�rV�%�
�����
����!_��[4,��U��҂���N_Jg8� ��Q'k��������B�Py�S��bD�b���R���69��@�8��ϵ��ڊS����7Vn��t����Y�q��U���ή��1l�Ӓ˄�a���ջ���+�>��}����E&^-vE4������O�d,ĩ��ɟ��p�7n����2�
��bX΅�ᆳ�03$i���7��ӿ���&���K�=�%�h������{~C�:���G򥧪�!�m�1.^�j�2���ǫQ��62̹嗕U�>���[x�#�����x�C�v�G��-	����pa�ճ�9��%M�8vN{��֥��q5�q��K7�^�Bg-������Qd
�)�U��%�*�k�F���u��٥8\^S~Ӻ��o��-��i�L��b=��I�����q�^���j�I)Gy������C���1�N%otOVȫ����!�������{���;$�C|�YAR�u�m��R3�6b�:����=�
��;L-��F���ZR,7?��_��C�''�/��] j��WaR�8ZE���͉U� ���h����K�eS�2�p��+L辚S�f���5*��r�5g�3\O:6��t!4��
����b�Wغ#[��XU~�c5�J��:��ۥ3hY�W�YL�a�#�zk�	78
3m� G��m����._�q28-�p~	C�L�W�w��%n&�A�Qn(�/��5�9-���1�gR�0@5gN˸�d����`��9R/!�d�N5H��;��:񇕐�U��ϙ��aƢ $l|����̠¤��n��aǆ��� �z�H4�2���g���lf� Q����B��8>gەK����0949󭓮N��M~�/��G<�䝉	դ<W�EA�[�J��x����NcYwou��8J3�u�i�d"�c�םW6���������8�r����mEl"^ɬr�������7+���`o
C���\r���S�ݦg<���+���0�JI�3nr��Q��IK���'J�tXP's�G�2����J���+"l�����$#R�����*����W����<��L��-R�����OY&�NӦu}�X<iQ{㺜!h�	��0���CNޮ��U�Y8)�P��\�Gw�k듦	��(��Ve3�v��]t�G�J���fYt8;�sD��i_G}6J�a����^Փ�4�3���}p1�V��#����>�~�k`�"���#?\N �
Ж^)ޣ���ɗx�\rc�F�����
�C%E���I�kn�9�Q�trgi�B��`�'>ٙ��5<磡��~���Rdm��Kp��K�/Tى��u 0�\����C\y�����]�<9�+�C� 	��S0�yG����뷌5�#���vSu�E6v��ϥ좥kؕ�*�??�<ݲ���_�c�"��(���2\��Ի�4|܋*�翈d�+�x��L�1�[�j��ru8S��UG����@9�����HA��=�����*�~��<�C��������$��wA�����S�xɮ����.5<�ol^m����%m=�^�-��;�o��<�G����"uT�cYZ��YV��K?��}O�Db@ �(�g4�).�~��,�tɋ���U5����b��_w��sk3lBl�������+�d�f�M�s<�|���P����d3�ϯ(�(�c�'�A�v=�F0�"�[������ȁ9�SB��P��!��]���*ٌr5���_����/���Ӆ�"L���,�����~�F������y�m��O���/v�][b2pN���%)�"���a���6��������5ׁ�mB^:�U}�Gxv�N�#:k�MC�'C����+�K����6\���ImE�7f��o[wʯ��#U?
F{�ݜm��"��0v����ԧ���QRH�GXʄ�kQ�=�`� ���b��]�2^O���%bA� ��@--颳l�g�t����a��V�Y,j���I+�f�{^Bv�	e�3nF�B�΂T�<�0�4�v�M�/p�b�B���R ��H� U���7��q�d�\o�O�Cd�H =�Rl���I�=�e��)g�2��o�
)[	|uH���g�~ʛqe�'�� ٗ�s�W��W��������J�.�\�H^	��q^��|&H)�e�)�9þ��
��nk��ME��0���%@{6)�e`Z%������pl
�����P��x:30K弃|d�L3qO;b����ߧh6�.����%hz��?;��%���{w��1d�aK�U����֍�2� ఁ��x�z� ��{�ߧ���'��1����k�q�㨪���#H0H��y����xl�s��	��e��m���x��9�C�4�_��K���׹A^�tP�ϵ��+��U�V4�qMο�^Wj�&�Ż�S\�^�<����F��j�Ɉũ�|oϒ�$;�����MJT���u曻�>�r��[�=���fG���9�Oɐ��Ts�!��3���O*N�(QT�Uгsn h�zC�B%[�ƑQ�M����@X�A.h���:�i��qt���{t��t�� B aNb�y;kP�#����Nd�9�QS6�Xs|�>+)U����aښ�\E�,J��d�"���DX	���(�D2�
#,]s)�;�O)�a����:���=�w"��/�5�o|1���7ɄPO\At�6N+�̓�dq���{��ZJ�bj�E�4�s��Q�Ů�<'&���E��,lv9-8T�ՑǺ���UI�n���y�E�YFku��Cwy�r�D&Q^E;�]pd����z�,C�+\��-d��`��!N1��������(ܯy�����/�gK��gG����(��l�]u�݆~ꇨ0�[���;U��E{&��S��5Pm�[)
��C� ��㠦P���w���B%J�����a�lb婬E�v���+��QA�$�|�"O�d�jW��^\*m�)A�^�G?e���B��b�:�X^��&�O|�W�Xii�Jn���C4	����EwQ���l��vu��K��C�	g�k}��jhv���GՄZY6��Xd�p~=q�r>�=6l��G���V����gٖ,8.,V�����X���䘵�����
9�"L(�`�_v�#�����4����;���D:���-�x�+��$�{���ͤ!�kt�W����J�������N��qD٥.�%��`%��綯�Q���3�[��~.��_͛y����f�HY-8�HB���<��jv���f?���H������X��xʇ�cِo�'��>�$]Ǖ���@b8�E�{�~)�<Niµ;ً"BX�a'<hJ��~$�'0s�Fn�/�K�tH<�z<��=�O�W���'3�m����Ƣ/U��o��w{!��1g/�Qގ� �6�OU�����U ��J���|�Dk�Wޟ��@j���������R7���qM4�:�~�VG�єd��k���|y�{E�{�;'T����=���  G�19y����]�8NQ��_^���yS�r'�>ԁG��hJrzT�i:�V�R����/k ���_S��0�
9���|��w�\H��b(�j�pJ˸��qs����*��(ү�������8�n��+����%�E���t��vR�GO��4pު�C�4I�� �#�!ĭc�k��ngq@޶RLjh�]s�v��f��]]5�z�ȗf��7�(ܼ*U�b�vS(+��ӽ$���0�ܧ���Yw���Pi�mT�UC�|+�����YqވP���ˏ�Y����Q��b�J��C�^��=W[�lͯ����Ñyb�ĘeD���Si�-������u����W�z�N����gM����
!�9�M�Q�:�x�㒔ar�V#U�`2܏}���1�$��x��n�$���6ьM�-�a�(��0�?ƬA� _�M�V,�\��ϐ���sio��h������.6Q�D>l�{9��=n5��d���t4pj�*����ty�ڳ{��Y�ٞ2^�wч�ڣ#sd��Ǝ�5؛>�9%�y�6�-~U�Vr�?��n�<E(y/��f k���=�M
>�)U���M�̓�%�eL�[��& ��������cTZg�רM��V�5���y{]n"Y�w�p��=���8#Њ��$�L
����	�r_���7Y+�t�Oxc��V͠�Z��K*�}�]��HIS�!�=�k\�af!11v�l_+ou=&�lW��O��@��O���/x�Uܩx�Ij�#͐�$�"�O��O0c�Ln��x�+F}�}�ɉDɾ�N]���P��X)�<@0��ȿ!w{7$M���4E3u�Mq�=
l��Apz�U|���=�Q�i��J�{J)G��͌���]��=��(���=WՆ�K��앵7�)Ú�EO�Y5|���j-l�ݶ���
	���r�e=Q�p�'TB����M�0��p.K �c��j�=~ c�7��	��ǀp�1|yi\�pùk�uj7�!��APN;У7v2�M����H2=һ����Nv�+�o̬w��a;�zC�`�7�"��i�9�)���n'�<�{),h��ɓ�o�u�i먰4ڹ��$�5b�{�����!�|q��ɓ��=�3p��W�#.�Q��/��(���0���<�y�NG~��T!q�y�i��\