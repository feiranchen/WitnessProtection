��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�o��ȃ|s�Pq��T�����u����. 0�fb1�30�M����m��l|�VoƅG)Ϳ�&���d�d��vf���K��ev��a,�Q�Ra9.�r��ƿ+]��ܘi�1_%��qt£~x2.��ķ!)�P{��Qhj1!p$�N�m�NAj�ur�N��F��h8UC{�A���[d�j_������ThM�����X�����ʨ�����-�U)۾GOL�s4�/�
WL'���	�!�8��3E8v����~��/��3��,��6b�͖�o���������0���a	f{k�D�gEn�]�%�sý��w7[��&�f�T�ś\���x��%N�!�HE9څ��Bi1�����Jz���$ٜ���	�A�FS�T`+"C��%��d]�	?s#�j��_=L���FvM/���92"qF�����h���h��Y������><�@BhԆ�'�]�lY"�7�#5<�Z���ә媀~L����R
ŗ�bC�\�~b�!����jDuخ�a+��HW�J��F�j�`�l��jm6Y�l2���E��c���)aɔ�J��c�Yuһ�!�����:ڸ)�9HAc��Mzee�5�� �]ԑq9x+���<�����T�KZ�I|���M3���H]����Ú!�Sl���ة[���L��?�j�My�� �h
�̴�|��Y|(WĶԄ�g�%�tWM�>{��eVV��<���;�d�W�ؤp�8�NJ�'���Z5������A%H���:J,���U��C�?��1�~�G�0w��<�2<n�խ�j���64���FZ�l�l~�	��Υ��9�x�w�hI�rx~)x�l�a�%ک~|�����{+����	,[��ɒ�#��, ���Z���k��q/��Y��d�g7�ﮙ������_���u%�Z��g�(�`qG�3��%t8�H?�[�]�sW�ܨ�ftt�θ��G|��e'������}��1j��J�Ԍ��_�8��r$R��7Е��aS����U���GE����.ŀ�pZ^;�N6f�GM��6�>��V��1��`����"���q��r�Z��	!���*&Y�#�T��{`8�K����~�Bd��O�g���wZ$��~�c]�f+~�KD� >��>t��&=�it�U!gVEzTᡢ�|@+��K��"g��_c)�<�c`�O��O'�P�y����Z���!���mY��kt�2'E|��p���(�p`��l��u%����H{��փ��,$C�o�׿�P�ˉ����NεP���A��9���)��aó�3�j�sU�H���,U��B�� �3�W*�����&~Kp��Q�ѐ�sBD~�p�da�}���m�җ
�H�p7���%Bo|=&����{��NOFiL*��FA�ɤI >��q� �S��k�	 :g7�,�	5oĹ�aډ��Z�N�HsaC��T�e\����<��P��YF�V��$7Yъ����w���wҭ�e�k	�c��Iݔ��+�n�_wB�|yW'�H�Hj���8�huѳn��y��ņ�hC��j8��:��/������e�#������ a��O��:�	$�5%;	������E�i'�}��|Ox���9F����!o��ޣ��Ǔå7, u�~����U�"M#C�3�_P��;O��_�z�ud:�-_�cs�骤��(`&{dMD�B��-���=�4���ǃQ{����{O\����'���S��j ���p�/M�0�= ���� `�n�����7�=����_:;��'��>>���Uĥ�b��f1tZz�iX�G�|T!#��.^!��_�#�:����h�L$S~�區�� ��]ʦ�g�>�v1�w_�����rE�"~P��y�p�n,���	��s1�Z7N��Q�#�$�;8��D�҅tLش��lz����1����B�/}���R���ɠa��{���OS\����:)f�`��N �Į,��)��q��G;���^k�D����������_���(�SJ͸�":�R�q�m6�Y<�{f'����Mn�w�ky��>#�<�j�O���*�ݎB�.P� �}�J(�#V�ea�Hȡ�l�!pc�}�Í�r��!x�I%x$9�t�)0�ưD�"C9/��:�Y�8����Ene5�'ݙY���j�͕���=ɓ�0��pd}�|q�dT1��#�j������;����ٰ��'�4n�����*
8f�
8���+��p��Y��˻W��N5~��Rq�t7�r���y�gf�7��� қd?D�^3/�[�7�e�P�!�qn1D1�ȍRӠ4�H������Ai�\��]�7�.�AԬ��������u�k���*V4& J��T�Sx�n0��o�f�D3��C�0�k}���p�q�(v�=���0.r3ڥ�� L���,DQB���,D���a�!OO]�^�K��ɗ���)rtE��NK�ӄ ݡ�:v*o�˦�ƿ�<9�q�M�� nUJ�l헏����G�/4����y��Q��۾�A�N9"�P�u�
���B�1�`�����,�`&&�{�Ըq�ʛ��=�9;������{6"v����`�H��$%�5��y�gp=�8�#�7	s�:����/������
T��V�-0��e8��Xi8YRR~�␅��\��ա�c'|�W�"�VD����z�W��� ��&,�x�ɿʿw�j�Z�	�|RV�s���>��4ݷ���|Kw����5�+�i�-H0&J�GmLd=�M(0�?{�{5|��H�ͳu�3?a�D����s����[��6=�C�A���"z�b�)����� `pU����^(Vh�F�k}���s<(Xz��)��u������4���!�U�1��:��)i. �W@�+�n.���_�o6�J�-�,{��`I
y4�qBfu]$��aT���y�B���$"�{򽀛A~��3v\(��}8Q�zN�Iǵ��Ҧ���hY덑>���&�"8�VC��Oe|$%�y�X�K�|qߞJ;��J�7�Qk� ~�9̈́2HO�Š�˘�Z]�
�8��Hx5̄KJQ��sS�`Ҿ���XX�͠��r�U�Ve��y�ޞ�$�)���$=9�U���<�/.��æ N|�{��j�eP���Xn�O.� ��v��P, �n�%�c`5.��]��Uݖa��xx�N�BU�I�N�������[*x_fJ"_��:F��5��7PӔ���M�xX�o����xu�둌���9F'2'�)~9�в�^�$62"�Nn4��EG�G*U7Y'TN_(Z�U�`.~��v)��b�V�p�%J��&�M�)0��Ƀ�U���J�;��H��eF~���Σ��$;d�ۘ#���Ȼ��Y`J� ����:���0��*_�"Z�����n����<�棽��+���0˥}�0�F���w[��z�UT��x�� �G����i�h�P.#Q��� �udR�M�C�������NS�@@�
Â*��o�88J�A�Ȥ�.6:�~+�EM��^�J��D��L���X�=s �8����}	�C �Ăݧ��o�m"�F�/ �ՠ����Ce	g;x�lp����z�o�P�C/g�PN(*a��׊/��+���C}�y���z�xCbqn[��RQE����p�N���(Vvس�>��E~��x��џ�Tl4i*�/uCcK�&������}SK 2e$YCcI���ǎك+/N8HbM�+(�O�{�N�3�y��\���;Ls�$�c�鰠E�9pYэ��:�vʑՃ�  �.�����
 ��y�Si%:�)��V���k�i����_�6z�������X�Q3)��#ݲ�a��s������kR�Տ����ܕ��1�����Gs�^��DI��ܥ������W�h7��Vڡ�M��q�]�Jj�S��ŏzWBL�iyr�1�3g%�6��X��gn���xz��� 8� �_1l�o
����-"�a�C���]n	���73?9<d;{�d���v ��Z5Da�c���f)�N���)�YX�>����ݯ3�kF��,XO��Kq�ǂ�A��� ��/����K��Y�)�AGp��/U�zxL3wq�K�0�i��� *��ΥSk�EKL�e\@�n�g$6Tj�í�b�IT`�/��N��R�ģ7����/ZO$�5�|2�`q�_�lِ����6oˡ`��$R-�%���p8,5�2w>�m4|��\Y�C�V*<�A�Isb�Q6���ܗ�L��7���&�����.�,�tk6���,(�I/�Q�t�/4���AǷzӻ' K4�����~v=���=��+m@8|ߺǯE�eQ̓��S������Ȍl�����=�fe��F�ʀ�װ{ԁ�KAc#uE��/�J;>#fV�RB��) R�DgZ�a��lD�C��/zF,�������{��oFK<-�d�n�R?3�Uo��Kf?~=j��7�:��v�@�������T��P'y;�����	���[����"_U>�=���wq6r��[�DOf�>�G.�PE�������x���si!�{%#�X��n/J�yڐ�ܩ��pE4�����&�㰳��xt)������;�PYii�p\��40������mlŒ���}��K$�RqR�����w�����1���md-��[��~޵�fW&�`�� ����_F�13�8v��-+7�4-M�I�!o�کg'B�������޳Z�Z����L�!�(��I��y+4}�ɯaI���	����P\V�{yrȵ�8f����m�S��gl��]\SP��&�-�v�.FZ�@�i�۟2n�1EVW�11=�g}XH��y�w��"E�6i~VJ�T��j�9�[�j�$IX�꽨������g��>�% �\\��:��e9�伙�5���'�T����,n5��Ͱnay;ﹼ4�n���~`�'�_�,��j��I��/xƭP�����?P��o��bT�t�Ѽ����h%�e���l�H|`�ݴ	_qȖz5��u ����ݢn.u%G��nf����"B����B��=Mp��l�ݦA��,d���k��(M���+��~�q�sƁe]/�M�o"F�V��[zWP6�����L;���FR)�*If݄]A��*�\*v^i2y�D�Jy��u��C�=i|��������hE��!�>�6<��T�W�����B;���'���n������8Z-��X��,��	l$�Pļ����]��8��%|�� cJdS��B�Uo�π*]<�Gv�ƄJ����2�Dp�h6G�yy���N����Ơ`����5�C�p���r���\�c��'��f#*��i6"�$�e�q��W苙�:u�Ԡ��J�{��;[ɔ��Y]��)�f�o��`!�}��2�HβO��B�*Ȩm�%1��;������W�����"f�i��no���-s6�a����ޅ����Og���,�:��y���>�	�&sţ�;�������̗B���@������<P�t���9�tRy�8��Ǹc��LXO��A��^G�+Ԧ�9��M^��1�����U=���^��R���	l ����ᖮ	�&b�Y�j�Nѩ���o�_Z���z<��r�r�j/Tz@HX RS�T��F�%��`!�Ib�}���ir�kΒ�F�I�L�ǳ�s[�1�8���L4�`8�ˑ�?|V&��Åܮ��/�8:�#�N^a �Up���d�cD)��ր��p�~��d,�l��	Y�[甉���D�n#���J�����[�ׄ�����W��#�hT�b��,����c ΅دW/pM�+\���g@��6��/�W4���HD�Y0��!I�,��t����+�F�_ݶ�,E�X�QaP4<����۶�±�g퀬!�����O��h���3���Y�<w�Msւ����{�I`��
ӯ�KC�rǨ;�NáF�3X�G��N�PN�m���.uI��T4�c�����M`9>�P۸��a�G<��R��x��%�2cJZ��cs��D:G����Q0t���ȳ��G[K��J�yt\H��PD���}�}1���(�of��Kq�ѫ�$������6�lǒ�qV������(���tb�TS�"��y�f�H	bׄ=�#
�	aC�C�o_�4��фj�i�`��e��g��[����bj�c�z*��G����cn��L:�iAqK}�_$�������_6 �Ay ��Pot����XA_L���Y�}��7�R	o�$�������ra�>um�_�1'�z)��H�;���s��X]<7&�̆���0,h�q�נ]S���2��t�w�ӓ�-�ނ��Vu��BևriP��%0y��g@�}��ہ�jyǠ�/c��*��\_.��_�j��5#W�iqy�J���<8`��Z[���h�C���x�Չgn�B�%\��S0���d��݉Y��L)��=6�J7'�cH�����HWs�W 9�,�J���Xs\�)�۩{��y΍�.V�v"�B2��yW���nx�ſW ��Y]S���̻UHޟ�89���k-?	V��W�P����t\��;/��M}_��j��J2����_�7����
wg8ʗ���x� ǅ?�2V��	u�)���ֲ7D���?N�{CP�@?�[���p���9�/�����X�T��{�l�