��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��M���h"��;��ږ��[`���u����b�gt7URVSStγ"�SD��_��WM%����$�c��d]��q�$&�T�*��"^a��OR�|���k�j�����螈�	m�o�ݨ`��?$Uw��HH�4�����XA�,�لK%E=�tiL&n�8��l��HZ�F�SX̲1B.JG��T�v_[ �A��F�,�t�eΞ�ď������L�E����Uڶ�6ji�Jp�D���Gލ)͋#�"���I�
1���0n���~�����0��Ԫ�y|ܠJ��TH�a����#i�G�#Ѭ�9��k��1��8'�mW�p� �uh�ty<=�H���*=��Uc�/:�ǽ�	��v-�ܪ�r6���b�5��k�-L	8�-�;L�$O)��Y��A��]!e��Yy�ˀ�>rݕ0���ӓI;h&`9T��*_�VR7�k=�k�NݖS���Oq�E��y�����?|�	�	\�X��D�"�n{Ԛ�U�,�G<�::�4k�貆�a��hI�)%^6�r^'D���j�/�S}k��CM�i���&d�k���ć:ϢL��T�d`6�E9Id��0�NeP���e^Ψ�I�{���˹9ʦ�w	˻@fn�E��Q��M�E��.����Zp�5���t���A�n�� 2��5��SD���ZSɯ�R�N�t��L�ng�ѩ�oy� ��$�g�sL����C�E�>�TAB��3����A���-ɂ��� in�7:���1W�b`Wy�x��}� ��Oh˖ �[��Y�x�]���+&�HR��M�� ����W�1�|����It�j0�lI���m�"�Wp��I	,��#O(�aA~�<�P�[+�>��L!k|����4����%1��f��t�Y�*����+w�
jE;?��<6�#�d��<,�,12?�����'�j�6�|��>?P7�L�JP�fz 腍\@���؃%[��L������~�!:|3��pB3J�������&n��uWX;H�����F�ܿ��䞾�C�f�1pYzI_��j�|W ,�6L2+l�V�Ŝ}�xcG�x#�ǆz�6�Hpo���E�n&^��fum�g�˞M��5�ٯC���g��_��`B�ɋ�;�И��h!�X��-�~"��mIa���mk.�,�� Jc�fA�	�:��;~h�����韸��^~����dM�2h|Sc����_|�L�/[�Ox�ʹY��K��Ĕ���\���7��aX�;g��)�P�f��A�H|�3"�� �ګ{�v�EE����3�	�����~	$;c>��p� �	�ІzV����X D$
�g��8{�d�GnS��E�n�W�-�2m���-�F	���f�		����IS�_�󠮭�Ok!%,�E��1g�H���+_�[e��a�=�D=Ƥ>Q�a`�8M��U���n��,���~hL���1{@,�h�7M�w�Bo�idM����W�V��:fE�s����Ϫ��y����2�D�Hq�����P즹Zx?c!���Đ
t�r�c��>���!s��C7B�2d堥�����j<��G�m��D�W��)�?��)�Q�v�+�����J�S�w�V���T��� �a:�P��^�h�J�Q��c�'к�cwI[���}U�Dn�\��+�6-%�@�+�1��UБb��h���O{@5co@A$��r��^�i1"�K�[r.IN���<Nq�����'kaO�" 7�w��D�&��5����
�S�2��OG��J�-Eq��Sݮ�?�ΰ�/I<� ?��bC�8mX1�|v��T��_A�?F;?.���b��n�X2
'���Z߮_K�W�#�P������7�YObT��6�ˤ�) k�B��Nd4#�I�Tn�:n0�
=+��B����(��S�4@��}�(n1��_�:E�Hh�
�!�����0T�WD��*/�=g�-�۟2���T����G��V�.3uA7+n\]�Y$4�+��T�7 `��؄H��c��.��KK�;��P����B�2F��I�S��duL�C���S�P@?���K����ܣ�?|j#g�t�i?]��**