��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�O��?A~'�m��ʜ�w�3+��F�D��7�Pդ�#%Yt�u �	�����&��ؽ^T�sc���_B�`���Q�Em�*uK���on������d��}�B<&;�7~6��K��Q��
����Iy�f@�9��m�T�S���g����A;��[���_�g�Hkgɜ뱳�y����K��1ħ�':l��	�0��t]�:#c`�]��5���U�E�,wZ>I��	.xګp�W�y!�ž��J�[��n̻9|3�	��d,����u�-���|���MB��^j��'FD1�ojtI����`ܑ4�,`3���-�?���
��)��,�f§f�p�[a�
��Az&�Nb(��F�񩎘���K<<g��i?�3�;�! u��Qe����	ۨ?-M�=W�/���K �\p�<����Q)��@P�O$>Y��j��=	yôK���,}ؖ�PŇy� �C�5�H")�=�߳`�;�ئY�����A5|��Z��Q+g;��F����N������}ga�`1�?�=(
	b�~��狍���a�|w��~be �A �9�.-�����2ǲ߿.�+�}08M�H��9�$dY.�O��!���h�������%P�O�Jj�qX���2F�9�2a�h��:J��)�.LCx-�An#���UP�+��N�;j��6-r1B���-��nP�������ދ��yY�߳��p7s����LP_.�1Ȕ-���%N��)s�������?x+�ٚLh_��҂ae�k�m���E=�)�����^T�>��-X �I�owq��³>G�������Q&��^@��)B�*��q�Gf����
�Eۗ�@G7i���\�ySǞ����70��E�U��賄����7��dj=��v�ѥ'�z��KS$GRa��������g�T ��I��W)�^��[BI��;" �%4"��sF#�F�_Uk��-�X4�^�!�Tj�kbt���e���?�(�`&B4����� �_G /�E�<(�̫*�zl[\`夓�+�����q�B\���h�.w��;���~k�t)��[X��F4D�á���a+���z��\[��_Όr!�u��0p�{�X8�ۍ�@��K%�J�͊H�s�Ȍ_`Cz�p���+~w0!iY�p�i���_�3=DB�
5D^����*�J7�R  ��(�^�GY\,�\U�MG�D���oj�R"[�H!�N�+�\I&DA�j����nH���Zf���s "a�;��aZ{ͧ��h�T'��,������8W�`�JъeD:Ow�Q�z��Dei֚ع� �������~,�
`��OOjj����wu\�5�/��`�wd�>��������-;t�!8ə���)���Ak �"��K��e�.�^H=�p�[,�Uפ�4!w���4s�Q����s��u/պ:X��mB5��nJ'*#zN�$<�$�p���%�n�x�� ��(d�b��|����e���~g�o�$Pv���*T�w�iC��6}��L��^v>��v'�А�V���_' 4Z�a�TG����n�LF�,u�1J�p�d��%�Ȋ��m�>өj$�.槤���,4C��,�H����1Q2��(����\�H�G%'�I+�R�Tϸ�����0���C�1d�c ��n5D���!�-;���6q3��YqxZfN��n�Tř1��!��;m������j�*x�����<f�2!��EL�ͭW�0B&��Ss�3����;�MG NHc
�7�V-�k�R�X�� t9�*�n	1�I�e�����Y�=&x>����S�8��^l��J��Њ�).�k�x�ǽ��UR�;��|*^ a�;B|����ȕ�Y;�������v!��?�)+�r.�gU�y�0�j�*�`	ф[��m�ZW�:2?���[�-������Qk����/�Ze~绦1�̇5��ߚ.����Pc[�yzx �𡽔��HE��]�id:3�6��� ���^��J';��H҂\��oN���l>�nOʺ��kz�GS3�[�U�00��ZB���(�U�j��_7 qlH���N�TX��[V9Y|�]P��ςV�N^v��\M6����T��Ly!F{��0Њ��UF�r�R�>G=S#0U�D���k�$|������4#���<�鷄6���nNl��r��-K��(_!9�$n��ז�=���%i�X&֦��u� ��;)H���!�b(H&��o�Nj����i��T�ӊ*��@7n�Ux>a_��w(vݠ��&��DfV^T��h�&���wd%��;�q��(;�*8���wΠ��,�`�\�G�Lr��ʘ�ޗ�+���;���G��q�'v��~ k��nK|�i��V���P�����ۣրP�	�k�m_�:!�[�۶Z� � �I��r�$T+��}��g9����w�u|v���)�7Qf��F�K,����O�攸��Q���#m]�z�^#7�c�ۆ�A�SgƜ둻_��Br���gx��g0��Ϳ�P��5T
 [�3�d!���iY�D�|!u9�k:&˔#�J$��9�kn(�1��3��<-w�����une��X��3˷q��x��ʟa[�7?~]B~T��������lg�8(�� �-^d�X��8x`	���}��w�'�YT�H�m}�(G!�<�\��u�'��g�J���+a��������I��h訶ɜܑ�O�a��M�P�h���?W:�0	|�>�[��px�>AR���5���v�ҕRًV;��rX�:�鹷�K����ܽ���-�(߃_N�K�j�t�V4ܷX
ޓ�ݐ���u��}q|u�2#u��8%H���},����F�x��N�F?�Z2� 7°��t���<��k��d�"�_!4��{���K�	,3Y.�v�3�!��D�`ξGPS ��n�?��8��Nc�hʤe*7���oYN\_���z V���>"�>�0]&G�)�B2����L	��d�A+�ޞ���t�I��bf����J�������eT��K3WzYYU}�gR���q]��<�J;���y=K��k�����7��������u!\��~�R���*��EѼIH�[V�klZœW9FVK���\��V	��e���v���<dEf}<�C���>�XSr	w["�U������2�ǀM@K������>�\Q��͹�Q�̀b����[Z[e R��s�3E\��+3-S�`䱾)b�
���)��Q�'*Z���=&C����GYn��B������ZJ6i$����Wh1�^�,��M�0�׆ |��P*�kbh�'_�h���W��-2��eh�;��?��VDY1��	��En������kKTk��<q�V�=5��_�� ܍�����!td�9F)���x�����X?�[u�w���J�pvLc�pL��X��8�	�����9P�z��@���~�2�m��N�� +��S2�KV�>��d%u"{0!v�����[�eM���yQu�-������!İ�pkhY�,0��ޛ���b'?���G�P�R6��N�|��$<��i2=p����$Zzk�{�~��w8z�#1v+�C�:��#���e6'h��qDXc�ZeP�.H-���	�~���6��ҏ��@|��v1^�Od��:��,��%BB��g�n�iSJ����6�ՠ��t�.V}��Rj��F+D�s�}�*��Ps*8蝁iR�X���h��D�%/��2�o�7�Y���v{N�KW�3���,:8z��n�R��eUR⹡q�3"<�2��+4V0���?�ܞ�tb���Gg�Yi�����B��.%���F�P�9'�@��&�Z�}�o�����7�&�V|Dঊ7b��e�U����@��e��v��,���q�HL-r�n����g�^�"�"��g�A��β���ģ}KzǨ�Z[����U��ؓ��ݹx��]��v�NfN-�����"�1��}Vd^β��%FM�P��[���ƟN[-|��K/C�0�"& ����V���UL;�'7�@�:��=�f xDu�X6C�A�*���z����B�vr3�jRζD)'J�r+*M���R���)S���P!A�����Ђ~[����K���� �l���6r�����<�z�C�S�Xw.��)<|���_�۸:W�����8`<Ic��_s)�����S�HV� z�o�Ó$N͔��fmp�m��O�փ��$�Y��4!𾗸&��/?�l	ص�aͻNjg���� ��iB!/�\ǕgwR�2.VY�g��6 K���A�]|Ci�@�#ʭ��}���T��ni�z��+A)��V�ێ��i�ȶ�Ij�^;(p%0i:ܐc"�nu�&��(&��7 vv��c����#����ԁ=��0���.Q��Qr������]�Ye!�0�bE{��
4�;���)�������H��f)s�E���F@)L�!�h'"PG�R1�s�&
���]�F�"$F�nGR�J�s7�
Mk�2`�A�w��(�y�dԱR�*=��ZZ����d� �K�b��{�O��V��m�l�����Bk]�Ȁ�yD�X�Sƣ��8��:d8�ѵHEŋe^-&o�e��5�h]:>�*������#{�J�~���LT���t]����$́t{S�g��Zh����';��z\ �a5��V�����&�|n����$}���p�Ogc�LZ銟�߿W�.[O�����v������"`����#|�swD-���Q�J�ΠS��GPޡj��=���J0a�$�M!E�	~�%�^��F��������u$�����(*�`Tc�6���G��qSnT�m͏�4�l��y�b�
��f8�3����]ֽ�G�e���x�^F�R�������&3o��Y���@���Z��2�=1��v|^-�m(�8�U�  @a��!NU%�Ȝ���1_�g�P�XRt����	��&�� TM�