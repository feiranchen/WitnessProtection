��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I��P�/ǻ�9�-��Q�4I�-~@i!�L ~�5i�u���bJ�g՚�G�j�b[��Dپ�mN���_0�>����E�kJ]���V����M����ɀA{��7+�e��ʝ�1^��|�/:��X��I��4s�,�,�k��HTY)�6�D�g�ȵ�4޵i�1NB!M�����Ǌ�V�,Ɋ[�.��l#������ܝk��.}��^sQ�i�>o�����)�Mo&����F���8}|A�C�F��!�������/÷:�r�BY�PY��i-h�#MnW!|���ƴ�`���}�&wK�m���Og��?'�#o+��:�-��+����#��^�Z�J��?�Zޙ�T�t�v�F�03���a�6j�_r~U�\J.x<�E��l����_`���U-t��p �D�޵��?�5��<�=��t�S#�8U(�'ʙTS_C�ԀAEg�/�d�ZA���6\�����~����lQ��%��V64���"�e�5�;w�9杣�u*�ޜ{�&��eh��u  �#YO~.�{�f�� -���kg�=D*M�o��@)��ν�Gc�{��?�ܪ�2ocX��C���[����̴!����3E3`2M�냞n]��)
�}z	�`�H�>�)f�B_f�Wc�C�,����0e�%!!��$�#x�'7 ����u�c1>B,XX�T4�ңZ��A�ܼ�]�Q���i]@�tF�B	|2 ��>��K)o����|HNQ����_��▕��Yi�ےq��[�Ѭ�|�(���*�w���UX~���J�	�M�p�G����6��0eVQ*D���4��!n�����Z�v|@%u�ƽ� ��b̚h��6��u!� FƖ��rr���!힪M��9�)S���[�j��G^)
z�,�
'�|=�R<��M�@���tXp������HJ�m'�c
0��| 5��Ѡ�R�����ij��M9��b�����}n�QU�&���2/\m~��]��K�X�T�]<��� ��i�7��Ƅ*�u6�ǫN`l'����f��9��g�qv���:*ѰǬ�u���?-؊ �0R�2��g	��(8�y01�B}N��	l�$����E�Y�O���n《k~m��yW?��\Yi{z�U���h
�AwŻ�����EL�`��TJ���p��n!P.@wۡ��jY6�?/����nΔ��o�0z�y�vEt�5A��Gy�<��`V_�!E���Ryv�p�]4���-�~3CP�ϐ�4좤TF�
>V�b��}�2<׌��pw�z<Tdm��f���SĨNV�u��t���:&^�I��JvA�ʨ�SK=�g�A���.,�WG����P�Ɲtd>�~�9O�.�ҍE.��o#'r���C��� �_��(:���}�_��c�?����}ۜ��D�ѹ�h�V���YDN�\q9+�F�