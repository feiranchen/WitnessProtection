��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T�K�b�;���ʄ�/r�S���pd�͚g3���q�a�)��s
Ѕ�<�sl�Ƅk���ƽY�����xw�ԏ�L�J�������L��J��1�'��̦"k�����~����g��/]i��Ed��"A����y^��k��%�_��&�V��A�l�u�ݭ�d�l[`�+�8'�/��i���~朙:�Qڑ�`i@b�^ |�]��ӗH�T;J���1��� ��O����r�vH���Y��aL���v/�EG*��CO�<�@%�~�
B�,c���F�L�7-�S�W�������s�k��Hl�=*
W"�[T&�
t!r��T���Wn��_kY�.��1�
l��U���D��e?p�����i�����4꾴���`u�U�s�!m�6t�3�R$�=ݬ��~����ՔJ!�i� �����]��n���-�)f.�!�u[����m�!�c[�"Ѽ��"M ��*��
'��A�Ln��,�ZP������]Hz�ق̄8G^}<y�]Vb�xRm�R�%�R�@"�}�8Z�i�e�R%�5��#���`�sn"X#�����r'�S��M8Բ�qRJ.��sw%���שԶ��Wk|:������O���U�8�DX�X�{x'�ڀ2�elN&���KQF������6�k�g�B@�k�)0���������e�x��٩Z��Z(:��l�x�R����Q��Ȝ6\��������"}2r/Nlfd�����
��8�/��=$.;q4@��~�x��?K6} 8�ΩX�in6�Z����ׄџ08���y7���tA��~���^�4�������$��X�ߝB���O�����w蔎ښ�Į[Ejy E���4��{�׮az��5�-�w��Y{3����
�#�-����0�q���@��=���P����Fę�����P�̌�q��8,9���y�1j.2�O��tE���:�d����=ǈ��˞G��W	�gNT九x��z�f�ifnj��<ix;Q��M����2�At�I4�o<|:���s_Gl ��8�nVA��'�H�L�i�t l��B7�	;�%*Di�&٣�T3�<�H����̽����gC)��:����N�!�C��D'�9��g�d����8������P�h���#Ӎ]7�[u����,(�aL�\�J Z[�Ļ����Z���^��z�Q��z`�����ƓL^3J%����`lI#R�5o-$�R\!=`!���5��4���c�F4�.(A
�f�h��wJ@��d�Ţv��Ғ[���_��@A�R�k���g���s����Fr�-�-���
�E�]��� o��E?�%���*/�E�rrrk�����u���A
�N~|1�*�(C\�1���S�W�%!�hP=�~;�R��bئ���u�Ė�d�;PQ�NY�����k�-wC�mQV`7��5�p�	d��Ce2G��Y��y�b����\.n��
��K����v�!,ڽZγ�7���j���ib�դ^eޚ"�ɦ{?r�B�����>-�e�ζCPN�nx�bDH31gZ��p�&��r�'*���!3�&���-����9�ftػ�9����)��F	�zq� �X]����0sn��q��S����DG�Ьd�0���v����Fgʿ�,z޲>��x��t��T��$��k\���>�J�ȓ�!�yuc�Sm�e���z$m�>�\�
��f�*�h�x��� ����y�k� ���;>)�K�M��.�{Y]oY�&�(���æSK։a��s�\e��`�1�����0b�k���dݥgnG�as�r��!���Hn����IŁ�=kh�_:�1�O�O~R&m����J5f΃����6���#�bu���)�=�J�E�x-���`��qϪ�����Ԫ�aG�Z�[�5��Zv�
G1��h9	�MfB�;o���X�'C�����.,���fN|���,����B��R�_jk���+�"��j]_H^��ͽ��1�)u-��E&��Dn�Vl����_f}��I5�"�h52�Mr�nļݗw|̗[ӥ�Ev��Ad%��Q�<͋K�^vbjN���|x(����
���.w3O��?q�m�)�:gO���#
�6Q2j,oH�
�^lzG�d+�c'�'��Z!x�(8\�j, ��C���f��(.ȿ1�h� ��e:K,Q�lʲ%���6a��T��]`�-�>#�<�	�����d�+���ؘ��������_^D�}����LE��4W���ƛ�S)�����Xӊz�#�0H�#�qN:P�?��q���G�p�ċ=_�xh�~���u�e������>��'�!l���XT�%��Y/��:���u���T�AO�&��]'��R�:�j`L0Gi���}V�0�fY����6g ��%7��<']�)�Lh�8E��v�-)�o&K<�{�-�y��g��q�mɾ�Q_�J~��Fع���.��3�f���B^����A)�)$��ǎj�OT��
��uB>f���ɰ�W�'a��tS	��]�?��'�����d�(���gt��� �4���酷ӄd(<��px����b�[�曗sB[I���֯i��:�Y�h�E����Jx]Q>�רm�81�N&Ù0˱��!\�(����g���R����^7o�Q�8�� �c�P���������x#���Jg��u�w屙K6��7�f�$�.�d�q�n���ρ�5��}Cm%Hy�$K�BG.|�Om.[�@����L�Ak���+Fa�:vi��+	�u��u|1`Ad�����o��.���S���1!0�m��7�L[+�c�M��>�Ԫ�ɰs|���ޖ������������L�ژk^�s�B7R��P<th&�p�+���e*]�6��L�_F�y_���]��0�VK/���	�:eQ�<������3���N��I�"|�vlVt������xl�#\�����r�y��E�C6ت���n��6RU���^=��v���#���BB�=�;�Z��.n��l���|?1�z�� ��0����(	�Uʪ�|�I�c5=��L���5���k@�|���c����2�Fs�o�nFGl���:��i�G��޹sqi�ͯ�������g >`���JZ�,��Iy��xiC�|��B9�f�g#�WCب�Y�%��Y�z��xi��⮬	���w�iYeX��L��H�J�D0��%�U�^VV�e,p��Z)UkH���P}��զ�y��q����GtR?�z�����5�
��+��,;F_��Њ�7U$>Y�	��17�oVg�shҾOF��
���~��.#7>)c#|y��o�M)�_�T���>e;�*���ѠH�"���������C�,�1D�JT���m�&'�g\��,j�gp�Ԇm��k�,a��ve�Y��*�@�Q+�dY���� �����Q�*���/�ݘ���r84)>s���'��/��c`F������г�̌5 �+��62������b���8P]Ho��xZ'U#0!�)��������9�w�~~/󯳧(��E$�C���� �l�S�X^s�����Ǯ����\�Ֆ���z�p�ڋ���HS�o|d|��t&̥�,��pL��]8�X5���V�Y?`��$)}�r�6;�;��C�_�\w�Oj��.��4�Ъey�=Y�?�1$���Շ�w
PΑ�UX8]�+vGjxJ쭓釫o�F�X�%Z���t��}'r��k�����T�Oe��A������p�ݟ1S�[f��pOm�����]0s�9\�dC!/���nf3���G;�{w�s��i<�u�<���<〯J)l\���>�6���1W	�;U����@�L���_����Y|g���Ӄ#l���*�#i]JDf����M8�x)5D ��P�����t��r��OO�IV��q�H����p�n��@UǽQ��d��!_U��!}��۪ۡ�S����z�TH��@�f��٭����$�@�F�TV�{��g���ͭ�3�D���v����ʭYdp�/��d�����K)��nf$�MJ
⛝�?5��ʅ���4G�)OW '�����'�|���3�5� �O�"�'� �
E:Q���=��6�3
S�t�|ʼ#E�	��i����" ����S�u����b�wԦ�17����-�ޙ��ůޚ0v�muT�����g�s��]���N�eR+���X#n�h�M��ö9�z�n�Ӂ�:7Y�QI��J�-M�O;y9HR�����E7�d��EI�*�J�����;��L7Z�a���Kϧ�wˉ`��� M<��l��$ل �g�8#&`\7Y� vyfKtL���y��eq}���ὺ5'YLd:K��a>M���eP�ѭ��߳Ԧ1���(��l�?�y��>�2߬�֋'�RG�ܶy�p��-�rT���{ͻ���m�7Y�'�,�;��tFG�t���J���EI�8�^�HP���N:W�D_�/ٿ<��
�y������s:i^���&>�J�s��ˢ��͜װ0oV��Y ��H���M)2�0��xu�HMĸ��9g
�l'���{���>"��K��c�i����aa���kԷ�1�e*�)���b�5 ��T�Dщ!���/#feC�ۛi��;�g͔
�\%I�r�M��r�����z?=�Z�F��al�X��El�Z1�G�0ar���^�~��
��%{�6&����恰�ȭ�ȡ|��M3O�B9����5��_���4�0v�����;P�-y�7��o���u!����	�u��'�?A!�S8�7�6�I�\8�v����ڄ��O�ԓ;&YD}�* ]fU��f��������X�;�N$����F��X^�N������ȷ�"���U�1��1���q܏��~ �[u��uU���ҡ.f���=�_����]�P��û��W%�u�y�-V��i�M�X�z�X�,e��֗��N��݆Zj|�W��_���H�w&�S�{��$���2~�wxAVgY���j��s�
;��%�2& ����p*� ���m���5��e��r �׌\��E��\�����a�	�Eq�O��FJ�=�9�|�8����Az�f�]��r���m���L�Ӄ�8�>q$�)�{X�c�	��.~�QC�l[���jW�e�6)�?���ւ��6�8>���\���9|䳮�|�	�;+�|̊5A#�e��� +����j�p7�7b׃s">�5�RC�	��p�Og�5j���C���9I��̜��Ѭ�B��r���
`X�R/�f$1�5�#ƞ���ݸ��E�������O�� j�*�Z�B� �Sb�4�w荫��#E�r�u�@�J�%<+w��&N6L4v���6�	�
��e9ιA��,�����#VE�3��E�����';ߎ��%u���+is������l�&[��%�������*H�LY�(�:T�L���g�drO���u�����`M���J�[����1YP��b���}�%��4��(̛�+���vM{d�V�#w6i	T��;^B��l1���=Ӳ��t:z��C�u�1�sωk���$�I���b��75��$WK��ʦ��@*�D͏u��r	���	���b��\)] deG��������s^�f>G7��.l���
�g2fh��	&쁓��J��T��s�0����zf}͇�>��ݍ�(����c�j��[�u����c��U?��j�?O�vF�m�m�s�2��uzTr3�i~J���;6	_��.8���V�	��l�>�ؗ� �_�`do�j����)�)�Q+'lG+ ���bL�y�	�_�"��\zp#V�Id�"2�i�x�}7�b.ss�w�����	x,����y�AW���+���H�Ѻ�o����@� Q�H4�����=u�1|˙r��7M�'&�W/zr-���0�O!6P�vtr�e��N�Qy%DU��_��;3����^ܺꮑq�����K�����#p�{���S��a>U�J�`笻�RK8�c����'�;ϐ0䬳�3 �d�C�E5	A��as�ze�A@=�"�\��~��]��{���q?���� ��U�0ð��5��!�	��/7ޥ��Jܳ�� �R,�U���λ։����I�\{1����hHn�Ù�!G��9�����o<���A�J�"�+�k�h��N�9Ѿ�Y���a7��['���A�PC/9���ƿrmc~ʟ�C�r�(���u\Ǹ�(;��y㼜�O�n�qB��ۘa��A	��:D٣z�]i;чeE�?��<�6�`�v�-��p{ܠ��q*6n�-o�T$��us���n��HQ\E�Y�H7�n�a��B�_�j|c�˳���L��!���
����@^��R��:���%f���G��;. Xe2o�4�qe:l�hcNJ��}�[ ��+j���\[2���hfs_�O�a�1�s��"QߺU~��E*(�[}��Q>rW��s�����H��ug�΄f����РLъ�:.&{O+����!e���t�]'��]ґ�������6�)էL?c��߄%�>�qBzO�p&��h4vn�/�q�n0��*�ehڣ�k�D6������ם�iO)��̤��;��}���X�S�N��d)F3�YS�^a�$��[(F��l�1oI+M�����3���/���LU�7f�G���I{'����U5�8%��3�Cn�ԢUa:�HE�cL��$�#<��}��Aw�3�q(��O��p;g@5뺂�w�}�������db
��	������ɘ�bz�h��>m����1g[�4b�vxŀp�� �t�V�z��	�8�'?!�.�V�#&ZdƙCʾ"q���װ��*> ��j ���"�+U:(ޖA1� 6f�1��b6Z\x���m�3�0���h� E^O��՗�1JSuIq]�Ӿ����f�8�D��7C) ��!M3K�ʎ4�A~U����;��Fv6qE��@�3��K��'$���9���Y���?~�j�αݗ�ç4���x(��O��鼁`Ɗ�N"ZN�]e?-�cqLD�s��7^?��r��ʡ�9jc�