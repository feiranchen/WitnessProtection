��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O���u�E`��C�g�"�~��~�<�@{�<��Nּ��~�K5��o�=�^*����q_�u�~�#��*��Yd��77�U9t) ):i��6�"���B"�3��`��4E�pI �jpRxDB�-}/9I�Fn���K�TW?�7J�����~��Mg�QʭO�E�x l���T���-�/K8֑2E?�����*�ݞ�1�4-!��U��=/���,C|ͼ׆���.��K�N�=��F�;m�\����T�[���?��=i�}Y_3�%]k��'�HA���g�$�4�j�}����Q׳��}E'b��g�}�;�CW�6
�����f�H���4�_!= �	����)`����A��Z*S^�������R��eXx�z�L�$�q��ɫ}�ڷa�;�θψ�t��՗Z���=/P�v]D�����+(xۀ���^ �e��1E�&ȓx�DE����U�/��]I�V2i���f��A<�>�}t�XJ�$`7���ٜ��9AЌ���'�n�k�M��D�� �P�9����6�%{Y��|鯲��Rt������l(E�G1�l�{A��J���͆q�k���\wɋ�G�<�b.�8������j�C�-TF>����H`���M�g�OR@- k�k���r_�<���sPy>[/����F�Me���\��������G"�v�F#�ę4���RUz�MGz���`�����t��
"�O��	�{D�|@h�dة<b��҆zF�_�6������7�������l����`͸#�^/ȡ�u�	|'<#S(�C��/�*S�K�&�9�yO���R����d
�����n��lv��L�l��A\�؀H�>� '�i_�5�T�@Fʩ�¹̄6��S�c	�\�Β�!�)v�.������+����y���iR��3���m�Ek�-@�傸��to�he�[���-� �,@��F�b"��j��e�F����̠��lv7�PZ� ��S�\Mӧ�aV��}��.Q�c�nV�����)�U�F����:̆w�i{��^�?	�=ӝ�<9A�M�F5O�[����~&���r�%��"*�T'�
��Iye��&fشĽ�z8��L�Z]�,�
��SڗG��j=o+e�W�\��gɜ���ąBZ�M��O�`d��+NE�~�YB�w�E3R��2,���lϩY8�6z��/�.�s'������Q>��/г��Թ�<d�:�H�Nm��C�	���(J����c ��$wPic-9u�g�tOg�q��	
���<�uBc��`_�r'O��Ή��p�3ܜ?�PV?��]c�Q����lka~�N�dZl�H��rw��T�(��wb /�~�$m���]e);fw�4Z�������V�:�<�����C�ꗶ�X��,�,���`;� ����8\r��̊�����Q�P٩�mU���E����Iu��+t2�^F�.r$HҦ�!�Uv�`v�����gj�-�B�`�I(���dږ0CNE똧%�$/[�i8��?���h։o������`�A3@��Udo����a�Y��_
C��P�];� 8s����1�7wFvS��2F�}@�����{�:v%�)���K�Jt�a�E���hzݸ�d�P)ӧ��R^��Wp��@���:�"��{R����buZ��D탍�ߨ_
ۦ��{WS��V��=��g���q�ֺ[8�e�2�}QR��#�m>Յ*�ױ�X�R]��y}qa�Ÿ�� ەWL6�0��.��]�����n:|
�o��~��:)�k ~��T��.�������(�g�J?�H}��u�*�)I��|��B�P��$ڜIr8�8�b/ǚ�·ʷE]�y�����>�Fc�y38��`M�Xe� pW��b�VZ#x�H�~p$s�p�k4�?;a�=�\�3�ZVX�����
�F�Q��	�H�N9̷�s�����'_�-D����]4��T�c�g��3|;�'��KŘ�e�I�vE���9��=-�7�+w��Q�W]�M���y��W3�gt�#,Q�VՋ�gܱs��#]�1Al�Sn��Ĝ5�	�B��p�
9��-�_J���3������i�ކLe�_��"���*��N�*�6E��?-�j�Pl͓��lǫ��#��ŊbV�j��F�"#����l�v���/�,3k��#>�֗&�����3 ��{��"��Ez���QÚnG\����[&�����q4�X\i�Љ<�6W$�6&���%�JB8!�܍�c�7�Q}�X�Y�����ꪑ�YOQQ���Cw��J���;	*��k@���^)�-���,��TǢY�P��[��a)�OHZ��!Ih`�$��f �[�ᑊ�e��_�ǙwjzLk�H-=?]�t�Sl摥	Z�	A-wLf�������:5�uI���]io\]��#��;m�U�n���9�l�-^��M�4������2��#�>����*�;8�NJp�]M7��~�3D��{�m<A3o9#�����*�L�������ۿ�O�5�,�6�;Z��8U���َ�� �NO�~���'��єr�g����d��5T��*�Ьr���\���6�-T�D�!���9� ֚ jtT�le��64�u�:��H��P,����΁K�&��>d(�a��@����M���w�.�QSo�:;��x���V�6�K��k	��:�Ɍ�]D��]�-%���V:����3W�f/����l�����ķ�Q���-�4�@-�oh��	���?f�	�a�"ܽq$�Kәz���C��'��k�ՎF��s��v;���tq�ز�k���U�d�M�F�@�Ds�e}8�����1�Ig�[��h Pέ魵YWX�-q���xQ�_�(l�󨮩Q\"�Mϙ!��v��)&��vvG(�}�Y*������M�t��X[X/�A����g�ArW/�=j�k�S�6�����J�����'�I	Նw�>z���
�X�o����~c�G������Z�������	�������c����AVLXO2�1���)i����Ri'kV
�z���"��j ��>���X6|@��c~wM`���*�ԡ���"��P��Wwƀ�C�T�9S}o�������k�=s.��T������C����B�k�v�XF�g&m((&_�f ˤ5,���P�@d�$b����+\S�����ʳ���#�s��>���z������[�n��`-��c�G�-�'�8��h����=��
�X�PU�ϊ|��Q����Qg�g� 7�콤Ս��FwD�YìD{����[��%�R��7���%��R�;���xS"2�l��}��3��d�!c��n+��!��+����l����4�`Tٜ�5z�����-���G�GT��0��ݙf�y�P����0^��P��W��'����>����2#E-F��H-;P��� ��2W�4�ݺ$u�`�ƚŶY�2[�<"o�l���f�z<g��Y!,��x�d���/�*L�
8(ՕTA�7"{�����h��괖�{в���a�QR�Fv:i�3G�N9/�3*�]����T�	N��ߙ��K�Ϗ�!_J0@�J�
��Mx���c��������5�9$�*�=�Bޚv�(��GWm�qkB�(&,�����;����Hq�;�pU�˯�Z�l{t�zo��x�8�+�ߒ�s�T�? }�Zl����/M٠(�}�=|�j�{�I�~o�ޮwb����#��RϤ?��&�N$F�%#����gW�Ɔ!\��:����_L]5=���~Z�&}��X!��ZXB4�<K؍�������ػ�~0k.Z�A���CŇ�=Y��:g���%|-@���8D�b����"���^��9W2�MY���QnA��J1A�&�%8Hy�m���2�e������  NbP��2z�~^��K��N����92� ��e���7�VP:;u<��s;������y��"P�oSYW���פM����ǆYV8����f���~5%��W��E�3�717-a��i)B5I���y�t+�Z�JP�8q�!E��;�
���Д5��`s�vT��`���D.�`�[i��ǃ"P&EY�\1V1a)���jV�{��*�"�LO;���������
�lڄ��~� W������K0�"|I�&L�rC7H��y��t�H#!���Y앨#����+?��F�g,\[��e)�&;S(�!Z��{��]kOd��i���ۙ��r-�2ݑ�[���������y� bb������&��x� Ry���(��t��X�ғd�$�tZh�� wY[	�
jO�ϟ��z�dZ�p���,o�@��0tI?F��e�����Z}!�i���eH�pij�'[�I��,p����IMr���2I��� ���Fa�nzsv� �d����������A��U>WX�,�����Ca'�!DMd��.�+A�����շ�ą���b�e�8���q��Qws���5��h�	�"��ۊ�>b�M���~ޞM�B\����<j����%��)Y��3q��� ��]/�����*�4#��zF�/"��=ɡ���J!��Y���2u'-cC�Z�>�����j��u� s����r����j��/=m�q�%��@�P���
�V����F�ݶz<�ny�Xi���=3�g��G,�g�dPw��j�o�>����(�|�%3����JF�b��s8]ͣsǾ�8)����pvM�l����R"
�$�
{���|$d-������@Gj�MF��P��s!�BOko�)/i��\���Є����%
�f�}����8���$ɩ��Ȓ�.�(#���'6��oe��|x�O5��U{�t��N�<C��օ�4N&��i�h�(r������I�]���W6[d^�q��B�I~��v�S�>�a$B4��_��~|O� ���h���L������/��p��	�Ay�ֺ�dh�|
������D��L�Yݥ��*�+ܡ�(�Ŭ�|YV`�"�J��h���WNؙH0l$,D�L\�ڻ�@=n$�]��ח��h͹�����掱�eP�|���O>��qM}>�� w$l֩a_۷�JXpl1Q7�&�<�^����n���-�&��� &[~�c��z@�z&'�ls
϶���8k�yF���^�� @��4m�+�V@�ǰ�e�� ���X�d���g��T���$��.�+��ݝ!�n��PĦє���)�@i����ow�𫔄�*R�e�~PF�����PM�p��I�>�SC8ϝOz�>p-�df%�����Ul����l�\R&��LF�e��!�SQ*�mm-�^��֏1�ޙ�L#Ì$e��h�W��^ ֈ;F5�40P與~��mŽ�u�ӈtKe����n^_�p6���!�;FlHHBO-�uA�-~�"b��gO���za��NV��I[��k䴹5���w�A�2�tV�+^"���H�q/P9y����n��L���i�1,�Lj-����^���^���Bb�iz4g���4404�(V	z@��y�bI]��W��ӄ�vr�p��˄���F >~T!����Pzv���B��ﶻ����&�Z���"���D�y�������v�١����]�U}ᆒ����w��0_,�V
v�𚖌��,��C����~��tj�q3�J���ҵ���k�i4G������vͤ��=�e���}n�><�b��_i&[��㸅6��6�-�Ԉ������7�[�i�S�X,P��m�Z6�@v�@�1�˚��I�O�o�B�8���ma�{,H���/�C��!���2�a<BC�s�Z�b��7H�jڄ�r��߭���5�TV���(��QZEo�'��K������Ca��+j��c���Wix|`2���o�e��FQ[Y���|P%�^�-E`\���>��?J�G��Ti^	�=Gc���`8�Ef���{㒌�t�(�>���Ӈ0�C�?Mh�c��d����2��x��p|� ����p����������o�4d/��	2eG�i�,:�
�V16+�}?�i)��/tS�bڊB0�ǁ��+�;�̐A�"�g�9<U3<��Aؚ1h�!f2��E��@�4Q����1�ˣJ�5r�Qŕ��������K:�r�$5��/N��N)o�Gl�U�ru#�f�,b�w�����v/'@��d���\���_=I<��{�3c��t�ٍf�uF�6*r5��2���d(��e���o�:��\Eg1k�Jpfc�[��z5:0b�pF'�t�w���m�?��އ�ڋ��XʬWQe��m��iu�K����~!3j�\fd�y�6	�8���9����B�3�x�"!W�����vr��+C��%ɓ��`r��F�Q���>�إC;V���GKJs~�9�Jg��n,9W�W������V����"�hNC�~�Q����T#ʊ��ݎQ ��PQkԿ�Nr��|�o|�U�ҠݱB/��j���P>z�0oCzI�uz�r����� �����|\�v��ѕ@��-^�NC8��w�HB4rZ�3!cLy��#�����8	PZ����[���q�h0X)��ȵt�:�ޔ��G~Wb�m�� �}�|U��9qP����"j7�S�P|P��Q~e|G�t������M=�L�3GHb!T�ʻvd��8���G��(�TSѶ�*HG���S-� Y��Ɩ!���4mW�	���>����tak1�U=0׾zsۼ/�Z`ET<�SFF!X�o���T�x>*1�*k��G�NjD,O�.-}i٤�r��xKKr�Fۄ
�#v'v?�e֜�5�$G_�V�M��¨)Ѭo[̝��V��A�p@���р�Zl6w�%]�'���k�޾�o���v�ECޫ�#ؘ�#S6&��ˮ��T�M�l�A=�I?́�1-���nVl�|X�uJ�0Ҡ�ی�Aw��h
�����G��S�����"��4-+�KJX��f�w�W3K��'9���p �}�y���
r���TY�-�'��E�ve;h��U�M�i�7��AQ�Yyna�;G��y�E3�"v�*;m�G%���YfP���I1�~�ERQ������x}J��e�g�]b�7�G��9����9;mo	��gS�FŞ5�|M�U�<�[g̍v�����Sx�*j���x�����