��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ��N��������*�%�rXwl`��|�1�Ev}�-#t�1 F���?���%����Q����V̇)p����yzoD|~<����$|Q������֜�SU� ���0��Ѫ����n���O��𹄯4�<�b-���)��c~`I�I�)re-K��)�bo	I�X�J[�'�1�b
i��$��ŌD-Ca�����y"�X�p����A-O���,�:�=���$�����^�ߛh��ܺv�K@��!aް���И9~������7({̔p!"�h*��|yk����L)8�(�=��Ģ�<��%�iI7+#S%0cP�<7Ͼ����ӱ�$T>�7g��n�!���~����;�QW�����x4�짡�)�s�*�\�x����#�5��0x\C[�2�R�
AN1�ԍ���Y��x�Uo�����y5�rY�%^x���>:t��Ӓ����G���,i���<���1�^�Vx�>�?�"5��-�N�蕎F�x�s�;K�D���� ����,������f�ąĈ!*��#�{�e����=:��c��d��S� ��V9ٮU��j�r��}�)+�-"oP�/u ��I�MA�ޢ|��p���%�� )c��?Jq�O�
4C��ϮA�_�v�|��	�-�cY��CG �	���#���:�Ĕ8&�.Ľ�E(d@a��W�]��&cݴ��ƻ��b?K�:l!U�7	(+Zzף&Щ������n��͙�=��5K
���}jsx_D�����֬qw9��9�K����
��f��<`��rX�~���|����JŤ�4l�Zq��"m��]��J�M�\+3]^�< Ew	����|�พ�~����c��^w�&�'��%L�c������ ��i�!!����e���⼾���Rc	&_��q6m����m;���RO(ؾ��l��>��X��b������t��猪�Jj������������DJ;�j�q�#,���A�Zu�/s����v��������N�Hq&���%��mF�w��Ca�H(=�&!}�UM:��8�K}���������Ҽq\�(+��f�A���7������]��,��nM�R+m�l�Cg�>�73�s��}\���Qt]�E��ƶ2���%������:l3��ȉ�d���h!$���2f�������	 ���G�:M�Ok��̼�Qt��h~Q)���`4���rC��CJV3>*J���}�&����E1������4����α��^CsE�+w֜���k����;�������@<���:U­���xR�:�B��5�ri�<�㪹_0J%E���Dػ�0�iݠ�e���\�]�7��4_v,k�-ǳס�//퐽�4�~��߷��1�7��S���cFF"f �����r* �������c��Y/�����H/��g�RےX�"�(E�Lv$LT>�o���^��c��vC7��?�?8.Ws�3��#���J_mSZ���]��ʏ.0�"�'�8��_X��|�M�Ahj9,�	|�8`^�K��Բ(�T���{��	��?.�j�ŵW,�;���w��c���]�l��Y��Z�恦��d�L�w~�$x��K�@!7���҉��1_��d]�K1U�8<سބI��*8�0*��IY�W��o�٦^�\��k�� p�3%՟�\��=x�#)�&�Jۗ�k�e�3��{.B��i��o���:h�p���S0"&�n�k���4���h�,b���ԝi'��s�r�&����������wl��%m�� x�򻥝�0�TQ"�%�@Ng�xr�WҜn�tDkح���Et;b^�k���h����Y�ȅ�]D��:&��2@�`��)<VI�Q-�\��9�9����J��"LV�/���x���Vk�#�z�T��i����&� �P���5n,�+�V%=!V�;X:�1��v�$&5��hКB��K�KP�iڊ�Y]�ȿ����*�����}d�ߐuc%9�Y�q�Ϸ5؀�;���6opY�S'`o�-��:)��V���:KeP	Y �S
^	����9�q��2�)�s��{̕l-���"%��[~�i,�n�=�9�EL�X2��G=<��"E�4=�[�*;�W.����ҍ�	�S��2�I���m�q.���T��� �Q$Zm�q/>��se�����.kY�*������阇����M5��yp@���C
g�QǀQ!Q�����"�t�k���T�m��t���ؖ�x�X9ω��cg�e���g��P����`����rg�?+%�"��>�i"�a��!�:�?���6��7�=T+ȑ4��Q�,p���^<X�$�C�l�T T�w�Vmt�C�#q�.u|�Z��Ъ)#&W�D�H�p�1KdԅW�(Ӈ����H���-��'y��E�����}\hp�����";�#Th�0T(�u�N�Ugs����{�\ug��!��)���%��Ɖ��5�'�z���^�
�ѥ58�BBm�<)���g�W�����,J�.��*Z_��or�F����	�*m���B�>nxԓ����1�s� z�y+�݅3Q3���-)W�7�t����u��-�&ֹMi*Ҹޞ�A2L��z�yᾝ-?��q@Y�'ު��1��s���X�@8|��x)Ec��A.܁�	*31f"l6���v�Zk�ۥ���������@1���fH�����i�>dI��F�H�x;�(m��,��5}�L�e��P|�Qc̈́0��C��1eD�v��<q�7G{i���֬F���3���v�8=ĮB���W�����Β��B"Ōq�V�k]��H3���cWp���d^�]���+�����<�e��*�c��B���HA�M�z���cC�
�Js���g#�#����.��`��3���I��a��߿����H;+6և���h0\���)��d��"���2WWI�xr�bW�cة�4^Z�j�e�H�*jf#vT2��w�˄��3s�aϼ)�R�D�E��/$��2Ț�d�s���g��o��Ycx_�m_T��!��;EwG箎еȣ�V��,�=݅���M��w�����Jw�r�Ow"zg8 �� �����_&m�L�[ŝ�p��4S��>|q!I،=(@��,e-�x�K"Ms���.�wa�	(h��ֺS��bspc��WH���op��
Y��D	n��lr��j>|�D��A���Nȟ���y�����b7#�q��d/�R�"NLƲ��դK����<������uj�s��j-��e��	=*Y��OK�:P���~#�R����w�{���d^L��}�z4����#�����H�/])O���D8C4�:\��%��c�&L�d�7���h� �c�|$����޶����e�R���HyTH;gY�^�� ���.�1�S��*��L��gѬAf�%���My�E������(�������xv���|���*�
bÖx][�����[���ـ��vIKW�H|	�|7,�OO����ſ�����i@��u\��'d��@3���k�1�O~��@�oPCH��)dЭ�.l�h��k�\<�q�S
7�T���E�AS���#7K|�
;�C����ɈE)湿�L*���A�h���V�"�	�p�|�nE����FvD�Ʊ EǬ��2���=�X����J�g������Yzj��1�*�8!ᩰ/���6�����[B�T	#�N0� r��Gps���(-�6���f���U�iv����d�+7֘���%��Ψ�1&t=��a�h�c�;6#ˑ2�^��P�ח٘1��j��y�6!t}o|�cS�B�uI�=݌�v�p4�����p�<�"��z�]�'�q��w��:��j�$w��Aઙ
|��h��V����'X�|�$��/�~綋8�n���(oC]��u@��xʸMI2�f�?�*�B��o��9\#%�q�3����f� ���0���݃�;n�;�=�I!��R_�(н�����ؿ���Ђ;��:>�<]���$����������"����uBUtI�>�\�e/�t$��D�5n�����hNL��֐������\ܐ��vKD���b���r�{`R��b\
N(O���3}�f��c��ƳFwk�M�h�uy��crB��������w�z�>�̱��T��޿�'o)ؾ�9�I�d��ص%Sym��a���$p�ͷ;D�ea�xlZ�/������b�;�q2-�.���@�HW^���-��d����`����u���������	{�S�3�.
���L���3�㫥Zd�%��)���"C�&$�#�������7?ē�
�������E�OD�%S<L�ũ��Wzɨ`�9�9����.+ы�0ԡ�x�qܳ6�[�~Ɖ�:U�;�κ`�Qu�ǜ��/gV=ijγ�pI�p�>�;@~yu�k3񈌊�Tp�X���l\,o0�x!� �f�w`9�M�]��R�t��n��ɕ�����Rc�Q/�ʽr�����c�u�N���:�h���G�o/N�Zt���0�x�D�X����#�JS�0������ʧ%��W�oҚ�p�tG��'��1����z&�OQ�u�AL��ɬ�5܎J�nW���B_���Q;-�� ������R�6n��V�!�"�:�H0t1�}{"M[�)2͕`ea�����`��7����x���7:��[�-����=�v�#�=u��]�3�#�8�'�E�£���#g9�E�w��_�AD�����i�D�j;��(�[6��QݬS-������TS~1��P��� ���������7G0�r���)��c!���?���Z��n4�čE���Ś��l=��xe����+4v��f�V�s5�����w-�T�xߪ�/�4���o-y� q��4Y�Y縷fR��u��4��Zuw���3%Z�jt�d���T�o̰_%z�nW�S"t�4!��_�.\�\��cŎ��;V�U��]� ���.����0��Q�MQ�,-��[
���z>�\��䚫-���X��v��ДQ:�#FՋ�w�.>""C%M�Nn`�H��82���=ǱK��_�9����W��W�T����h����:�)qm�K��8�hl`�hq�p��`(q��6{o�Ӿ��Nj����\>����ye@���l�7�O���p�r�I�n�B�^:��x2j�8������G��Ќ�iJ��A�S��y�q�9h;�ԡ�9J��)�H<�J��Z�G���j��tV��`���x�4~u�ѧ'�C8ɗ� 	U<�N71ڑw&�����XI��XW��|Of4�����Di��6���H��Κ�����c���7�8q�g����s�pES
ACn�L$��J&8��+�:J��;x��'�ր(�k�#]C��Lm���'[��]
��ط��b�fE�|�_�N�I]Iu���9��j?��w�d �4�����MS7���`%ѝ=�)�þ�6�_6��.� �AQb�6��G�%�m4.M�.	v�+E)�әZ����4h�����5�`��p�Q��5��an�J�B.Rkhh����usMPZ�7�i�DwTE3�WWkb�
K�����<}��T�<�g�ʈ�z�h�[��u��p��G&��S�5N4�sl��M���t�;����k8��>����/�`p�&�U����$��6�|��	�/�M���|y��
�/0���@��s�&���ʉ���9tS ���s���}(��D1�!�������n��M ('�S�*A@I3A���O��F=D�����"_p�REM�����5Cb1-PGU�Ʌ����F8�۟/�'~ �aU^U��IՊXD�+�]����Y�l�/bZ��׭�h/�d�Z�(>Y��%W
�R?�|C���o�pڸ	����M���VV?����	��ލ�*l�,��t�V�V;����f�>�c��P*��Y�K�Yq�:���Z�n���ֹ���ڻ<�eQ$��v�\��\`�\f�a���ȵ6d�F���V��g�5�f�����wfMxZگt�\�k�뮔�a���N�%���ؘ������wwq��  ֋ت��5Ml�V���[�QWj��S������B	x]P�W���k:�ik���z���W�^E"V�S0T?P�O(�Y��s��˅*=��Ӗ<�Kpq��v�j�-��_c�K�z�� �_���C^�]�q�D<��yzN�oH���f5)u|Rb6�d���ᕟ~�:�Z�AU�Jr�b+���h&|@E��+]~4���R�h���"��IfQq�J2V��ojN5��D��7�ߎ�?@��̅l���+Q.���4��#��z>�7�����Ĝ�o-+�@(T�Hw���~���gsƁ*��>g<��˘U��� l����󚹬�fj�X�;^т�G'�x��W������k ��V:
�:T�hOx/��bG�y���X��X��I%��u.�|�8�÷
� -wF���/!f��\���1��N�6�:��1+��zw�sJ�]���٠��3H�4B�U*W��A��X,$��+�K����!����	L��#v�7�`��
���Knn�dJ��L<��"�.�}�Z,uF��%:YÜ5������r�?���l�JA7[fuǍUC`���,�mC��2$�Z7��*7c�k��Œ�ZB�k���Kd�c�g���9���a)�2�摦R�Y��2Rdp�����0`2�y7��G�7p]<dt�4�=] ��5 �|Ķ���*ŷ����ޤ���4�[��~�^�|���F���!�e!�BPKB����=��zE��S
��<5�РS�����5����Av@I���*3��$�b����[�"gt��A@I�K�v$kI�J��!`y\��q~z.�j�V��7�L�H6�1����u1V������@������9hЌ�o �<�^��,Bqn������w�����R���w$�Y����Qi�u��0���cNM�M\��\� ��F*Ic�%��Y�I�>^A�G�o�mS��G�ę붯z�r%n[�1hrR�nu
�aWm(;��pZ�oC�Q��+�l9 �ma�*)w����O���I�3%ra'M������M�gYP�?E�����x�(��&g`���3E'~�/�A �%5�}N,7��G�7.��+ՠ�i6L�y�
������;�n�ȇ��_da_�by��UA[t^�>2��؇obQi>�=��� ���e�0���%��=@G�,�� ������/
�B����}�щ ��rW�����5Y�!c��,b�0�H�R��-�8��L��2՛��~�;����X݈���\��� �����q�d �~ �o�E�R޿q�f�9S����7	�_ߎ�e}f��*כ��q�yEx�Q����_ܪiD��z�}��l�i[�q����}������&m�w�)����T�{�~E*������6��� `PSn��0�j�4�#ʱ;�y����C��`f��1�!"8��e$���72��0�[�`~�>OxR���4��k��37�FfBvo��,�^=S^�КyI���NrMb�����ڲ�^
�(���ͷG�φB�l�T�r��W2)uq�Ύқ�T��a4� ��B�9F�H���,��|��I�0��A��>a��Nꂠc%W�m�:z����(ͨFĦэ��W�UMEqd%�ʹ��������d�1@s���(���Q�=�&Ē��Q��������d�2	�����w Ȳc+�.A^p$LAE�������xa*�O�S�Jx]��1 o/�`?�@�+�+ <& ��ds��sl���5��"vx�����j�y�B� �$8,[=F�&�.�Q���,@���kOM#	��n0�eXM������$��%[�o��Q?����
�f�D�](\vC�����Y�����6��W:� ���L��9��|{`V�R�!��$�**���݂��d+�k�b��$RG��(�v����)\:L��B�}�C��1F�	�Bk�b_����v2�ߨgz,^�69�7�x�$�M��1����f��?�OV"w|,O�FW�^�/�+
<�_�7:����Ƿ;7m��D��:�'���N�HfZ���0�H1���3��'�&��C|l�6!�FM	��� �W�o/i0��?��慯g���A��[�T	�`��6�S���Om��,=����S	�4$���
B\�*���b�ǜ�!�J����d�;�Z��@ {��EgH;v��i����5����"���3�	SDw3���D�.��qw-��)	pE�'�+�D�vzwb}lzK�db@ ��7�+lr#�v����_Q����
�(��x���BTT#L�i�\Ub�?3l�(�;Ca_�e��J����J�A�t��y���܄�ڰB���ayS7�b�ᅡ�<�&�+�I���a�o#x
H��w��Q�k3�ba�PvUE��d:C�ღ�@.��r3q�RC|!��#��O���M�,"�y���)~��8ξ���?珥�O
�6����-kC�u�D�r)T{*�.f;�w�u��9�U��oT�0���@6���-@ԯ�AE�]��� �Q#��a��3�&� {W��i���|G�4E�ѕ�s���~���ts�Q�A��R��&A�����Y�Bַtb�a5��R���T§
�}h@�ˌ"_��zS�W+L����w<�K��%��� !�-1��Q��!��4�$YX�yj:l�_��Av��i~fE����']�(�Nʌd��}�Zd�[���	%��9��/ʶ�����B�L��'�����4nu��.����T�rl�'*�.V ����?�@E�T��晞�x��JrZW���iM��N��/�nr*`�=�Q5�"|�r.`�js�=���m8Z�}T!k�����\���3�}�hJsr����}�"��D6��O�tn�q
ma6��j����Lީ
(C�&�z������ @R�3B�Xg X؊��y�Y�Wϝ�<	��B�[��m�Q�cu���9�)��	ΊH.ᡏ������H#���e�oE��g��%D���wƼ�
_;f�z�����F����s�W�i�)i%}�� ���]eT	�#�f��Bkٛ�I�_Gӧ\]��{�l��-�jo�u�({������Q�8�}\Et]d�J���1�<G�?���W�-��ؿ�@r2�z�~?x�T��%�c%��d�!�_G(��������-�x3C�o�;vX��@r%������C|���pD�B�&| �5��t�ʜ(rV^t]M��� Y&C&}h,c��gO��;�H�D�ب��Zʃߦw��o-�U��_�4��/��Q1{g��r���%�R����#�e���<T�=�b��4R���¿�$���p�L�I�o���tEQ+���J%G��Ƅ�E��s`d*�zD�z��
���W2ҕ�}�p�Ǩ]46�
�}�
��*;xl�H�？��%�v��OP%��䬿�&��+1�U/���(0�"�a�+�%K_m�j�wPe��9Hh����3���YTR�9R�0�ݓ5]F⧆/���Hb_�Ga���ݼ�w%�'�w��Př��XZ�/�`}z	�Q��IR@֛GfGY!d]zL���u�>�/>�{�ӊL�_&�(<r:z'���˜�G����i�%&����d��Y!�C�/�*ɘq�xH:��g�b<�-��S-);΅��U���%b[?Ӎ�/o�/���7|�9
���z�2�~����~)�=���ݺ�� ��	�ǟ����ɓ=@�y�K�ui�'%r��9H���_V}^�7��9qr�����H�	�3Z�Js��׈��s��!�|)�᛾�vߎ�����)���p��u>�衑E�U��X�/s�fT�8���<]=if�`��W�֞���]����8����Pz�g�Xc�q����i�m��!{�睝��p�����y8-1'�w����7�P7�C��ӿfì�����[�/���D(����l�D�������J-�^D U�|���0�jP<l�S� 8TU<*"�A�y2��l����3\���\+�z�xu��,���

�����˿�W&�h������ol�/��b !'L������U�Hˀ���A�
���	������Y�w�+N����B���U�sG鸧��t��mD���1�{�������q�Hy�8�(vF���Fl챝,�r�&�d�}U筝\)���J�^��̪vG��t�F�<��؀�j�|����d��̮��aa��8�%��"	�O�&l�'��i��h���>�O��W>{XBF�HI�1p�!��6a�d!��,7��M�� 8�E�e���D���y�bʼ�u9Ѳ��L�`������;\P�aUj ��Du���R<�x�I#�$�[F��̯A����9(�Og�P��qR��v�p��R��}���:ҾN��Tr�9B����!R����=�:��=ˍ��,ί�_��˗ǰ����&�W���HB^~|*�^w�V�:�+��Y\��6�ND������{*[���[ �A�"p%� ��S$П����V�����Hq�mYS�M�oi����?�G�6�q��0�w�J���3$=��T�a7~ɗ�b��J���t�;�Ⓚ:"�i�h��m�6f��3ͅ$�e�a�O�R���c��B��O���`�m�x^�L��sw�bSG�<���m?{V�0s��#o�2�'��v:r�=i�`l��7�!�<�U�`e��7�̥���΍�xySL�;-k��!7��ь�(�b�QX�,'�u��Ί?Hl��8�fh����.�Gv�%��8n����q@����Pt���c`	�M��~uvKaT��d����#J�/��N�`-{P����f�����8q��;�#vl��й4:�
�ɞ�Q.y��֟��?���7ķ�c�7��d��B��`��T�>�5q�f��
���XufV�^?<C#���I_�%��t并�NoM"����0��v���Ap���L�OO�������ksj�*�_%�	����&�xFؚ�G�^� ���ict���S���z�l��+�
e�����z�f*%$I��ŕ��ye��k> ��.�'jP��b�aEi�{mJ��NʿQ'��k�	2��ԡ�Rd�5�ļ���+H�k��Ig�Js��t�V;�;���p �~⳪�/=�49P&ʃ�ŀ�8�k�N�"�2}�j�lr�.�5��Z���qi�#��O� 3�>��������-ǿ����MJ��A[�ev�x�=���Ѥ|�1����M������qt�/qD]�9��PBr�mj���������hK�a�v^��/:݋c��8�PDA0��!��1���54��e������G���'�"`޹=s�(�`]2q�����	�l�1��3)^}=I�#�P<��8٤n/�mZ3]�����D�r`�8$�$rU)q�y۩�=~O�?u�
x�������_?C�����d��774@k���k�:j�(�]hcVO��)o�x
��KBє�p�O~�����q,ŀ8c
,�V�X��ϽLH�Z���t��Yt%�}� ��7|ճM���TO���b�?���mR�C��.o[����N�"���'���$��5���0ԣ]�զ&�!1��UPs�ԧ2����$Ʒ\�W�����.�#(?K��-GA�"h��e#�y`��F�CC�h�/��{���`��A��A9�a�z���j:w����a�\� �=?v�~�Fue!�7�Rŉ��M%�ϐ��}Ѯr#~��3�O�N��N�B��r�D�FX��=�t0��2O��:q�U쎒2�YC�d�mb>_��Q�Bs���^����
,��5#�6��Q�˞��(�c�d���VG�v�@m�f� ��0u����?� �4ș"K��|���F�6-׳�~�c���s�ʬ�*g���ѩx�(���oz>S���l���������vϲ
d_���"��)!�����l��/�uf��\�E���}s��̯)2���1���Uw���>�Ƞ��z�^�*����P �t���)3@�
[	mA��B"�h�2��0��""�M�Z���kW�$�.87�B
ǎ���~^̼p�B���'[�迬�4��������Ws,���C�x�p�cԍ`UCD*�֦W�\h��
�1���Y�0+g�w��E�-C��yE���J�7��א^�Ч�Ũ=�i�	~ղ� |��~�ٻ�{�w��]j�-�J�ri�;��(�h]צ����r�4դ�{��*�����E�oEr]T�d!QN9��.
VЏ�sFecȡ���9��נ�,����o�i��ݯ��TWޝg�c�
`�8L�0�G6���8��֩+;Ĺ�������@ ��8�G
~7׶o�ͱ%��cgA�al.-�2���9��:�`R&M�U|�3P��	�'D6�Va���q/�`�J�:����5r� �!F˜;׽m0E��ͯ�81�܎�΀s>�����5À(���ȼ�˾H��V#��\+فy�G��i�]ŋ��j<�`�9�O
4	Q^䖿 1t	�����~�j�2�Uh�v2�����i8]dQ�	��%Q����BT)��hΘr�"��#ۑDE�-,z؍��2}�;���1
�v�Q
�=�a�Xǒ��a�`w���Re3��|��CF������^R�w�
P�be_њ�I��
f�3Cc%Q��_0
�4!z0)�38^{62SA@�3�T�����3.p�g~��"@D���몙��M��C�eu��l��z��Y�"� �)��bs��	��U�Xơ:l�|\�E.@Q���#�pfY�m)���ŉ����Yď�A�'Z�q0-�dY�E�d�ON<ik��F��Zo�Pb:Fjܘ��g��L	��թs��)r��&�fh⢕Q�K���;I|�����EU���;���xJ�GJGj-��瞙�?�yΡ�eL9�4�k0���S� 7�?���f���_�!�Xt%��� %Xd� mt8W@UQ�rS���lchY25��`�`Z�� #	Ey�(���2�q�$�Ez`3�(r?ʗo�C8D�c�w_0U�9g��b�ʑ�#�m��I>Nh�|�#vX�v�h���nb��C7��Р�}�Hy=uH��da�ny�5>��G��7E�B��i����g/`T�"X�� ��q�s�]�Κ�%��p� ������D}��2n�;fVrõ�g�?�:�hk ���*��,��3��m.�U�R�5�TK̘)(�
şx����%��@���?�#��h!�N��	��r�l�l���,?Ԏ�s�B�멧/�G��?�;/��Z�!��_��Vr�~�Lѡ���t�տ���I�u5Y2�aؼFc	F9�c���W�}����;�}A�XeS��K�=UK<m~��*�A�=�ޚ8���	�iK���WZv�"��un"�W� DeO���-�øX�E�1y�� Z.&i�pܐl�W\K4E�CDy��w�_{e��ą��k���ʉ
0�3'c�ŭ��-��N�\���m+IM�8;��o����I��7�Git���q�0_��+��z18��ԏ��">��F���=�wnÞ3���[�hC��4N�]ͧ��d��j��Dy,����z5 ��җc�����,���X�v�Ř����4�D�1 @�横9	�0�Qp�]B5;��]�x�X��8�N�Y�x���U���Q�����j��?Ԃ���(� ��H��Û�$�j~Q�B����?�U���5�iأN&qT3|f�;����|�<[��tm[&XE�7��U��غ���q��w��c��nx4�;�5��J���T	�L+M�|�e����&@�5H�6�%��,�>Ɋt.�d��o�)78�����(ǈ uo-^��9�z���)xxmIVFrR\}C����}tU9�dy�����n�2c�Ϛ�6�Jģ`��&MU��s���i����Z�ѢR~
?m��VX�r$TmE��HwWY1���o)�	O�*Ӿ�l��"�?�����RbHF������w��F٩{s�����p�� C�*�}L؟��H��EL���ݚ(T�a��΋��ml�,����R��g�>���h�`x���Yw������\�H&�����S������XW�ZT�DT���0"�z�=�~j(QH���J�&�8��\$���>�P۲���>�oҰ'.��)�Lo��6ޛ�>?2q�K:!@k�P�$�{\�|z���&XZ�G�Nݛ��d��%X�y����и�(&Ȁ��)��N_�"q]tv?Fi!�"�t�!�r�Ԣs4ͫ8Gف��Q)�A��*Q�����X�_Bh[ #�b�7z��cw�y��l��h07Y�.��LMp-K�Y��d(�"�\�������RFs�Ψ�e�Κ����)('[�� z��h
:��� ��������|��/�9�;g/l�aU�̱�.�CE��2��ss�o!�g�$-�F��H���25R�ж',es�����m��(�3ea�#�9��Ulxᚶ�"e��7�+/TUޣ��[z����6����E�ȋFݿq;0x��-[l|�C��ސ���o����܎Db�g�h�]Bq��Ј�l)B�����yi夾`U~�Q[������P	0�{�%o�r���0��COu"�0�{8��L��mf�+���f�/���PC�=a`�%/�J���rK��b�G��QmOsd%�Ν�M�K8~�����^���L���(�!Si�[Kw,�b�BI��i⪈$z��|	F��3"�6.�b���)�%�y�jR��+�Im��AvP��m�.��p���{xA�9��q��6
3�+��:;\��n�d-T�Y{X;�2��q���^i��ݨ} Ŀ/��ӔT����D\f��{R
�kUҌdڏs����I�C��P�T+
�a#�� s�_�ɥ�Pƚ#`��s/����a	�ly"v��l�ݺ��WU0��O�!T���dm���&��j5t�S���>��D�H_C�7xI���vq4ԚvM�v�بh
)M�A�yà�B���%���D�O�F��k�
>e���4.{y�h���k���k`�;#��"f����Y�݌��5�b���|h>s ����[Q�"��mT%�.��cJ���l>H�BHL�f�<��T�wd�\�>����.��VY �CIV~�7/��9i���uj���h��XM��Թ��("�cN�W�f�e���_*^��r����0��n%��éU5��z����7�� ?5���4���6�� �A L'�����Ѷ�M0ʑ�	b��O��dp�c�dt�>�nM6B�_�rrr����~�@Ŷ��_�o���J��^��nW�YA^B��h���]DQ���� ��ÞK`/����^zh� X���}��\\ǀ~8O�5�V��RKg%(��C�ћ:�^�5��6��31X�����?�1����.�j)�q)�f�H�����)_m������E��Ŗ�MtЈ+�C�'��������DM��﹬�+�;�GB������x_�5^̢�<�����<7�H[�L�߁������ErIz�
�V�끭���̬O��x{P�X�'�vH�,8D���b���$����N�ZK�a�����=K�8t��\|4�݈$LT�H�}�IM�wIrO��L�9�ⳅ��0t�s�����b8E�L�P�n/
�	���	��`)���J��a��H��Γ5%�WMA��cϦ��wv!�.��h|R�:7�4V\{a�}��Ii��v^�7^�|G��@�	�7u4�`�,��4�^�^ �[�u�^o�L�b?c��M�ag�z7��/<i���`��v�B��}��^-��/%ti��V�y=�t79`�v7zj��N������	S~��[\����!_�H�0X��H��Ej6*k�<2����cz���3�9�d�6�4}Ǳ��Y�Z��U�0�����M(��%G��R�c�AN�8��4����u���>��z��;.�R�#��`�ZN�;���Y���X4��5�����Z� ����ʳ.'�%
��q7w���A1E(��\��z��¯�#�.����k�! ,���@R�C�V �%�z��a������p.������:�����Yt�;}�CH�5���g����@�Ș�7��$��r��/��ŷ&�[`S����\~�e�ʆr�шU����<���=�W"o�4z����+��8O�vĚ��	�v8�%����p��J�0�P�����M3���u�8,E}�!�[KofٌD���1��p�#�Xo�Y�NH����*\�0$oh�SQ����(�]b�j�����ۉ$��4ĢŹ�^������/M?;��H�Ҹ���B	Y����L&D�Q�̶�)-�1���V5��~
�R�H��-B�p�5 L*ġ��D��|�)<O����l��hW�ɎUK�u��d2'N`'�T/����śSyNu�8�V���Q!�2��\�D��EaHۢ�[X�rmX�Ǩ&W�n�輁e�C%�b�^�����**D�����c~z�nK�c�1ԓ��3���,w�Ki���A���?,��������� �4�$$[�Gh+X��:���/�}]��Y8��LhO$d�
��,#$2��v �`�Fs��zO�B*(�aߚ�@��B>�,<�� ��=$vj,�!�չ��j���m8Ayl�JVi	�A���Ls����<W���&���c��v�Zd%\#�04��˷.�N��`���sv ދ�^)�	w�,I�!�i�]��զX��U�����o��Y>��$0M9�e?1Mq�aG�RW��퉕����?G9U����t3p�:.����g����c��ZZ�c��ݑ.�I8��*���X�*5]::��� 1��:�йo&�jv$�����lֆ�����z�Dp��&_�1(jY��h�-�V���(�<���=��>�񅙗k�h�e�{�>�(Mgn�STMJ{�����n1/Pey��ma��w�!ZnqY�����aI��*9�N�B���#՝K���*��=2�aO�$�3��燁�,xSYxx�~o��z��:������DLI�#�8h�B]0��r��\M��VĄ���*:ާ/?W�L�2�:��5=A��y�ӳ���vq�];G&��q���l9R���cQ�*�b���%�P��Q�H���%���o7N�j��3�:A���W�V�(B(��4CͅF���g�Ѕ.'��%��&�k޹��OZ �\^皂����S?&6����w7���Z�(��ʛ_�����B
̖+�v����	�q�X�4W��GJq���h�5m����|:�KB3�j����~F���=�\_�0�h2���u�̹��4�<&�%sr&HU��0Q'����M�,#�ʿܽޏ��؃�k�%V����8���؊0��i���`d��%�&w� �}uj�O��qK�lH��cgw��Ġeg��$�e��v�z��9� mV׺�Wo������WjMr�"�N����߼����-��/'�; ��0~�J?=����@=�W�B�9�/4�7k���a~Z��U�@���������86��m�
���٭Z*����@��Y�`'Q.1��5҇�����������~��g��R<.����c��<�4�ؘ�!���s����+��W�� �(�$`�����W&�-��Fs��V�֛��A�h��BY$���_B*8�,k��[ă��e��%�V��!r{ȳ�<Ìm�\յ$b�q3}�b�0K4�6a�pn4}�:0 _�1`�Y��5 �~�me�|��6��K��Hi���._?OJ��|[Шv��x&��a��үp�U��o�Bcl�tU��mgAy��� �]��	MP��?�TH�B�~�Z't��ug�Jq�����#Z� ��Ll6:�fB �
�#�Rv�O`x��[����m5AL�2Or`$H�X�G�i�Q2��Nb>hEseB�'��p��f��<c��΄EV��׿�<���:��G'�Y�1%G�c�w�F�]��f��-�Ӵ
�e�������-�&�(�e�f�!�
'���4b��"�>ELUq�ou�������\J�)g|T���:�fY~��ӭ� !mCh��ξ��i�WIj������[w�ߞaC��?Ԇڥ���9d�)Z(�6�ۻ�\=I�t���h(�f
�D�e�o��gw��M�iKľ�\O�
X
�:���I�L;���qVtf?�t ̩���'r�K�f�d�"�4��+aH�#�Wئ\O� 㮘�'�%d�#_��M�	<8�R>��)�\ŌZ��Y+�O�Jq���o�o�G5Զ����h��ҵz��P2X�{��n�E�:�m�1q	ڡ��ʈ���d�v�3�0BT�a�a���@���h�3U��5�r3!���s��
L��x<G��O߀���+�n�����oi������c*�qE��4* oni_2K����"�k���c��^`?�Tr:"�q [��R����hĭ�UPN�ґ ���kv6��"-�1@���H+�Z��m�ۖ۹�ʤ��v������蔗g�����V\�0���K|�,�	�C������F>�P%��3P)�^J���e�D�����w�����	5~���PLXF�z��E�Ƨl��^����'0B��"����|�H��KE�rS�ME����C�G������O�·Uʖ&�R�N���g��)`ޔM8ۡP�Z�H�$�ky�mU�;t̟!��x����*@�L���T��ʧY�.�+��|�,�@��U��aѪN��x Yʜ6cUP�g�� y~��|�P-M+KB���:��&>�[�v�.^��G� h�@���B6�a��9|��<�.��9����UbVS���&D=���Dl�����?^�?�j�l#�4,�-0�Hȃ�vT�;������n�zNd�5�_�J���<����{z�H� �l[���,q64R�2~P)`�e�숖�
���Y'��źb����љ>��x��[���8����O��V���Ev@��w|�ؖ�6E9<'.{���ʈG2�`=�qۦ]�g����/��ǰYj���x�/�#����F��	���a�A|��J�!FZs1�!�`�E�v��t8�(��S%Z}t�7���SR~�}?��u�`����1�
��](B-\������x����"K$���ɨ�-�J�ï�>��s��<+�Ё��H�&N�5*���w��|=���\=�f�it���¡΢2���΢�/�5�=y{�A�j�r!5��i?�)\�)}h*����Ćq(#�.�WOsW��D��&%$g,ؗ�~!S^6B$4�������̃�U���V�k��RY;�e�Y )|����_��������7���nX;c�3�� ��
~����N1<R�6u{��U��˱I��æ�z[�Y���?��
���?�ہImt�@�����H�ca���\fw�+\C���2o�g�1U��AC�xS�ɚ>�[[��D�ɸ�I��(�o�"����N`����d�]<���[Z����9�ob�~<����A�N���<����<��teZ�T�G�R�]�\'�'xK��?||f��M>C'x����e��(�,L�ʏ=N���\���`������"z7V�ψ�;�lS�K�}wt�&��z y�~mЇ�Y>�HO��#���^�裨�0���A�a�o��7�פ�����e�pw�*f�1.�"4��/���O��u
oIYj�Q�F߶�Is�A�K#Ϛ�#��sr���8�̷7JYq/^��Q�B_M�h��������.���X�ݻ���@�3��`c�8�{���ret�O�pE&���C�H�)lb'��}g�?�kG��c�p.�Xĕ��Q�V�pv٦�u�$M<�4��ӖU��D�	X���S�8�������m��=z[���ܱ;�H6�տ�${�j�q;�A���g�\�dK9U�<�v��Lf�d�����c�d�w���^�;.�+���t3�M������e�wiwXY��,v�KV�~�<>` &���9n-m"�����4���m������ῆU@̠�8������:z�X%�8'�t����� Y~3�4^v&�i �YI�ʔD+��%��z��ٵr�gc�NrTC�E^Db��0�߳��y�&@��8����w��o���c]w�I>"��}v<b����d�#f_����g���I�]��]1�M���HL����8�c��H�(����!�ƭ�X*�1*��QG;P�[�A�Fy�:0w"��86A�~��❊f��������T�}�ވy�9z�3��c3�*D��7A�C�b�9�n�n� T
|�.���l��j��|�����n�f4:�y�.(���W�LЗ��<E!ؕɝ;#��ÞR�R��yj���T�T�Q�hu�6�Qاc�sO��� 2����h�n(������o)��E�b��r�A�gev�����գ+\�����7A����t�Hmv�1���XF�9��^�dl�/�����v�s��=R��/'�$�Ǝ\P�v��5�>���O��҇��x��]/�_������U'h����r,�!ӊP_����"����!�Ŕ���	:����5�wmqT�5:J�o`:k�{-���x���ͼ��=%Ue���$H���D�����m���L�OY�x+p��<f�nNl׉���CV0�Gn\�����/|���a�d�w���fá��R��&h���hF�"��]~|c��N�.[�&�r��*���/�����Y�!셏���]��hH0��!�,"�i%��cy��Ł�G|��C�J���%�5���kFo"�%�V�θ��&S��ʃ�Z���2m>�=X�n �>�ɺ���[���V$bߟrq�v����ݷ��$�ѣi:�������� _f�qU1�����Ao!��� �9m�(��z�K�S�:��G�fn�*k�)C�܋�v�i�}�#�-usy�·���']�����?�ŭ�)
��A:��:��tZ��C(�IxI���ҒH(G��C�U��ʡ������;��ڿ����t���!~�{2���&�""���j��z/kb�����`#�\�w��eq�L��<�I[�çc�D�A0�U����y1���Z��D�UY�/�.����샑�Pô��TJ� ���\��~���`�wGc�菉[WM.������<��];���5�:�$Mq�X�����4п�eŊu��� (h�����)�/���S=y�Z�S�m,>���S*o��(���]\�y�Pڔ�!�unʼ����g�$龭(`d$7����r����g���y���'.�N4�0��/����ڻ� E�g�� \Ĺv�W>9L�,ᝊ#�p䓳�g��l1SUZ5�ʃ�}�.�9ey6���
�i�vp�j��L?�|E�a��� ��a7��(\N���?�YJ���iU�A��5pڡ%N�����G���z��#� ,������G�c3CK:y�h���K�9ʭ��/��ّ�E���
]�]_�ۀEƦE�6��h��$]Z�9>�@�[��p	���i..�dr�X��/��5Κ�i�4��?��3#�pC�zer}�Կ�V�ʋ��������1��=?�W�@�\ſK2�r�"�ҟ�:ס���^P�u��_|�RO�'°��z"�b=W+_����
��X�~fVq�_Zrp��iZ:w�I鄑��Ύ����l�o���[�_y.]ٌ����1�+f�e3iAޑ��Jua��K#�����d�� >I�˒ 5�=js���
�Ї��� �f���M1̏�������!�b�z�ڦF��h�w�NpB�;��%.v
��v�7�im���0ĨKT���V�'��pH�/���	�e�R�۱�?eqi��s�O�'��x���7�=+��������J��{5qD����P�P�n{���y���̷��H���q�ġ|���%�R���f���\v0�[���}��ccL�l��~,'���@��&��������1O"�R���Y$�)����m���	(�(���{(��Ut��XzS2����
Ct�׹n-�	�:��~:Z�|�#�&t8v�?�<pm�;j�8��}��8U���?�Q��3w��4���BQ�]B�Z>��ѥ|Ŭq$ k��_4���B����:��=ܤ���m������{��T[x˓;��޷m����\2�� 
���/U���t6*�6�o�,�ܙ�LW���Ac��^�#��.��������6��Eu�:�hI�'�/�Ήx0r�}���!���ٮ��������ԗ��aS����C(�=��^E��3�N����@�(�Դeړ��q�	�&t��PIj���*g���+���)1ylbV���ަ�*�.���W�1wQR�2e�n��(��-����(g�����O�o֑?�l/jr��X����v��6����>=,ad͇T����4���\�r��`|�Ny`|�7=$��G.X ��nƶ�t��P�,���JB�^Ђ���{,�K�s�F
"5��+>+e��k)7O�[L�� 'M�":\����3��4x�/}Wg1t���m������Դ���,�v�@A ��hkgQaݐ�`�8Uՠ5A&����G��W��'��Q�Sn:b��|�wk��)k���]�W��;*�^ôi�2��)d��-^�%t��?pT�Bo�S�=
�fp�Ա��"�E�I�ջ�!k)�#vj���vG"u�y+�OH��*4>���'Į��y������ܵ�ZRw�?8)|�}���Z�m)��[v����Y�����!���N��~}A8Dfq��l�đ`���\ZDI8����H������T���rz��3�`ƃ`�N��>�h����s���]��Mk��wI>q��.���u��X�긥ԛ`�;W�Ꞽ���U,��C3/7����g�l]�Ƽ� �˷�T�?�V�r,%C���Y�����ƞ�c�Z;����� �[^����c+/��c�J�;�JƎ�fՓ�4�h��~��ܕ�� JZ:}GdWt��*�@{��B����ة����B����o��fd��j�? #�v��Fe��ަ�un����2Ȧ���0�PV�ȯ�@�"p8b^Fd�2W���~#�����:lp�a�L�r%��&��h�X�E��4�2���F}�o��74���ͽ�ķ�.�O�w�^�w��yy�����C(��Y�u���"��Bˈ�3H��[�\�wh�sw|>J�e9��2���l���u���6?+&�4J�*t�*�%A��"T|����sS�'�h������YK���	�~a�"�3WT?V2���P�g|�dG샐@(�u
>�}~^�A*���
Ls.���2'���4���\�arh�����{M��v�Y=Ӫ��u �N��/����p�����[;�sb �΢��uВ�\���/�����h������ڐ.]�����TS(���آ؀x��*9S�f��p������b�-x�����;,.�JFIF��l�a�m��u�2���U�o
'^D!_w+�X��u$)T�!�Y�2�SG�.�od�^(~҂�|���&H��Y�_B�n�Eu{XLaO/���&#5��`���M�u⎫�P��'�-���9�3��{HFecl���8� ����᳂�`���ȳ!����� �7 -<ѽ�ΘS����c����f����R
([���a��	��_Z�|H����{+Haw(�������d$P\PE���KIo_w�[�䤏�l_"Z��rE?x8B)�`4
uo��{�J~GS�Ҩ�\ك����EA��7�~��t@�^H3�Z��E��b}����}|~�6���6IC_[�%9d��X�d���J�@젤0:��ln+ɠ_RZ«��R�j2[L�Z�a����p�)˽Z@9�Ayo����'��!�]�����˗wC����Q��F�;�OH������s��T��)1���灐ۛ�P��ځ������}Ur7�{+%^��g,9���|��{S̥��*E�!�>p���%6g�A�M��\~���D0Y��_0�%��H�bo���R�}����}�6#����?ף���^��o������v血��1��S]�ԗ����Pb�\xcB-����_$&���_�>�a��:wz^A!��r;�ԦVx�J͘[�i\�WH0H<6�N�q,搪u��]{d5A�ԟ!q��A�ȕ)LZR2}ɷ;��;�f�����B���X�,�V�����w�Xm7=��<��	�Q�?j�!!h7�G�*(-*#�&A�l�7�3P�F� i8a"_=�299�r� ����H��e�G��_W��')�V��#�	\h����=��1��%"�A7j��t�<�Wξ.!��D��5���@�L. ���_�&[��sAH''D�0DC<Բ]�V�pJ���Vљ!D)�*f�G��	@��<��~���8�o��N0}`�A�X[�m�>��.��T��2�:�4�>��y��t��M'����z4�XX�F�]��-��D��&E�br�9�dMkH�tD�A���ι��x�mu���|�,h������Q�\Ç���DDHJ$���<���پHsu�i��ʇ8���?�� �K�4 g��YG�.����-&*r1ҔW��Q#�Zë�@���O0CY�PhEw�W�R½ׅM��u�����9�ENy�[���������dK�2��a��"��~�!/QL=�u ���Z���鄦����%��B�e�c��X�OX�3v�	�y���?͗S��N�w��
.���F���-��(���u�_n3Hǰn�1M��8���?��+Y�b\Q�B���7�@t���{�0�$�p�Q�(�%�b�ͻ'���S�m�[A�H��_h�Bv$�4��&_^0e�i<:�`�e9�\p�����ͫ�<Rmrz���]��ږ��7�L�)p&k�T�}IMfj;"��{�"�U��H�~w�U��V�߹���z҄�Z����{ދ�ՍH�����@���ᣧ�?B�����~'�*�"��P!9R'���I�_ȪҎX�`4v͗qC.��\�����ø��`�QFor$����|*`D*q����[A�
�R�N�A�:ޕc�o�
���1yt��E3�9깾+��#GPWhy�A�^Q�us�B�
fu[PÉ�щ��nr�>���>${L�\��=0 ���j�5 ٖnzҘ5<ryL|��N!B��7v{{M i��)mP��4uO[����n��,�V-2	pyq�y�I��ቆ��b��?�ӊH+�MD�ޱIǏ 8�P�)N��MG5eR�,2���FU����"o'�5��&:�������;*�!�{��m��8l���J)g~JJsH�j����[��
��Y��Sx�AD?�SW�w렚>8
o(єP�i�=1�B`�~܅)�A�H I�wE�Ӣ�Cܛ��\��L����^ܫF���mŃJ3u���_�X� ����:ϻ�o���M���6��I!�(�P"pti�4�{;S"]�h,��/��-�W�����8���U�0YQg����Yv.G퍆-�W hU��l�^���ldEF!S�)V�V��Y��g?l���]��d�O�)-������2��#/A�����a�-��mR.�f!���h-v��51�㘒M�2C�0��k{��zd&e������@�ev�ׄ�&9��w<��;U4��>N~'�▥q�s��{�H�#�� F�£Ǯ6�,�ϔ�V�W�_�@.OZ+I�svF�U����ƅ#��4e*&]3m"��6��b�"A�<jTre�=[7�%b>�$�v���643�n���_�;���쐏��"G��IOЇb���;t���1�J���%<��:���0f�C[��)�ήS̼�s]��"��=͗��ׇ�̴�E*����qr?>�gb_������֙�K�G�H;pdr�[g�;,b7��?�pL��妁�� �B��X��K
�ZՕ\�T$��t���Ǘ��-����X�4��gZ�;E�M_xu�΢�L"hL#��?"j�0�c'�Ϧ����>5j�B�C�v.��.�F��^�q<	�nx˦�Ќ���JzC��Y��D�4Ō�
� ��ZYS�xL0T�z���&�ѧh�D�~�%�ݜo��W�a��;�+��-���)��{J�ʈ��n  � ����{;��`	Z�(�s̘j;BT��� �?@XZ�}��߾��]��2�x���<�<v��	��:��ׅi�����!h���Hs�!b�y�K6�z�K�%	g��m��.���XB�2�.��[Q^Dk�lbb{����]8�n��-�u�(�E߆�ZK����T��W�s���׭��XVx�(@ͩ��.�~�FdGo'���=h�f#ߵ{����ۼ�����<6�zxD������D<G<A��Ne�'K�-�!-�J,�3�t&14��?Y��B��~�?z���i�L*����t%����i	�B��י�R�%�/��3xt��Q���0�mn�Դo�r��,�.3��R	��.�����P���������HsB,���Dw��Lqp�g��:CvO,�ڃ��D���6a��h� �!p>�+��#Up�N�4>2��!g(�҈o��Rܱ�*3�k3ƭ[vɨ^@�LgZŶ���8��h�-�*'e�-#�����N�G�gV� |d�̝�(�\�����.�TB�k.>Z��7�<v*�x��[Ɵ�=���)����7:���D
 g��<D��5�7"¹�q���h-p5�H��6/5+���^�o�"v��xS<~T�!���ϗЄ,�\�ػ'e'U�i'�h�J���d+r��+�0�wT�ڝJ/��cpH�1n]�?�Cy�2$��E�>Ǫ_ ����}��vF�f�"]������}�)x�椂x�BT�:�7 ��� ��>]�j�!�w�76!�oQ]�W+k}%]�zS602�(�[��{�*��#�Z� ��l�RGݛ	�'�/}R#�J#+3��hP�vҺ�CY�e8��:K$���tHp%um�H���^���x�6cJ_O*e�	#<p�	3,58�Ґ��Ԡl�,i����(=�a�(`�
������ӔY�Uӧ^���lƵB���(��&|���>$Sn�oW�D^Y�&yjgȝ
@3aѿp>�؃���K��٘]��l��G[Զ͉[�D�*�������Y�\O��8�AHb '����b�_7�/��~A�|�n��:^���`ꦢ(����=�1KG?Y��r�n���1�X�lNџxR��[	��-���l�Q,uF	d}���Q�O!�_��g�l?F{���.ՂT���z��1#X��Ф�ݎ�`�']١�G��P(�z���0��"ǣp6�}���2�uV��t�&�Q�Wv��z��W>&#V�3``���
?�]V�o��Pmn�u������H( =�'*T�����x[������.�)�$w5�ރp�NV��h��`C���m�@��q��q�&� ���z������4�7�IѦ�s�.�\��%H���^�?���p;�7��}������:Ck�&߁�4���-��=�./Y*���ɯ-�j'� p?A<d��ޔ�0�Ӷ<mF�XSkP���H�u�{���+���A�� �j��?rԫۍh�)�>VJ �OH'�WUF���f��i{uS�e058�~F���Q��Șz#¨8uF�ϖ�4w���)�K�Δ9"��TU>�巭��c�.�W9~��yk�
�}��$>�"��zc�,���H�I����K���@j���R` ��''�^�@s�����/w}χ�M9����7�9!����1�θ�5���~
s�r�j(]�N6XINQn��=�<�Ź�cH��]�^�07���({����s��VZ�٧�.#���9Z�7p�拼�?�h����.?�W�������i)$MP�$��:�
��j�.Z;_�����d���[�o��ӆJ�O��E.BZ�j �+�6f��.���<<�Y@���)��O,�eI�Hہ�D}:��d��z�8�M�$�}���Ɲ2�M)nÇl�~��@��<F�Ѯ$p�}6Ҫ�:��W��'w}pZ�݆d��O ��Y�xE�\�4�>6��_��- ;��)��a�ao�x���A�|������9������auV���w�s�4'ߺ����l����3��Wy�/�;��&�@�ذIyp5�%Jg���#)�s��(��.O�@�'a<s�e�����n~Z�>g�~<���}t �������:�.$*J�8�F^?��.�ZO8 W�)���rLaZ�ͬ���M����̗�:D��d�I3����x^{�����Ӓ�Qu��kZ�-���9rm�ԟ=���5g0G��*�>)&�C���f8�R�CԐqLEy�U�̈����z�eOW�1�6L����Ѳ�r��d��M�q��$���_�%��y@�����q_���iX���2�TH�lu1];b��1A�r���J����T�:9��Y���Q���gi��ѓ� �:NsVL�y�ND�2A��.Z�Iz;���$n�ϳ�Z�{/�maMS�>Y�(<s`�ME�h���&7�����~DjI��C��G���Y_�+ei����K����Eڹ��`�q�T�0�o�; \��Mhb��S�������@�����`r���$!<R���o�Qs��h_��������K`,}�/��^]#_C�>r�֨i���&��&� {�vFP�v�|��9E��~KeK�Ccnu8��s�Մ���KjOZ�&�=�Ļ}x��XE�a�p�� ���h�!���� ZO|٥�W���_Ѿ�A����O�K�֖���߈��мKH��
�l�z�0C(���
`ˣ�ε�l���ie��׸ͻ,=�8Jl�����v~��5lĀ5������W1�WHa(r���έ$�J�����)E˱��?�z�X��J x��;��,��IZ��O����hy��c�:/6S�.�?)e�?q\�_|%��Mp�˼��w���O2A	���+��3 ���uƏ:�]B�&�3OE�3xn��&lQd9�~� �#�XY͝�p:���~}�֠���IUȤNB<v��vCkY�k���Y��w9c�+I� |�.
��J/����N��ss�)���y�9�#��7+��e)�q����V�\����&��e����o�%��B�W�{�P��q�W!�W(q�Q��822*m �\*�cԳm�Sz{��-\K��Fh��{�5ㆳ��`|�Xy��j��Wz;���Ej��ʲ	�gV{��/p�+�X��q�!oIf�oGx����s\�ms�{��jP�����t�����Kw��+t���*�����#��M�vS���Y����+��[m�W�+����}Qg�����"��Nm��gO���T<�넲3�$�s�P�=�V��ʜ^�bl��R��4���w�����J7a���E���V4�K,?��<
�ND.�r�����|��y������m�o��(�ݯ���R"�1{P��:?Oڝ��]E������|�)���������oJN�4��$��M����F���x��|}�s�t�&�U��~6��%�fb��^�y��0W�����hhG}�b��iO��L�����ZY�RA���0��
=�{�=p�hL�&@=�
E�7�cRx�\�`D�b8QSb�k=6i�Q����9i�מ�_��GkNͦ=��F���MĂl�,���9��C4U���o^����� �]��6�!x�{i
{T6�P9Q��;⾳Y�fBsa}#�8�N�:{�ˑ�'�!�®�0mƀ�B�C��ְA���r*C�����"<��Z5FZ�"�?��E��X8�����snJ��e,�y8O������An-z[��'¸��*��ll��ϓ�/��o��'��K�Z���Cp)\ۊ�����9Ջ:�(�FWn�z�]�_V�~/twY��8��b�H����nL�/���pF���:�V�ݬ���a9|ש��),�r���i�~vXx݆��L��zؠ�C����㙽�.,��B:>`�hCq�%G�w��D9��9��O@5l�E�~�%�#�-�� �"�b͊@���uTR��H/3���3�2�2�<��Z-�����>�3mf�&�*.�_e�����D���mW�1B��j�_`$�p^�Ŝ9���y�������WW�N���`_�e���k K�	����!3�3DT��8Hʧ�f�] ��$�m?��ʒ�����"���)(�q$��+�гN\���)$w=ו=D4X,�S�JR����d�pk������P|��X�c��/� �5v�>��l�,�P�Q���,81J���~~V��� ��v�G��nu*Zlh��RU@\c������X	z����ZE��!�sT'�^.�PK�ݟ��|u���x��h�$��ni2�tN���#�a��=�n�T�a��@b��zpu,9c5©1��g����~�z�Ś��Pnܹ�2��nr�����1u��`1��:*M����P�IG!K�|�:�9Ƣ/bc�軨������S?4� ����"�@|/���'��s����YY��B����p3\&�ܷwr���2l�J78 W[�?�؛��A���W/pϾ�pȨI#����]�p�5���&��;f�1)��pI�+�-�!BW����{�1 �긚zw(�]����
v��rs`ܢp$p�n�g��7�����4s/��ㅦ������I�I@����I|�7�QK*���Z��E�Ý�8*$z���7��.=��-L���@�������S���oK5�qE�	hs��|��E�Ɇ%�+�\�߂�+��MK���c�|�ma���FݜJ�&���Y�9Խ~	�����x�-W�͸�6���c���o�ns� �kXBȂ7�@�C7��0H���t�E����uiu?���X�N����������dU�����c���sـO��{�;C�	����1I�����I��f�4�(�� ud��=iw�PiqZBr"�}g�(��8֓,�w��ϐ�}�#��JF;��25�vV���_����0���1��l?�ٿ�H���.>���X	�
e)�����~����9�;]��P���0��W0uؠc.�� � :��7�Z��pΜ��}�;Am��pB]�XJ����s���"?�|Ǘ++���厫����G���m�����A��>�!}D��~�fY�� �%׈�wv��W<Ș�;O���0F���ϸ����a䏐�9@X����l18�h"�o�K*�[��?��rQ$oo�>=�z����p�Xdі�Vv�*K�l�( ��6UߤUMF�U85KuK&�r9u��7]��+	p���9s�HE�#p��2d��\?rGr��Gx���\g�B�M6�i?�np�&ͼ�t�����z���V$��*��/�iG�Q�Btn��P�y�a<�*�� o���7��YD,��6v��``C�n���r����kw&�}��2W� �8b/o���wjH��W�)�\[�v?�H+_m���Hs3e¡���u�&����/M^��{���A�K<Aߞ+i���:��0�k9����kBuY��o��ޕj\�{h��"�)B�8~8Χ�V��,�1��_�2� �t�:�?Q\�/�h� �%���M�x� ��ӓm�Irs��_��кF��Y�Y��+B"ʓ!�扖�>�ZGq!Y���P��V����Z`���Z��F���(���g�	��h�]�H�6�,NE1!s �K�i~4vH�Ei8xf��`՘��+�QC��79Bqؙׄ[���9���0²�^�NgA��GC��R*�a��El�K�����ت�l⶗�����4C�VH���G�;Ѷ� =ߵ�J��a�(��]Fw��Z`Q�>z˪�q� T�G�rYrvf@��}�hkG��9XIl�KUO�Ij\�O����ɢ�ipF��g]+��O�v;��2�[ɜG"�]&�����9��j�zӱ���lH~e����6�$�յk	n]�+{���)8	�`�qGb~Ё��_��aa�2u���
=|=v����ϊ�ġ��s#~}��?ߊ�s�q�ؽ�ع���N�Ub�~���H��[˔�ǉ����(c�àW�-�ω��଩l*��e4b;)�K��ȅl��ֳȁ���`6[v��O��.�[��n!1rߡ���n˭��g���Yy\���z`�Gsq`
�)Bo���V��P�D&Y��:�'^���^.���ϋ�;y�T9�O�n<L�\��;_�%� �7��(��v쑃�8p�����yDL˺��u��6�D(Noҍ^am�꩔̰y�Y���#�(�=Ab}�Y�&g��5gA6��eL�Y0o&��&`^[r�``͉ �;X����|m0�P}l��{�� ��˹���~k�;
~Z&_�V\��&<��n��{;l��S��8M�S 3�?L[�Ҍ�1���!-��E]<�O%�Ko��`)�J��c�ln@]C��cz���\��K�[f��a��X��4�ځ�Ɇ.?t\8g��'�B���{�xe����9���ʣ���h;a��(�;*�vjE��]�MF�7���_��}x�k[Ad1=>^ L��s�������QD�Z\d�hZl�Ԥ��2��G߾AK�����qh�s��3���'�I����-�L����jkj)�	�L�����������\2
۽��,�����;\ )��n��o[��eGJ8GC7BDe�E4��e���l)�G/�~����v�2���y��ٰ:��n�K4��gcmذ��Xb��Q�,���XD"�29>2������'�"��t`��5�I�f��c��P��
\��#�H$�le�q��/_�g&�	�z ,<Ђ�`�,�g��w�e�?z4�c�e]�C����Iz�%�>�g�)�����\�ì����YJ��BA�� ���*��X����}x4�rY�9S7�C�K�7-y�2��!��g��K��Ô�PFEQ����Ec��VG�,B-
�AgP�Y(���)\�yQ�_�� Y?)���/��;,�H�B�x����I�J�U"6�4(��PI�-:	���x�%�oջ�7^��V�����9+/�	�~ ~?��I,ն4G��e��V��">=��ҠJU���D7�k�w���o�c��z�cD
��U5�F&�(1O�&ں��܏�
#Z�`��V�ua9�)���n_����%�S�'�=L�p���z?�3�%����� A��T���=q
.�� �K���mr�^<j��(�'���lC��]b�y�� l�%jyS������V�`���*�2�ӓpX6�]ۛ4�e��cT6l_��u!qܼ�m2�@����(�ObJ��[�� ϟ���O(�6��p"���#����
cT�A�@g?h�!�F:���+g�������f[�����}��>l������9�2\dqI�`��"Z���c?;+��'��e?9T������걓y��uE�H�`}��z^!��~nޗؾ
5%6���-?�x9���m���cn�傀��˺C��֛N
�욼=�Um����w�d�Q����eu{� ê��\���@
l��+5��YlI��U(�n.G����qQ���&?+���yAD��ȳ:
��}�ǜ�f�fP�(�M~	���d���b� ���&���K�ihG=��݃4�o�;R�g��+�T��g�9y�$v';;���Qr�����Gd�6(���f֭Vkb�Ǎ�����m���n�8Vzf)
�N�]#J_%�̣Au�P��6C6�1����&�o2q}�?q���^��r�ك�Z��o3���2h�\
�"��j"O�Kz�Q�����7�O�g�w����ɋe��
c���>N3u���n^���^�"6"��e=�"{�sk�➢L�21]��
/��iD\P���8ܗnhj�b��6�\}
�`7|>�P�6aQ�F��"�Z��`V��\�ERJ�ףּ��̪�=-z_�Q �!��U%\m����"MO��'�.�Cd�q�ؼv���el�U^��cP�4��&�y��"����{� �� ���'�hL*c?�66���ۆnz4�%�*���\zgmuvQ�����:�����L�uke��$nF Rq��_�."��FU�#�+EL�+�=^K�Dj靌(��h%��J����nT�;�l�X���x���s��9��O��ҳ�¿��wjMy^�},j�^�F38v?�G��mU)��O���$��"�[����{{w9�>N��T��ۉ�&�
�*�����ҞV�O�^����R�Xc����Y���pP���]�\�6�t��LD^y�5C_�Q���5iyX���0WA���+S2�_����p���n����c��g0\f�7���	x�-j���>2�%懮o�����v��Y�>��űX���;x�j���<��}�7�"��h7 �I��n>�G����ٟ���G�-�^;�F���Z{3w
�~� �-�.�OՇlcGg֠nX�lkT�N:�IfB��������A"CV@j'�}`�U���;	:�������i��!O��v轸4v������t��Md�v?��F	7B�o#kR��%.��z,�K������yJ�'���#��g=ba]�Dnׯjo����gڻ�'G�\���j
ܷi�1P`̫A&�0n�|37Qު�m������u��?xޯ�bq?5��e���6��J`�e;
<,EeJI�,7�Q��Vl�$��1ܲ�4(�pH)��=��'�,6�\�T`
�:�s���=�AvM��g*#��R��\�ޗP�*��:&�?�����i�{���������� �_p�O�����Ϟ��Sz��D}��m��7,�up�+F�����uR�&1����ch"N�5�nJ�>��@Dċ�?_�Μ�\J�Ϩ'��G2�s#��Ǫ�%�!Y�/y��Q�5A�\טX<8��kLEŗݼ�w/�t!���Fg�	�5,��t�h��D�r`�+�����z6�X[��VH@Uǻ��3Z���,|�`m�RϠz�
�˅n"��u�V!tV�e���֜ �Ԏ��)�9{�Y� ӊ�!hb���_�Pw(�hu�\��u��n�=�w���d�fU���b��	�cR��w��d�����@�kY���<�����á�^l�jqD;S�4W��J���e�q�z�؇v8�'�m���ˇ������:?Q�E�鼥P�H<�NS&@�xǘ�c�� �����ٞ�a�����yB�2I҈(��VE�E	�������}�J�C�ԡg-RF�G��ubo&z�qލ�ե��vP�A|"�Q�;���@��c.��=��蝈����4l(��֐Kh�k��ɝ�>U>m�`�Sd�$�'L|���y�wV�ǦMD���K9��H���͹�?�B�2R�i����+c�4�qUNX����i���x#�ھu��'&��S�������D���O���,��{������.�e�RԷ:n?�wF�|_J�Ь�D�w24W�T�7��)�)|[�>_~N>9����'vy����u�]$��#��90�e�7�K�_�m��	Z?�/�g����)YCZ��]vk;��}��G�P_0o��_�-�WV�'l1-����o��ң��i������"2$��^V��[r��kF�?�I�}k�&��M��%��~�C
����j�apnG&�V�fQJ�^���e�������	=Xb�U�ƞc�%�Y�q'��b�R����%��ߤ�8�4�EuB������qth���.������+P��v�PY��^�@7B�o�Os� ϓ��gxwkE`�9Ȓ���6������-�n��G"��v/J3fJP�����\�!t�b��
"��\�"�3J(�MBpZ�4�O��H6����ѝ���L)�e�a���TF��=g���C^�ç{*�/��ԁ����T�O���\�H&�ݹ��w�KM��⤅ګ�R�E�K
L#�\�W�RH����1r&��
���Ζq��ݞQ+�Pr���|������kzD�����<�瘟/���[�����J흳*����w��lr΁��>t�o��<gyԍ�P�r*t'�&�/�B+�|MT_a��x��+�����jKZd�/�g�^���,���!jeqy4z��3�%J� �Uߟ�ӹ�w>��4G������J�k��J�E���Сؾ�Ť��hFXSxjm�v��ͺz[tj�g�}5����� :��(!@�d!�,O�(�}���
1w��c�0q;�!N=������?�V+��鐥rop���{�-�f��(�|]#�R�<�q��V|8�S��o�(K����C$�h������z/̽���^��T�p�����ϊ%�����ͼY^Mb���7wf��D��ſ��Р��&�Ċ��"w	�*T��ML����|�|��x��4�"1ٲs2I}���|En���[��|�ܕ���"�n������N(m��D�H�T����M��"��0Z�����O�Jŵ�����ޮ�'m��;�|@!?x��l۳ z�U+>��	OS7y�Os�x�#��>�aqd�I����w*�/����1,b��(� ��y�P�@���)�j� �:�z����[�u*����p���;�	�B�dd	�8k��]�+���,��LȊ�^w�@�Z��੅�\��*��UZ�&�]Q4N��6�(�"	kf�UN����do�0���oC���#�pT3]���s�����1�ԋ��T�ϴݲ���:!g�4�jGK3ꢣ��b��R���g�PU���̳����S����i��i��<���h�o4���:�.?��Z���_18i?A���g�,�E"�|cW�Fz,Z��YbL3c�Q#��xX��k���ʹ�<����+��rS�"=HR�z�f�0�=�:i͠!�׵���\L���,`Z��/�F��\ջ
���f����cmf5P�����m�(���Z�qw@
�QpS
ͰPh5">�:=�Z+�EQSf�d#�n����|wܩB�y�v'�9U��&��2n�����D�Q]��W3!�h�q��.�]	ZO�๶I��%D��핏��X��$�Y��?�� u�,��jF(�Cuݒ~��Ay��y�3}�e��%�V�q�}������S�9%�%�+��"󝋥6�iOԪ���S8ޝ�1і`�m�����R+�YXUOe�Ԗ���hoo=�п�9��SPQ��V���M��Z]�i/�:O��Ӧ�D��0�6(C�i�	��2h	����{4E�$Eڅ6�o��ݷ_�Q�g0}��'��I���M2�\��K,���I�%oK9ԇ�m������W��Qu�0�:��z,{����2#�j����K�}��x�q*���@�|#��M��J���J���%Bw�y�'�2;��ª��us!̺�7~I�����t�]���4��[�HX��@��@[����Iָa��p�y	,òyVB��~'����o�F'p��o���	��&�$�5&
G��X|R�|"O�mH�ELp�WrӴ���T�˜�@�>ޮ^�i�F��U��9�8�7���zwp���Ͳ��U��2v�����f�\C�@m�pd~.K���,8����/��R�i�$��z������oaI�HL
0�&����?�#�d<Ic����٥!m�U�����I^��ț຿�V���"�5��!\��1�N:��������z�ߵ�R�їLj���p/�0M}�b�wڰ鮖�� ��Є+��=���f��������� Rr���T�V��N*G6=��.�/�؟�CO�)���̽
�����d�� KN��h�ٵ6��l|=z~pd��S����z�	^�����L�e�Vt֮1=X��4�>�(���b�}�E�c����̇�}���D�_��5,7�Jm'���UBp�\|1_��;`�1C���<��mGN�\^�z&��拓�j,� ���%o�A��X�Q/��q�F���B�VCz�ם\)�^���@��h���dMW=��S,���v���u�;�suU�aB�?��f�(l0��j9g�"��)�a}��t�o�9��e��y[e���ǵAP0?`�>*K�}::K�ɵ/G�J�:v����L���e���8��a
�S���n�����3�Sp�9dS�ɸ���d��
�㥫�!���
6�}`�I�pj�y8�cޭy
K�\�L�8�iP3>4`e3���(�����P3��s��h�
\4X�{�9����!qL鑧x#��pd��1�k���K�0�n�\���Ԇ�H=�&�_�%_��� ��W�%�55$9�6j7ʄ*��N$�eD�e�H�_�ll_b�8�A��IU���6�*�\L������Js}���79CS7������kuDⳇ��,��=}R��mK��N����I5��!�����v )~ҹ�
��a���T�eU�"Q�[@F�E�>�b���_Z�֜�Qj[����P��V�6LTF;���(ջ����r��L,BHh��Rr$��Ԁ���dP�Yʎ�ճ�1�J�CL�����ю���
D������v�-�u�9:�s��LR��.�rb�Sb�qvv��88����>�6q�[���$�ؕ���	{p��KY�s|�:Dm\��\�T������9r���Wh�S�gr��/�#�� w7�gl��3�j�r%�@�47*�3_竳v�7�T�#��8�e�Lt�c�^,���	��jE��e0���nS��t��T����X�;��:�p]$�����@j�F0�Ek��k�Rσ.��WV1�[[8��8����hz�9�Vd�|`���������irQ7T"��;v�R�f9�d[�)�WP��`i��%�K�fZ���^z	j,�?ql֙��@���0C�����O8�<�ba��XT����=��|Y��`a0�)r���ǶJ���	sA�>�<�o�F'a�&
���hg����o(�-b�m�%�[���?Is˜�F�V#�=�[d]�PƇ�s�d똶���1t{'_A�fm��{q�/�����~��|�V�_���+���ϢgA!�՗�r�j��6�.�y�+�1Vw-U�A��/���Ztkc \֌r_��^�{Sx�~~�PnҚ���xlP
���q�J���\؈6TJe},~��3vŶ�s,L��5�DLI#��
h����}�����an��~�]�z3T�q|nक़��)�v�
a*
��	wu�\�2���Y�e�^���\%�T�*�'��2Y��.�e�9-Ch�������B�������և�k�:�O���o=L�[M��#��	;��;�C�;��{�}��@���l���x̰���(������ů!��VS�Y��8$Qy��N���ɯ,�2�!�[�Up/>:��������wQ�m�;�S{�;���:��%�:"*kqN��ޡ[	*TG��d�����̤�N�1�	���2Þ�.E�7�UH��;a�e�3#�����i�z��c0|I'����%a_�#R�Gyg�'	��A�4w'�"��\�ﻯ�9$���/���%|K��>t��x�tɞ@����(�$շ�r%w>�C�
���:�v�a��O��u������0pwK:��6
��+�2�?P��`E^^�ʕ/��	
��$~�D��nW���ߗ�&厀7ML������~h3/2���d\��L����m�Dl����a��id�È���b�8B�X̭J�F�s�@%��$ �N
��-o��h}��&���D���_dz�g����J��=ɮ�]�f�$!-�9cd����2��_"#X��T�-T�g"&nD�cmi�G<(K��A��UAU�KN�|N��V����N�Q�V��K��%G�����
��J���9N��7y)G��+�}V���]���*�ϑu3���G�����'g�ȃ�N��B�gEb,�N 4����TƩ�u�w�d��*�Ğ������x�OE����`� �P��c�ނT�x0Bgʾ�As�ؤ��\{bS`~���/�}	�?$j���*��g.�p?���(C��a��������xl\8�猪��1�=@EF|�E����A�S.���(��.��Q̃�q҈�����l�_�a�ܸM����b������W[\�E�./�����N`��Ɍ=h[,��Ӕ��e�{�G\�g�������.���4�e �`/;j��NBh/9��kzS�WI��˂�������3" ����C]s���������l��S7��.�K�r��h]�X^�p��$�	�3e�7��k����J�~Ε֞��e�?��g|�j6tO��d �R�j��Q�Qu}P�F�#t�`4�0�\��#x��L�$��LFK�K��[�8mw����gY���F>V�P���hK[���X���g	$���o�N����r���-�lr���Hu
JUV����l �e�8`#l`W%� w��_6h��:i�a����?��������]'�BU@����Y�O�[�]������ؐ��y�*8/�W���k>ܑ��4�)Qq��M$t���jq�@����n�Q�	7�f� vh�C_�|�n��E1�R7`�L?T��n�?� E��+�)�K!�mEX�
mĕ���!H7ޠ����߀M�Ǐp$)qf��Ĳ���}�G��qю��*��HB���mnĈ���DyB(���-z@j�X�yq��� S��:��B�7����!�'�b&d*|�l�=њ���yg.��et{Jp�J:��h��p<���+�i��ox�~�|Pבu&��X?��%��МL������e_s�9sj۞��-�y�N�ÙA>����Ŧ��[�����K�����JA>>1�t����9ݓEF�4T3�tg�@=�y�>�W*�vbQ�[�$v	���Ի��9�V`���47M��.��_��V4�â�l��j�N�b�Nߋ�9R��F`NG#�K��dU�'`5��'k��i�zw��^�K�"ݽf,�Z�⫛��.�n
�:�_�3�7s���vi�����ap9��ۼ�O)���}�z�Nu��黽�|�������҇q@�Dܻ�pj����Xlul�*E��}�^��;f�ؘō�?�<}y)�pl^��s��8{
<�+�Ƈ�>m��-��TTU��v��t�/Uh9���zr�N��XY$�!������XQ�X��8��Y��5v+�G�T�`q=�g]��r�r���.�T;."�-�_����9��9��+٘i�6�m#�JD���^_�r\��1��G�kz������j�'�3#�@!��[��Z�e[�O0�;eb,\�i@*s5Z����=^��9 �uf-&��_��@9@���Gfc+��*��:Z2�M�\��b+�oTOHiTeI%s���ݽ�MB�b�z�����}ۭڼ�[����?Ga�d��ꛥ}�~�
�� 8�RЦ)#U���w����{��N1�3 �����D��|?�M�qF>h�Fe�v�^��fZ���cWVg�<���#<��?M���-����� ������آ�Dou��eDH�P����v%S$���S,ø{��T�R��@��L83ܝ@�`����6A2&׵	D1��-I�<Wm%l+O�,���Sn�\�?N2�hhJ����̶�U��u���;N� 1������������-C��2�D
G���[�x����ba!h���s�}BQ�l���M:�1;��)#9ς��J�qce*��Q'�c�]LK8��#�G�4����"�L�.M�����F1����l�:2ٜ�Mx'��m�\�1�f�`U�<F?3p� �x�h����mC�M�vg�V�E�(n�	;ڨA�]м���VZqu���WS�!�_w�JXŰ��A�Ut4.�}�0G����ΉmėYX�1<z�:[��z5^�ޝ�m+�@R���	�����Ռ> 	I�|EOI:�5i�8�E
^b�ۧ��_{vΪSt[,��Ŧ65G(p��g��-���g ����R����9V�A����L�7��0��FP�,�u��{$Եa��h:��ӫ�7�?qv���-aa4V;�V�A�W�1f-�Z�7�WV�r˾���O�xb�.���G��r���K�/�4�RϜߪ�(&�t�ϐe%y'��@N
~��c�eʌ�&e��H�(��~�/&GG�y{�����R��%�"2�n&~�T���ͻ���9�i֯�����jZy�Ԛs�>�i�MҨ�o\2,�����OeL>=��A9dܘ�)���5)����c~�)@s����Aa��ܺ ���a ��t.W���jڶ2N���~@?�M7u+L6U\���;:$J5�IC���̘F�2��K�nf��9H�*�_Ks��u�������yU�&�^���!�s��\�b�a�T�__���f`p|�?1�S�e���o%��5#-AЪ���ʒq�� �e��$�K�P�x��6�1lOc�*8_$��r���.��nU�ufk����,@!w�E��=۹�P�[�ޱq��"��/����iF^�SW����:�l����$�2�a7E�4���i7�7�:�-�?�Orډq�:ڤ,@,�C��u�b�ܓIR�3&�zl�V1��1 �W5.�5��yWt3����%�zVE��{=vI�:ۣ��j/n�����_��>�&R� Qj�ߢ�_QǗ%����y�n
���T���w��`/�[�����v���3Ceϟ�� ��ܾ-�=���y��ڮ�NW��r�I�e��$��sW�'ׅt$�Kv�n:�\�\��4�=��x]d���i.��dfFK�I��]�7�1��ۮ�8�R?���^x>���&��m�n��!��qd��(�Ō�XL^����fO��-R�06���u�]���(�cŖ��P<����1�2�L�����T����壟�Y�l�G}����{C=Ȱ�D�/�+�Jә�g2�.;V[Т�1��S7��_D����XTQ��m� ��쫤��F�Tf�r(�`�C��x�]F��-ZMȖ��y��oJź��u�NC%����4N=��&Մ{�Ǣb��_8p�MX*v%���(
'P�
R{��O�`��!���h�?Bj�d�e}F�f�߅���͘�I��I��9Z(����T�J��P���Bn⼂�`�����f���˟�C�Z(���n+� �엱����2��ܪ�.L2l0ʙz$����}�͆�u�X�c��a�̣q� 3;�	sFBJ)~H�5/.��G�#/�R�|K�sB��x�fܥ'!��ж5�wn�{:YE�8qJ>�:is|DˠI��Fͣago�&��y7�OmNg8���e���T�ī�+��2i@�rq��x)UJ�)��BHN%Y&�[����
d��x����NT��][�&GL�S�C$S�����T���\����r��Q ɡ�ዅ
�c�U=_5��(�n_��j �B�ç���@�)*�)hL�b,Ux|�.Lb��m'����������F���L�J&�x��[ft��|ۼ����27ZJ0	�#�Y�ե���Z�/��;\�s�����Ba_+�AW-�s�U�%\:�ɇt��Ι3��v;�0kZ3�{C���+��~w�Vu�P�m�M��+$h�?֗�p��^���R:�°���� ���/� �-�zF6��5��~35 ֚F�?��~M�?�O[���ُp�����t�:�Q��qމ/,x\e��d �#�_y��.�8�D���M�Yϴ�*?�����H?����mDm"�`jF,癆F��ӯKE�N+;����מ�9x�E^�V���d��\�T��Ԓ���u���ü��&�/�;?�����BZ8�!��GRÎ��g����e�%ג#��e<VI��&3��H�^|�*�|0��P�Ağ�!x�@;��
�|���,�C�1�B���GEc:g�VK�2�/����(V���v��%&�8C�4g�$v�@�{;��6��2��+��}	U��:F�IIګ�y�R��8�����9C�]T�G�R·�����N� �m��%��K��E��7�9\
���5	��z��1���y�cb��gxHeٹP�s#�\b}�	K[�\�!�������ia�?��Xw?P㶓�({��+L�pS��
��$�H�o�vN�r��A	˨�G��P�MNSV�����i-�����&=��&�W�2��OW(��ў�l�6T���@��v.�蹿�]$�xR�~����вn��C)��<��}P�]ٻ��v�O�9��;]f��?e��U|� �O?����E��M���c��%��x�����"1��jr����bᚷ�.�as��Ee7"�|��\��3S����!4�#��}�y彰����TN�P�`<#��������+�a�U���%�~f�!��6�0���#G�gi/n�7���y�	��HF�9S9�o���	"�:�/��G`����(m�h���*�&��GUA�U]�pH��*Ғ�������AnwH�N�m��4�H!9��,%��>�)����#J����Զ_���ЬO��4�ŧ��x)k�lu~�=9����V(ߓ��ˇ�7��p��'��i>�\.���<Wc���X���ٝ���P��v�^0X�� ���7,S�W��`gp������涣��J1WB��Ã�,���{�kЕ=�4�~�������b�ɳl$�yOr��/rL6�7�bl��[��m���5|���%�{%��V8�ʊ�r�M�b]�#�(/�۶�B�3��x#,=��`'~(�i�>5�`�J�6�3���S-�e	^Y]B�*�'��({bo�7\�#�o�;!`(.��������8�~�ya���A^Պ�K4:��Vε����G,���3�H���9ZD��I 'nq!;��_��F�����*Np+�"��|��1G9(s�H��o��e�55.ԔSaÔf�_&-+��%�t��`	�ޠ4��[�'2����>7#�z�?��/� ��`��q>,���Ɠ����#;Ɍ�;7�lL���G~Z3�0�
�[��8����-1�<��y���Fc������c|������['g���}�d�F��� x\@9Ѫ��'FH�!����,�9�M�|�瞗�OwM�s4���W��qmOSx[�hk������9��ix�����J���0=!� ��魃�V��e"�.�\4��&���RR��ʸ�nsg����<��]����%&�61�q?�����O��wJ����?�2[�w7�����r�hj�lV��YmJ�)^NъQt��UQ��!�c���x`�]¨� �S{��2�^pۺ�ɝ�_��̚��Mtu���bA@�(3W^��'�}>��T¸X$�۩�I�C҈�b��gy睡�k���7|�Zr��0��Xj�_)v��{�G���@%�) �}
o�/����Q^|v�o���R��RNQ8��g+������+��=7Y睁=�����kEJ뫰�9E]�ms8�L�r>b_C]ӂh	B[��5����$T��+O��u7k�&�ŕ������cӀ�e��V���9RV�G�%$��	��̸5���1:SD�fz��R��*m@����X蟒H/%���ŋ� �tB�\L+&ì�v�|V������X{�u�<�?�7^}{@�ф�y:[y���9��2���s��K�����CVg�9[��d-x5�j�v���2Z���6bN�	#bR��{=O¶kw��D;�h���"b��>�Q4�ۦ�$3gG�p�C�N���j=i63��\�ڤ�?'smT��(�8»aM�'��_����+�Wd
�@�Q�� m�2����eh['P��x���Q3@l���V�w#�RY�(���ӝ�r��|Rv��hf��D�|���Qҧ~V exL}Pr�}�uy}Sh����u�N��g|�R��\�)�Ң��b�0vbi����7�O���;b*/-r���#��-������n!�%$Xj�����������3����j�=O��)XhE����/���_Q�X2!I�D�{�z�y�Z�Cˀ�.�g3R�l���Ǿ���\�z{*�aٍK���1�"l�^b�e�ؓ�h�������ݷ������D�z�O���ek;�mR#���n|n3q
��7^<�����w�&ү�:7w]ࡆ���b��>!���ť����(�0{?f䡴�^�\A��nJr ��D��W���<v�Wl�Q�x�W��8�۞���l��mٞA	%���=D�nE��1�V$�p��?�%[�(2������(
��0OYS°\^ϛ˓�����Z����@�ԯ٧b�zccKߖ�Q�jX�*��K�F�N�MX]��i(P�� ���t�0e�vz������X��������Ώ��U贤5vv�j&�o�<_65������ظȱB�1�AV���Ƃ`�H��vAqC��U��XФ?c��e��ԔZNa� -�z��EAV�?��p��B��  ��ە�W03P����<Z��E���R	�R����$Ebצ�\�#X�s�Ë`l7����^�B�q�*29�Vw,퉽�@�706�Z=nw�}�o-3�lV;s����Qτ�חzZ*�ѳ:e��JJxrY�/ni#���̽&�#F�	ۍ���l���������,�j>�R���<����eN��X)�6��T;��Q�F{iG��맙ߪ���
��8��ZByx�:=�HR[�#M9#�2	�'���Q�%��6k�'�6��c�K�q�J��=<��8�A�Q8��:!:�G��IT��>�13c>/L�v7�WB�i�P:�_�@~h�	G�}��5�8�AA���W	@]���#G���/��s�Y7���Ә��/˩�%ݹL��TBT�W��!�{{����������#꓄��a��M�p�_���Ԁ8��`A���^�w�����:�7a}�3ȭzڟ�1��r?N'˞j	�w������B�͕����uў��T�u�9��k~��3�,/O�t��g�]`Hu�qt+�v.�yB��3x�^p�-�d�����5T�$吖r�U���XM�mںS��I����P��]��%X�ln!ా��'��1@G�jWeت
*�Y�I�,W����{UX�Ym1��|;]����1c+�Pn+E�#ʣ�	��Ee��["��@���h��RN6�0�ߵ8ﮅ�(V�&�R��1dM�̵�*�@y��.bF�9#hO�$�8 �1!.;�)�3]��&�=Ww���)�h��������e����c�F��*~�aF[���uT�_BW��~)���/�q���D���.��'��P3�.�eD��m&�`@��B��gO^IK.��F^�vs��x�5@�5�հ~BxZ��

�-�
�v�I1�Ȓ��������>M��L4~Hy�b]Ⱦ7vi�2δ�c}���$��eV�W��.w�0�Lֲ�����"�����S��4O��K���� P��);@/����;�st�mu�("�pP�ϐ�@F�E&�A��t�x���stD�kz��S�z_�ʡK͉^��֋�+$��j�v\t޾�ݿ;1뎘��sw�n>�������y˜#1.Md�j�ۉŌ����=�7�G��%dK��ևLc:��BBCS�^+��`�*ii2~�e���Z<�Qdb�S�7Ik
ecD�[��i�Wcy`6k�`X�ɲ�T3lz���k��9z�U��i�A��y0�Z��(�H� ��o?}ڵ����*���s�˫��/O���=����BP"[�P�~22&e�Q�h��'��Ѿ�i)�e"2��WAAS �[��?(�Eh:��a�`ӌ�%������w
���k�9Oe�k�`�y��pOCaYk�p��g�ޜz��N>�fK@�3�x��e����l��;�0�A�g�J��f��Ӿ�!��n�UT��������6gG=����~v[ө	��4P�BVt�@{�Pz�`J�"��B�ig�c���xZ���3Q�1p�^�)v�E�;aUT���>t�T?��Ex�BG�<�d?�[��>�%���4��}����j��z
K]�='
ŶE.���7�^ζg�?�0��/�3�m/������C��K0���˚!GbE���y��,��U�x)��4�#E�	��S��V�MW�R�Q�S�˦F�����-�A��O�y��rO�J*�j�`}�ư�������샖ҳ��Gv��?Üx���Tk�,b#}
�,�+î\�T�(�Ԑu$1�N��:%�eN?�6�4��R(W��B\����θ�HY}Ѩޜ �ǒ-���g��N��� q%��mDf��>�Z�<�A��=1mq&�9�D7k����2_�f��DC-p��H	��X�Т���z��Qӭ� "���-��я�P�+�Q��Z�S���  ��~�(y��(>Xef�O�i�H2�5Ӧ�28&	!?s�#�+z�&�-_2��X:3n��ùmS�As岯i
[>�O���٢�l��!��~;Jʒ�ۜ�JAjs���.��4��~���Z֐p���U1�)Lu4d��|���h�"�Q
c�` ��2�S�^��%i�8)+�@���5{���x��%}�v�K��
�2ĢO�}߱ۮ��̨g~'���uO���PH	�TgkB�V�D��1VU9��e(���b)�u�U0Z|�=BT$������rErC�D;���Tlcbܗ�m>?X-�t�$R�m7DZ�w�=�3��O�������=U����_T�F�#?�q����#�^΋W�̅-��4	�dmU��[�YT��c��"��]���j����`�nV�;;�N
�`��m�_O<������3b�w�ǥ�Y�CjqY��+���_�T���׆Π�bK��l?��2��²����>�sYt�m�;p��j��o�ʧ_��;?k�<<����7k�-���Uʺ�K��h��S�H
l|?z9����B*k����Ndb ����}�q������=���wyf��d�(�Υ
�/*jN����}��0���J�N	;�1�o�/�ܑ���J2T��W�sR��n�f�_S� �[>F^z�#��z{�,i�휅��=���ۣ�:�-W�lA�>�;W��&�(�p�qn7�2~���N��6����X^��w�X0vJA0E���q��H��<��ۼ�m�{�(�we�}Z���NF���򜀡�5�qU�ҭSL�Ǐ?��aZn�E��璟Y��Z}�5O���a�R���P�W-,����.]�^�@��,IRo� ��{���m�t���P�'��@Id
��~�۽�w"fM�ז����?C��>�Cu��,W>��o,j�Zo(Lp������N�C�}��T��	�C��}��e4�o�2�e�n@
]nkS�
��*��l���\h�X���$Xp
W|މ��Q��%��[��_Ѣ��v �c�OབŻ2Ax�tb��	�ߞg?8��cf� v��g��Y�!��e,�x�TP�Y�5���gEz�B�l}�f��]�(�|�&bH�EF�7��}����ڕ���2#t( ؼ>?F@��|��ȕb��>M��"��b�m������?��)��p���� �Xn�{���f퉜71�֏��A,y������0w����U:��C�a���:��