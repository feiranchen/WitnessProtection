��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+y��mG�^Z�7Y
c��z�&��p��&���B���
���ס�9��j] �&�#&0Wh��p������[������Q��S�{"j�n�n��O�K���J1k�я��)��X G�4.�"Q^��kHS�i�$m�M%����@{(�i�|Sh��fv���n�`H$�S.�iL�M�6�@�ƏmpN}�C&.��/��g�_�(���JDALheMI2��vw?�n���/��ED��:�̴f(u��F�fҰ�U��,�<{ ��������8��Y_���?��+��`oH�To*	��>�20PIj�#z���6���nX"�TV��ȁH���>4@�{VT�O�4x7���E����ҥۤJ����ո^�D6���@}l]��1
�G�����5[H�L�6'0�_�2�ӕ�]������χu�f�F��[���n`WI$�A�FF�����ܶ�3`�+�SsFX# m�1փ�s���op����B�#S>b�t���E �j�$�;�����BW�xԟ|j#"R���bK�e��|��%�2�_��>Kh�V���<��i���t���Ī���1���Н��W�F+u;��@7(Nv)��T��*��%7�Ѻ9J,j�I�1�<1c��5�p�t���Rv%#{E��u��ts*~�8D��l$p��{����_�_c̺�i:i�����!�g��Y%��Č�v�
��P�ZyMG�3�������m'Y3����uo��E^홆c)��X��3����9"/y(�΃-�M�d�5v k��ȿ|#&c�n'�SV��U�M6_ϋ!,�F^WT	xu
�zV�4L46�I"v������^�Z��+��Rk@���Mh�ހC-�*3uR�����]<%��;�T:�ほ
�s2PQ<K9�������+I�ʩ��G��XZK�[�V��G$W/~��X�0�@}���fTp?k�P �
�E��2lY�?M���B��`��V�Kҵѥ/OVU��3�}�X���J�ݤ5��tZb�Au�=ѵ�-_ v�1cK�G~f��9?�,����;�G{	a�_�=BBI�U㘔d/� �/�
0��l��F5_Q�k��C+�z�1~�"�6E���x���j����]�m�뉚�b����Esi�U1w�Il5U�\#PZ�|g����<�����U�?��!�VC�R�[ft�y�)?2K�~l����7Z���҉r�Si�,���O.��uؘ���((��:N%����J2.Ҩ]�n�ф4_9Nfa�)yBQ�v�2K#U8{W$�.��S��7�2��O@:�|w�|UY&I�(��*��]�Ǖ��%�z�[ya�f)���B]uye��"�����[�HT/g+���a��\�\Æ��M:�{&���
_/�R������7��s�����+cH��Y�9
�f}Qa�j�l��ߖ�g�g��!�=�g	~�T��R�$��F���C�M�.&:�:�r6{7�9��!j ���J��o�pH=3�Wx���NeyC��,ԉ1�n,7BFiV@00ZZS�d&�� 	|gI��skğ֙�q�oĥ��L?�y���֯�������_��d�vZS~��CxVI޹۞��J�r�gN�vwQy"�2�p:�~���F��n�]� nE�ܰ\E4p��k�0����ci��`���#Y�Il�ka�t����i� ��%�j6��*c��pqS���P�wE�y"m�������٣�!Ռ4������	�,0��Q�27d&O>M�-#X��f%ɣB�_���\�y�9��|٘y����FZJ?x fHzD*�|��Uc�Dz=L�a�{��BmJ�Pn喇�m��;Xt�7$ɩQ�]�S�x�:L_���0���`Z�C���tZ��C!��/�ْv;N�s.
���U42r2�KB/�~�5���K��0^�	g��B�xC"G]��d�q�q����f�ɮ(i�_F�+=r~(G�vs�,-X緛8�*EH2o��'A�����p����Rn�1XI*��#G��f>�o����"YδϬ{��c��)oX(�������M��)�h��ʺŃ�]#h���pX�������=�x�^x� 7������(�V�`4�9�kD�<)��j�H�C�3��0��O(��� u