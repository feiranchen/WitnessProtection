��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
����F��':�ޜ�2̼ߵ2D�c�k	�?��lK���ګ�6�6K���}^��xF�u��hkp;���j�n���WVܫ� ����c������jɭ�L�5}��>��<L�=l{��	�Q�D�\V�d�s�囏���Qz��
2W6�ol��hX�| �/�������`����g%���9���/Y�ځD��uy��bPInb� �Zq����a��!���!����[3Z��{��0B�}���K9o�T�p��Zl�$r���^P�Uh���6��[�k(�3�~����NR)1���Nj*�:N>���y�5��-w��z��4�j�*HmĪ���/T��4��{.��*٘S"@'��A�4�Fa;hn��߸ň�Z�榧�m8d-�5ѻ�M�aSR4�����B�wOX*�2$��v'�T��V�C%�	���c�=��`a�0�f'�� �]�r�fb-]���Q���*y�i࿲l�=m�����R-�ĲXB���<0��\��KT��jEKL����D��4;�9
��}��n�L�2�C�o��B��LO CE�C}�gq�.��5�d�J�1��.���0�s�3<\���d%�/^� 2���o� ��M���������i��ﺶ�Fp����+�-0�q�0Yp�߀Fny����$1~>�)����m9^�sqѕ�ɽ��I�e\�g�I{����NoBS}�HX�e\��0]�X�yw$�~�<|m͐�����F��H�M|�_�!���/��*n�m��c�);��G9D?%(�4��e=�ޑX�Ra =��F�jA�S �Y����.fr$#��.�����C�d��Z'yV2��>��'u�Ρ)EM��"����bn3�B���{y�wZۄ�5���Q��{$�E�5�Ё6~���o�&�bY���|)˩}�YJ�6CX�����a*�w��#�`D9�R=���j�o\:���YB��1� Z�xČ��jMƕ��-;���*/%mL�Ե�9A6�¿E_Ub���)�H�}��M[��?�-�l:Z��%�t���&�o ͌��[�����b���G��6�:�7��k�%7�a��� m�t+c�Ԓ0������L���`O��8Կ�P]��- �~:,�A+F�ќE� =m)$�9"���n���!�0 4�	����Ǯ����3Tx��zG�Kv͑Eí�v14�%cI�¤�����D�ps��.}2�d"I�QoBHsj�z�5�*�tIV����ʁ�g�1�)"{���1�؅�ǭ؅�{�1�x��p��TM;�g�z�5{��زY�+�k�CA*�A��4��@��.�U��r�G����Ĕ�
�i�G����k#��JҤޗL����wH���yJ|�t�yџ���~�a��%���9Jė���Ekm���00<�ڦ��2�w{�k&n��P�}�MR�j5�tJ˄'	ʊEq��"AS���_f��u/��pg��ؓ�Δ�r[�"�a�.A	�Q�~���U��7<�+3�M2�
[��{-n��Pd���h�5�x�8 (W���b�U�61 ˁ���{!��|QRZ�9f-��[�����*@�J�*�/#�����>CA�w�%������W�ae��Hޡ����V���H�5F!�k3��?����)�a�`��ZP�������R��1�ހt�Cz���I�ܐ[;�0��0w�޲L�m}��b乎��+��[��J6��
�4�s=���-Z��S ��0��X�������uɃ��� �,�<��ȳ����ʤ�w1�����2R��&�щ��ĳL5��~�W�R[d�$�9���)�  ���e���\6�9� [�)��q%�"�6�lP�y�I�G�ZL/#�4���)�(/:u/��S!3������nȇc�T���ڐ��x՜��'zi�긔[��M�U�Y\x���F������>(���F��V4�[�Tpa���L�+]ڑ�hj6}V��{M�^��X��f�C���BW4���26�is�;�6�+Ht�Yc��_^-�O��@MS9��`U1�M�<���E�2	qv����U��<��
���${�� ˨���b��^r�pվE%�c�;�C��ƅ�O%JIw����.pr�p�I���"�򮄂��[�!�w(Q���ϣq��l:T=۵�е�P��7�1~7v��k�.�o�LmBɼ����A��&RrK��[�ɛ/�����zYŎ���T���.����h��t��ّXdYd�ݧ{3K�`G�.��f��`.�j������������O���>���E[\AE^D����j��U�ݝ���6�>��Y'`NO�Z�5e1�Z~�u�'Z�g|)��c������F�0T��C��Zp�$}޶�>�b=.fy�XE:�hD��.8,\`�B�%��5s\��_�:R�zy���Ԙ�I��`t!|f6̕6ǀ�Tӽެ=�6���RU�<���<�}���N���ES�a0+���`�δ�!�'����o�̷bW]�1��w��g:��gQ=<��/�&C�����A>��uJ]J�����$(��B�c6������v��4G+J��H�Ȯ�P�Ӆ���F�Gycy�&�J���^weZD!B�0��A� �t�=�:�Ǜ�?��#��'�jj�.�RS�j�ێ���Z��K"��x������\��(ҖZİ���o�	�GyC�z�&�%.^�$����8�v���"peW�P�9{:��S�q���ui�빘�9��u��@xl��>H�VYv���{[��$F�Z�����2��k��%ny�lm�ZT� ���]ay����B�)�����]BR��Y���s��jn�J�������#�m^��yM9�o�'�k�2Y[QL�rُI�浬��Jh��XwC�w-b��n�FZ ㏴ ���)Q�yC�+\���ķs�^�4��L�HE���Q^����m�̖+���;�y&�,�~M��e�q�,ʝ��J(J}\\��Cq�G��#-~k�[�;3o^�w�_@���H"xEk)SW�,���5Sīp/D�.c����f��\��=A�hڪ�
ĺ����9��Xz�9�5�{���V���g��x�\����{���r���M��0:VݪM4P�3��,�@u�bm�r�Ol�(4�L�`AK}o�з`�:xO+���g8���e��=Tl�6?(�=�sS�+p��(��'��h�a���䐽P� 2
�O+����<�@c�_�Q�=
%^
;���]6?��c�J_���ND�fr��9���۵�� �<�*���oYdLz�~,��ְ
b�+��d�]1lL}t4|ޞ�`?��w��7�u��w����L��ѓƵ1�x�����ߓF����-&�ֈ���g���q�]U'�SO��r5&�^�`���_����_؃�,�u�)�mO�3�b��8q��Bdf�*Q'޸�7��΂�vq�,���l��t���5K�,��L����È�����̩�S)��^��n ݹ(.�X�֒�|�1-:@��k���	�Da4��(�c�q�GZ_uS����	+�6�U�;����~A��3l�C��.�x�;lC��ARG�.<���($iˎ�'M�R�U�[�\��y�O�#�޽z��AJ��j�����8�!��9̉�#t8o�^����%�!�;���%Kn@mq^�VI�g�5	�Z���4N�0xκ��оRð�+���DwMz���24g��	��x��vPCL��kUF-�����E=�V�ǝ���ҩ��N2�0bViŃ�Z/b�_�'o��hZ�]������ڏ�A��"�uk4|ٲ��99��#_7��6'CT�g�-�9��H���u��������ȭ��G&�r)���j'$gL�^��M�%EH��Bz�S�.b�`2�!	�γ}��f�S\S�ĄL����������DB%��C�xی�\e��@c��S���tl9 ��L�*-l6��^���g`����9���# e ���( �k��B�K$�"/��{�eD�K�3o]�g���QO�m�r��*������$&<�
8��M�����M�q%;h�!eYf*"�R�:rA��̟%G��Ǹ�D��=����H�y�O� >��\�aK�[��P��a��\���b|�|,���2a�u��;A;�=s=4u���k�[;�d:C�xj@�}Q���PX_3�2|b���q~D!�G����Јv{�e�C��s|�~�+�^�W�;�hq�j���V�sr�ױ7|L+��ݠ�o�T���rg�OW�Fo>������ٽ?!~.c�S�"6��`���;���t�2���Y��>O�3	t~e.:ڵĖ�ɐ�����Ϩb/*
Ȟ�;] ���Q0)�Q���)��W�,�2H�eϖ�)&��<���琣�B��2�ϰ@�2�Vٝ.���I��h� ��G��l.>�)y��+d�@�a��+���jc���I�E��9c7�)l��!la;oI'�U�eI4_"}g����8�\*'�&v�#Zk��,����o)�Ca�lJ0����r�Hz�̿]�;]K:�{Bk��x��.���8fo� ��KyD���v;�	Η�4;��|?��ұ��1��`>D�!G��8+ ���b����@��f!�ݯxg�諷u���@� �Wn�Ȃ�������g7�i�n�ٍ�� wpku�]���C�C�f���z�GF��P(0�jL�������ΜL������R��$�j���r����iK��~�&8ŇW����V�?��X'!�s������<;t�O��F�xS���oHrx1�$!xB.	8�M8ӟM���ӷ
�`U�!`LH�h������@q�V���Dd�ڛ��R�ڤSM�(%�Y��/`I3�
�:i�Ϲ�p�FCӟ�哕X�C�ЁNRc�ી�����O�.�C7�ow�BqA�_S
������]
"ʱ0s��Oڬ��V��>�A���a�]�ܑ\,�=��a�HY�y��K��KGM��45bK^��)�'�H�x�>r�ٱE��F�c��%�(~�C��8�eRKc=��r ��=����y�4)�t�aʘ�Mbvt�-I`�I�n���;<�43�#꟩o��An=��PbO�������wL��WR9���3�x��<�VڕD���$��.&��Q����M�� ��]a�P��]�HY���	�K؊��@;�	�"@�̌��m������\�G$e�����t�HiO@}��RmN�8�G]��l��/�y�Y�Y����@� w�@@i����0��2�������
�̖�{��D������a�vJ�V~B���QR���*�C����[�T2����G�
!3T}������3�˓s�%�epFN�
�}O���u���0m&�<IɆ�g]�h{mFg�&!a�?�,�NP����n4
'���z��I����D˓ܤ,.��EM�����nd���7TƇd3���`�x:�������w�kB�WU�UKA �#�$ҹ?�c�3���	{�s�h��M�,c��Ê�Rk��힖efd��OC��o�蘛mߠ�mby��b�P���=�z��Y����ĉ�t��D܈IԻ��r��6���������=
��� \,�@��~U� F�����jk�ǫ������*d�kQ")#�J�ۜ@Ѻ�`��9~��|���h�h����ږ�ν�0^�U��1,0;����E]#��Ϧ�${uE?Py��h�)�YB"�Q��8���"�e����<�v�����B��ar'���D�k�@���}1@�ҿў�/<��׫q��&��x��� GI��b�_�ӎ��@!�wH�~e�R�u�z�V��Q_�}��9�-	�"�0g9tqC^"߰���;����\؊�����;h�	�n;}
�F�҂�CL	bX��f�\=ev?�,��	7�VsUE��6�&��*�d�赡V��%�\���~_��������F���������Rd��
�������ʖ|��+�eR�V��o���V[|c�.���x���MhauV�騳�`X�2���r+�BU��}��e[�K�J["��{_[֘�ճ`�xqS½�T��{�k��JA�5�ber��پ�r�(c~�������e�r�rO"CG�Y��8�䏛��Bo�t��W7�l��n��%E�A�)4Ġv�y��ǎ7ǃp��uE�Z��I�-�P� T�H����q�$��)OlB�55�͟/vx�͙|vg,c,#t*��d��4�͍�"�Ӊ_�҅���΍ueL�z8c�4[ɻn|e}(�;�m|�bE�M�ٚф1�q���vl�o�4���m_n�@�p�Պ�N��EZ�P>��6j�a�qJB����%�w^/c����L ������K�����-��2�$���pxN���U=16�X�V{���︡��Iš�05f"L�����_M�S�����r^6B�E��w�Jm�#�dPv�*��>���*B�A~٫������{�XȖ���a��fԠ)����A ^�=�rA�L�d8��(v��%�~�f�^eG��qf�8�aV,���H/��|����FIaβ�vP֜Ql��Ո����A���`���[�|��lL-8A�"{Pz�6ג���MP�EkA�Tǂ;��_�V��]�kO�O�d\\��_�O����=o]��9���ʹ� X�5���{;��>)sL7�G�|1X�5V� ��Ѐ����L���3������vC+����Z�����\��)P+���i����;/٨��Օ��#7m��t��[B� L�9n��J��i-,��Ҍc/�șS�K�P�����I�w�<�����u�.#+��į�A]t�Wᇣ������i�rx]WMCoRM�'f�O���&m�c�+���8*�N��Me���"��Y���gV��W�Z��O�ƐJ���3{p�|�lb�C���u}pQts�ƋI��q�K["�13;������D�4�r�]w�L7�l�M\޾�݇F �p +R-�@� $.�h�,��k����㮝/u��f�F:`]�7?G���r[���z�������c^~�j�������Q���5��ҐN>^N�{i7�ĵ^,�U�����N�92s�\��6�*�ߍ3?�
FB|#G���'�Bd�%Ш����9]i�6�V�-Tm��W(�S���"�?83"`�%W�T�'�X������c�J�<;"X��h��w'�}	#��������pˎ�\�g2�Q�!�vA�����k����e��jD���s�ޑZ?˽Ms�K_U���(�-<�>�>��ܞus�X����?�(w�i='���<R���ɨ_Zh���]�����ka<%qUJ����ո%�]GMW��6��\��q��~^��99�=Fc$��T.��% �@)Q��B��'� �"	��q7G~[�����7��ˤq�q���}�Yׄ1��Ҽ�|�{z�5�_��f���'�aَ+ig������|��B͞3�ދSq�#�*��\d�ң���8��b�g�]���a�\��	&��-B7�@茛`q~�&CU=���v�)�A����K���6؞K����M�_������T�V��.�ַ��7gZ�%�h{K�p^��X:Fu-� ��F�p����L{a�q�ﵧS�]���v7XF��g'^�+X���@X�"|�lw������7t]⯭gIC��`��<}G���D���OձL�?���9����������[7'���c0�B;� ;���v�����^�@C$�Kg��|���}gbrY3VJ�Q��	z������ۍ������_��tlf��FD�U�#5�fa��Xl�V�ߤP����~?��r��S��K$d�i�����η�9���rHӹ��nOa�wcOĠ��>�b�W�w���=G�/���]�5f?�)��7C�CU�I��8�nd�/���k��|������lao��C,�|�B���;b���b;
��r"s�.�,g��#29�G�)��
t���>�s.��nIGJ��k�?��^�����p_5#�L�Q:� a�e�<��I��?�����ؽq \X�Õ3������UYK5Che?{RQ>�[{o��	3�k��	{G�=���g#k�P����N�wF̝��Ke�I�_8GK���|4�ҋ&;Ƒe��u���;��^D�(�-T���F~.c�=Al��Φ1j�4M���ur�ء�|Zb���B+�/ԡ�}P�C�,`F��4kr�7`P�=�s�k�{8�ã��~ԇoӞ�Փ��a���J3�>�f_��w�,�X�����ܑ\H=�kx���"ϊ��8_�u�ze$���n���.�2� �a4{H�9��+��2�L��ڈP-�}�Z�ZZ28���߸��d�b�5q��pQ�$t�٩'�AIC��/��+r�%)M�x��{6�*�8�7p;��l:� $��=��4R�D�c{�z����R�[��?=�o��K%���o�#�#�y`��I2cM��AV1zz���Y��7��L��4XU�K�Y3�UС˺>
�ʘ�+���)��&<˝�B,1��l�bԡڠ�KIMO)f@������Ch���S,��Gj�ĥ�y5l�4E���aY�Z��/��5��.T�u5f[���v^)0���?d';�},S�F�[oR��Fk�����w�Q��پ�:�M�-�ʀ�@�iT���P���KX�x��/�F��*���A�+���?f26r���Ã�Ƅ��2ewcT�n�����t��$�6�J��;Xn,f�y�'�8�6ײ#��vN��oȶ�0"���SL|\	sI��R��y�$R�K>�I�>��+�"��`G�\Mws������u�r��ȼ�<��p¨��f^e��Ή	"0<��w v���Bz�k��#��o�̙��4�7\�	* N���Y]9�:��L��!cRO"@-����U���qn8��7��'��4� ~Y�V5h�!�6���UG��hP������7f�Le���P���W����B��DJ�;�2��)1ˀ�{!�Wr{�S�{06U�7��`^�.�$س��t�b��^>����W��Շ��d@�c/R
VT�aq�vwl�O���k�������rES�Q8�}�i��\�����	>_{��
W�U�U-h�<ݚ�^8\<x^���Hmq\}�{JT8$��(,J��X2�8�tԺd5bLO��_�I�̰H�R�J�v�`��p"
���ҍ��`P�k��N<��B�߈�XO�#��~՞�d��S��E�n"NO��s�����<��m���L�_`Y�Bb�<hn)M������.j��p�	�7 �������jf��  >sr�~�����������b�=�������-5��������N颞9?n�M}� �K���a�m�ݐ�Y2��QXbt��Un����]3BҼ��&��:2�4�b[�&��:Gˢ�!����}ńg���i�O	!0HE�ϡ�7_�V�
5��!��g� =ΕS��#D���XC�6eXl����m��Ga	�Q*#�0zk�RbSj���>��)�a��0WTD�|�������p�{��"z7�}J��=9��	ܩ�R@�ϓ�t�w�>Y�B0���Ҹ/�Ѕ�g�'gY<����$����ֈ몯���� ��0�4���=�o�#�]"���"(�/���)Q��S�J����Y׸�v������%�CuFʄ���͎�+���6�RE�u�m���xX��Pц��4U��Z��<1�����	l�趨֦�f������B=b軤��"D��Zn�w.�ID��Qъ5���bM��4L4�<t\�¤e��
�~�K�ߍ4��n~�*�lHcx]�T���P	�+�����}����k��\�������'���S�xL��ĬŘ��{�$E��25�ۂ��Ǣ�����aD�$F��4��f�m�  '������磆vi��M�qnmR��3I�({���ޙp�����C�.�Pl*�O��i-�
l<���j2�o�C�������mF��ر>(�;n�5��	kf��Jf�7����l!�P����-�Cu}[�OeSȜug{��-[�7��\u�[�j��H]�8�
�	zDl�;�<�AT��(!�n�:p\c�
���&"[h��q�Zi�Y�1ѩ)%|H~�F��X)�<����$���%RCJ�|��=�cX�}�_X�3r�Ew�A��h�j�}���%98M��s���I�)#+\?����I�Y����(�-�z�,��"(�.o/%I�q���&SN���켁-O
�w�ck����e}�*��q�r�-�e����@A���̧Mr���SQ��3b��I�C;�є�&�i���1�1k�)�eA�*_%�a�ϛ�7���z�x?���
<�l�*f��:��V�]y\�ҿ@f�ekX�����>fj(� �(�_Rۻ�K2f�֮MP�+�A?��h)����h��o.��x��΍