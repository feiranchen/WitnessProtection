��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�O��?A~'�}�6�xbR�v���m�r�K����n�y��P*шu���4I}��`_�����$��d�H�ِ� s��Y���<�N��D�IS*@gH @n�<3|A�]h�����;�g��Կ��=��Es�0�{9EW��Y�9��[
wςh��7Q^���������5Z��'B�:�&�L6�W�K�o��f��kL�}��:��RLQ�Kw=qS��kv'�]�H7��G�.*L����Dx�g�k)�5kw�Jy������z�����q��eg���ݽ �1W9/:{b��̣��f��(,>�Tv�	���!�rċ�tsqː���.���V�<$:��u�P3���*+^>���t[O�y������9�CtP���� cr�qk�&���I0FY8њ�=e��������M���]��/:4�:&���v�U>�Þg��a�h(iL�A0c���}O63�Th0>`�6v(wF�I!�9ACԞR? �%A:��)��qUZjk���	�0/�-��"ތ�י�IԌ��^ԫ -ғ+��Z'�����m��,�_<�a�h��w�)�̆K��������?k���F{O���N��l���H���DL�xk��]3e/һ�8��w�{����?c�jjW}ml��U0D��<�
}�m���4�#�:z�j�nz3x��??"�_K b��Y_ַ9������H�ēZ�X6-̑��փ�&�"��}�Z^%%}і-���G�.�йA~Dٯ�HH��l��g�~��@'�7��<`�<6��৏O�ah'�o�J˚� ��_>��y���w��rp�ADL~cS���a�9�b����FaN��d��t�	����-`>�.q�]n�Հƨ
\�wah���gڮ2N��ُS�8�s���%
�s�}v��L˘����UDY=���CN �x�7�Xse��Y�)����N7�@��\���SWG�󞒶�&�0��q_��CC�"I��aFJ[OQ��FZp����|��^{E+@��"�:�3۴��@����
L��h�[ ʛ���
��d�>>'�  �q�������{r�� �.�uXtl7���)<�n��GB��a=~�"L:���m�36�����ʳ�1+� ��?��֚֎ ���D��٭ kh5�<	���-��
gI+#¡�1����d�3[� �z���*q�Sl݊Q�Vw9T���Ħ)�ૠ��n:���inǝ�28�0��߭�j��,�K�<����7*�0n+z����]e��`�IAM��x������Ð�������`��Gm ��rUw��]��b����E��f�鯒�K�E9���g���G3ޏ��{���B0�{_�k�F-���-�����|�H��j5��J=�`ZC&>��V�{��'��)j�vρ�߇�q��ى;��N�?���󏨿Vr����C��Q��7���t]Y跤��o�������0�]~_�`�T",�>���;:�Vq715e@֯���{`ҹݯ�f�$�,bt��䵬�ovIT��oB�w����@k͠��V*,A�eǃ��'�=�^�Ip��{11��4/3��p�\���׶�2������8���Xkk� yz?��(�\��c��~� �V��ߴ��j��qI��^2�{���Wt�Br��F� �x����j�� �U���m�^F��,B�i�L�}�W�he�q���{�����I�à޻v��m�o8x$�����!Q(R�.�U�˶"k�E�� *�z�f�;�X�:�
����h@oZL$�' m���#N�����횟"�a����K9��%6�#�%��αTB�Xh5�����(�
ŽNz	����ݭ�h�.K������m"p� ��^@9�nmVd8��..�k�������pMm��g�O���UcV�ؼ	둤�7w�9��ݮۣ��X��1OX�N��W�ҹ�K��l�
�fإ7��s'=�h����^�|���K�҈b��);3�������N�Y��+~��	KG�ᇏ�a�6*��☮H���)8#��|P[|4�+^��6a�>��-���~}��@�D=�R���4�AH���gF���}OI�����OO��[�B��O�t�4. pZ0�hd�h~�7ȉ�l��R-��|�CB��UJo�q��V���o,�@��zP��9���a�YW���4�c��Z	�5�Y��Rrq�˿-3�j,���XU��Ǻ�Տ�B||�
1���+�ZΨ�<=��9S�����K���[�vŴ`���Dd�2�}9��m+���e�ݫX��w=z8���\H�l�tS)(�T���v��D��zOfBx�^"�ɹI�'n�7$��7�y��^	A�@�`^��1U�`�0����
ğ����l`h�nU�4=�꛴M	�p"��<�����~��g)3L�W
�x�Y?W�Z�1��祀�[jMn|�x?�����[���`��9P�1d] Kg�\�9�_���Z��UR�*1�yrAy����5��e��k�V9��_�o��'\��j���:-p��s�m��ZȻ���U�Ps�Fq�u��0b�1�_\+)�y+,k��\�!3����M���C9 �L"l!� I��;g!K�ku8�����e�%�V�E�"�Ϩ�;��S�l1��R"9L���E5�W���'�N���� /L��>t6mD�K������H�q_��	��iP�K5�n���T*jWjU��c�R�4��b���`<#F���Y�&\��I����*�Zy��
�b0�5�48p�%mG3�M��P�q=[v�,�����(�*p@�\=�tf"��ӧ;r77k]��(�Vc���k�ݳ��W����� ��ߙYa��?>g�q~��Go�,��<��k���p�����jl�En��Nq#YH��JC%ad
��������D��62T��A`*!=�M$
<���r�H<R�WI��n{���mr���L��u����C3�ՔSs#̧̭߯6�b,���!��D��-�/u������Y�xf�3��x�k�u����{.����2�9>W�����kLK�d���Jbk�<�$%��;�� J�{��T%�%����U�C̙q5�&�ߗ��#�s��-�)]ځ���s���	���xf�F"i�ɾ��d	\�K\n׏�^�Tm~�&��X�Ae/^E�x��<Y�]E�>>?7:�b�ڗ_�Kt�o�a��*��Oq�s�w�������i��xv+$�V��"m���ͧ�$����w8I��;}����r8KC�WvU����7�0z�&iYr��4,W�U��Q.�([��Wi
�e���L��*S�۩�*�e�\�&�&�� ��P��4��}:�VD��T�ȕ��s���:�8g�:�Y������Ƀ���~�QN����ن] �g�ɤ𞐻mH���4�IƆlBψ�-[J��)^_�k!A����2�H��L�+�x�i:{}�(�!S+@���݈��ʛ&�}�^�F������'��5A{`ꚞ�|��߉]��~|!�M<�y�repo݃�m=�N�̏���S	}C��O��{���o<B?����[^6����W����@|�E��}�@\֚�8���61I�a���YZr�ִ���t�&#m8]�aV�X��Л�m�4��S�OO�{�v�M��e�D������ 
��Q��Β���m�&2��f"Ef
 <�؅����,�|�ϲ�Oh�k`�l�����Po��z�ݛ4���Ɓ30z��Bk��Э�W��I������͇L��̢��Y�.d_Ҧd���Mt͞����������:&�6ڷ�O�Hq��R��-�.�cg�#�0���ʠ���KI\>W���EM�mbT���{ �g����~���Su��G���������4�`uvz���,*#Z�8찯A��׬����BM�Z����@�xyp.�i�l������˅���*'�U�%L��� ���NˏTU
�5��2 �p0�m�����<ן������ !4��1]�p�,4�����&P�����:�.h��2j���`����7nwy[�P�+V�����
+��j���P_���]�O�Y����N���m�wKUz�_g�r���812����`�w�L���m�l�ɲ��F@z��v��=^zT���iS1�BP�&� ���*GL�	U�ItXx��/�N�n�w~��W������AJ$aE���D=��(�|}PW5��wc�qŃ���b�/��� ��@�Eb�|Ꮾ�c.��������M2@�lĺO����a1��qg��зxytK}�"�q���k�Y�$�"��H���_�X�u��2T%�l ���U���M0[\&�.�i[�p��d���4s�	ӯ��e$��{�&A�Y����ڙ�R�,֜RG�ǝz�"����-����jjnɄk0{�RszXw0>kYBz9s����[�~n9��}��]l"��1��F������"�s>���=�/ F�:y_�Ƥ%���}N�Z1l`[�f� �|���"�7%����؇]jg�������P3Y��jX�#�W$5
���7��.Yl!�ҹ���r|,ѱ���"��gX�&�FBx�}۟m@a�4�ܠ��px+��`g>wk'	g=I�8�ϼ*ܵ�h�|Tֹ�(���;%f��O�=���R*5�=Fsp��G ���#����P���D��!���&��B,�fkV<;>V���+�@��i�c��MO��H��,�b8P��������RB��v|���s����X�&@�(`êw�����Ɏij�����c��5;p��?
��m��\�C��W�A�H��E!T��1�%��&�m-�Ls�ؽ����BJQ m�9��=�gS�7�H� ��1�u=�����yf�=�?>aD��f��b��/� +X��.��K��n���<�P}K���y��0Un$�5E��ĹV~�"��&%���ܣ/� �v��/6�w��Y�����Je
,	/p��h*K�BsB�(L��ܵ7��Xg.D��;���^����΃"}t���k�=��ʹ��� ���")9�lx���G�>��<��s?�7��v\nCc���]Y'ڼ���We)F{-��6����0�{Z�y���su��,������ �v��c��Z)��7J�!&ԟrKRЏ�J$��b��ځƐdz?�����2<�ч���r��٨X`󑉢̈́5B��W��R����[(5n7,-��Nh�n�륱R}JC�
�M����9c�7�h����L�@Ҫ���?��7����d(��	�^b2�0iS&X�'�����Q������9L��bQ�%�Y�*�g�������C�8�!\J*^t\�!O��k�ɡ�ֹ��ba[��3����5�7q��3�Q�h]�r�4��S濯b�9Ҷm7����mÊJ'�D�+�8��y�k�Փ� ہ�3��@��Zi6�6�AKn�I#��J���p���2���d�3��W=�=?�q	��t� ��N]
7�yb�z�,Kz~���(��xMW����H��f���	'�����-!Z_���~�fë.5��W�r����� ��� �nӓL	o��qL��5�?�Q�қо/WF������?~���׷������>�&y�´�e�Vmh�kfs���q�?�F6o�V�8�JP�n�;���Y�e��_�8.!�^T��Y�SY|����|G iUL+�u�f��o�/bB���لV�"�X��!k���J�s[�����k5�Yy�;^RHEx,Jf4.���Z䤵�����Z����휅k�$λ~��S�"'Ŕ��- �[�)���z�k���"��5�e*��>���
^h�*0�{���"�OŜh�mj��C�F�Р�Fܷu�������@^����d�8��Fѭ�!hO}h[�.m7)ԓTt�Φ�<���FF4��jk��v;R���2��H�GtE�P�W�X�$�����<bR�}cH�B��9����!?�ZozS,��ԭ�Z�:4�"sK)���2!��b������E5pw�'@���x���"z��TY����r���}s�4�K�6p��z�y�б�Jn��U�4���&��@�����[�a,���/��C��.焅]� Ŝ�L)���@s��"F:N����V�`��П�������ͳ���V����xWdY�a����ɣ-�����ot��	�w�ꈾ_l��Ͻ�\��dL@�4���0Z`����['cmr��g��9��:�/�ͯs�4>R�|J8��H�ĊI��W��b�2�O�}��I�_�h�J�)��k��~��7��ֺ�ɏ��f ,�M����mRk�qܹq�#�PH���y��󫩝M�S�]؆��.�L��������5�J��1XShZ�N�����x�"��k��� ��s]?�䂃¡L\-���ɏ.�k�g?B��{�WK���\��G�@Űy�h|V�o����
��ْ�w�M��ARF�*^�g%�e���X�"�*�mu�#�]ߍt1����a���_o�YL:eX5֥��'bW�
Z`k�_��wF�� dK,����FW���&���C�E?��Wh[�폧ՍX����� �iYI�6��= :LI��&\���z��o9������n�2���.�H����`�c��& f��`�Q�Z�MG�$��n!*{�=�^��0�����:�-�������n�����k�2?�o����<�$�q@i��t��>��^�A���}������v����3�M�&�h��[��LTw��I Yd;k+�3���=mߏ&�ñc;u���w;M��Am���h)��m��X��������6Oj0b�0��@��jY���*A <�������/=���I6���!IW�
>��qۜ�pdg�F�1D�qz�3���򵀴�_�&#Zu�v��-Q��rv��иk��:U!�>�`��u��;mz�ݫ!��E[u)=�Ȁek��l
#��,|y��-G0u-��'���YB�z#��d���Su��F�w ����b�D��[���W��"�s�[qP���J@41���%g4� �_���`{c���2����%�t�(^.:�C� .�V�T�A�2z&`>�KF�a���줞@��"/��8^m}R��]�[%*��Y�z�~��v��f�=ZP�&@R�do�YqZ@g����$>#�\�����[/�f�G�d�������Z�6��+Cq%�;�hf6�c��K�X�@����5�m�����N�C)#j��9�J��I��,�ij(f�P�ŔiU�仠�z_,ɚ䲩����d|^]�6�LE���f������ծU�vޣwRg��&�n0,�GtS:G�(`7I��u�D��#����zA�9��6���Ւ�U�ԛ.�*�1��p%9�!E�Fo[�9����k�78´����74�бw����~���q���v�������V.�\&��+R�c�Q���{P���݊p20���e�\a%U �,-��[O��pe+O�!5f�w�~xA��}^V#~�	��.���+VB�;�[H����Ѯ�}j�� S���"jcBR�1 ��|4l�!�w.�[�գ߲zp�y�.�5�׈!�t��K�#��*s�ͬ3��m��/�<|�`��|��,��w1Đ
��~a;�x��u*L�T"�fr�cJ ��K;_;<�1O��j{AK�τ͠�뵭[���`Jb�-~�����a21��s�bq�Zҵ�$��m�XRQ���Ò�nY_�ݲkH<��Eyu�V�ڦ%;^�ۮ8?;q[]�O*X��B�l�>(s��s��U��rxV����#bR�a1.ˡ���}I����)��YZ�34FQ����l"��G���vu^j���A����xl���CT����+����H��������_�=G�js�#�[v�<���f
~
=}�2~f�����ݮ�dG��[XM1߰�,�Y� �/R2F�kI�Qq,����;�i~��$�ǐ#t	y��)�Z��}���f#s�-���M��ނ�PI����D�y�\��@�Xk�h�7��A�.��V�e���<[�Сҽtf~�8!��N�W����ڵ��`x3/<H�Ү��p�_���x1=�[��l��lÒr��ZY<�ώWtY[Z7`N��`iǹ����#'�D=�VE-2����̧Y����P�"�Dw���4f?l/�.�3`�N�4l ?g���c~`�R���ʙm%D}��}����j�&+F�d�j}u��j�΂s����0Y�I<��u9�bSJޥ�F\&�k��eg�����R��/�+繒g����"�!��u|x0 �M&B�"���X�_���r����/�H��l2զ�m�
+��>�?2dwqjUE�T���n�v:֎]�x�F�p�A=����(��&��v��+�pP��Ns��iŴ�$���d���w�:%2�4~�8�裯� �kdk�|D��g�I�E��9uA�?����@6����'��	�D_p*���L0�t�%���W�[��X�B�����RK �[�:�Z��)(�^Jr`�������S;�B�"�7��H ������}��WH�{�Δ,&�H�^Bs�� ���w�( ���G�����w�1��cl� û��nƽ�%#L�-K�_��p��u�E�j2tB��hŏ)=+>�B��fE'd�xj�5o��?��."̟&�K�8p���Go�;Ve|5s�+��=�B⻆, ��ܲt�w	P�c	��ne]Ũ,x�b}��#����m:���D� �mCQ�<{�kV2�s�a;ύ�=��7��vB��m �5�%��@�&u������8n7{@-B�$7(���?58#������ZŶ�R[p����K�07>uߥ-E���+��-;P�=� (�s0Gj���C��nֶ?/�s�5�y:�ݿ����]#r@�WH W�T�gEb2�kE���G�\ .ޕc-�t��j0�[k�-�]j����㿦u��em��Ew,�Cc�a�H#E�6ϕ�[ޑ���n]��G7�8�~��$�X�U��uź٧��B���@v�Θ��O���F��b:�&��g���޲4ཱྀ��瀄����0�9�6&�DS�l,���� '0�9dȹ4�>3���z=cS��P���ǐO��H�������J����N׻-�zq����	�����~2`�.r��cg ��p��xq#�0w�	�Æ�s��	�=g ��͒*r�q~v����npM�2O-�Щ���hLY���|���>�(/���kHgI���n҂��>[�����v�3�1������f�I��@�%��4�1�m($��@:F�0q3�q��Y�2/���޸`ߦ"��@�Cd/�W��F��t����I<��[��������_�s�\3U���v��ଗ�3|�n\�WM�#���E�!���/]�/(��w2�$��pC2�G�	\r�}�sW���7n@���,lH��q��AJNm|�����b��K/�❧=�)� �E< "j��H�h����x�6�s;�s^Q���c���ɚ�$m�8S^�GI`� 8zӍ�h,`B�<먅qD���a�ӋE�EOW 7�٢�3���%(ZFɩ��n]��H�G>]�is�77��z����/�{�Y�����nq���#n\)��M[���<Gz� �N�z@�Sx��*ѵЭ��C?Pک����+IԸ�3Bo놟C;�W�<���j�tv���mۮ�Z����O@�m��^y�D�����w�OQ�#�-�V�wߙ�qAD��Q�h�&dq\fk�L�A�B��j��B�#���R~ֆ!}Q,��:�yu��h48���|��8,��|�A���˥�˛�\���9ї� �_���JI�_��<צ���}X�Oܱ��P/`0�!�-�������㏂��ۈ��4�E1D �N��*1/�R�t�䀨�_іp�iȠ�@?n��ܙ|�F&jba�%��V��  �����?a=zJ�6:�%G�l