��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7X,��8KI6E�2�
������V11X��b��v�չ�+'��Ѫ����a�����x�hiP���Ȧ8 �'�X9�rԜ^	D�n/�#X.�nQ�LgTx!�xf���E~̕�� �0�'z�x�]驏)]�9���d0CUT)�8L�m��f1Ò����1}���C}�ޔ��h���Rkg���M�=]��ʖ�%�����qi,�oY�r��	bbo+_j|-��%�����4g���("���^�oJ2樒�exੁ�7&�q%h����{��nRd�[�ѧ7�d$J�6,��Qs|/F,���!Q�`r�������*9H�$��ӂËi����&r�s�s �]��?MV�lĖ]��=4a *�Os���E�~��hC���F'�r{1J�cQ�ʳR��C��?��An��N�.��!�ʃ�0��Fu�ϙaI�sp��7U��Yp��\-�,�p���46�Lۻ��L4�.���*�qg�eL�el35D�ʫ]���\��N�V!�=�����J�T�mٗ�t��K%0�e���=~���UekR��f?�.����L]mɹ�����n%��Y���������P�1���R��"Q/����`0��V��VSi����3�͜�E�E���F8)?Xg��=�����Ɛ@����B�sI�+��!��MWƔ�
��y|7S?`�/5��=r�	��B�6q�l<�W�\9s����'����maz�A,G������d���Pw!-."�/4}r��V6���pPp�a��U�s��#8&	���\	29�r�\��媄��f-O����<���t!g»:m�� �)e����9���1@3��za�"�����J��yK1�F�o�ުEcoN�����^�c�W�w�7����������9|<�%�P����&���]����zv�G^�J�����r�U�OZ�м�s{��@bI���4�V�(%P�����/8*g2�'�$Ձ�`��4���w�������b=>ޜ�B�\��[Ƭ�+;9�g�x,A&�����`�Ww��8���(��xJ<UO�69 �ٜ0L߈�/��b*r��8��a�:�^�%	YWo��WP�NV��sf���/p�3����<��B$q'�1��պ`%?<~�HpX[»�C �(C�A2�9�%��:_�gV����YU��Mn�e�d�uls�@#u�@��x~v�� �h*D�ޖ�������h�������C�&�T����J�L�tF�S�{�?��χ�/�(�#ԫ-��}�r�M������?5�Y���籒�3�f�� �u�sJ���'��8��n���U�4J�C�4�R���ѻT��d�	�
&ب���ڬ�H��	\���<�y���`�6m�SZ�ہsC���'���B|�-w����ֿ�8��+�P�P��;̈́�Yc�I4c��� jcX�EE�.�R���H�w��[ ض� �P���4�M�\b_�A�Uv�N��e\�Pv0ȳ���J��8b�p-�8�!��*��g��<�M��w�z�
%�R�O�����m�ě?Xj����
�U���k�oԡ���b6���.ӺR��o@pn�]�5�yn����ʹO5ٱ�֋��q�zn��[[؈���m�ғᤉ,+�ލ"o��K����<��!�����瀨28U��t�G#�Z���d��m�S���.y�+N�?=�s�n,�Y�u9�PmVZ����*��yC8�˞ܪ�[x��,7�]���Q�=Q��u�q�v��}ȫ ��}��5�*!�g�%�w#m��;m�[a����g�Li��Av��v�ϣL�M�C��͠�p�� ��%J,��0��J�D��d.7C>=�s���Jl����nhta �dP|߂��((Y����&����*���&N��A��0�*��>P�)��T���������d�t�S�ab�E�U_f��1w��T�Yf������W<kW���q)���pخ�Gl��h��ؙ-p������zk���K����P�����	~ü�sl�>��#2{L��sF��D
P��wr����I�͑��e����B�r�mU;U���h_���wp��g��4�ەd���o���p�5�'ι������� _�R��) f��q�8��Y�����{��B����K���Kȩͣ���dE�;����{T,��Ν��!����y*G5��^Gm�o�o��!�A�UEqt����[�Pq���@x5�Yv����Ph��9�3Ѡ�pǻ�h}�"&B,���fz'���mH��VQ8�g�T/g�e��S�Ң�ͦX��r�:���ì�M����<n�����0�P��/���1+a�1ؘ�I��g��!�6u�;QW�4]�h�����q�H֓(���8F�7���W�=ZC��vO�p8-#�B��"' �n[X�XqakJ}�8/^�K�8rUS����
�;u�����O��h����H�5����,��	����'��o�j'���=��pX㲔����B�޲�JF�J���  ��HG-����,���ᄹe�k�hԎB�J�$��W`����n?��^]N�h�?����T1�"+UȦnp�8�)uD�����
#8$G
z���*��(��l6P�c�~7�&4�T�GW).���$P~4�a��Ǡ+֐o��{�r�.��j�Ծ 4�&I����|9�����&���N���Z��g�됄m{�Q&��]ͼ�������wŒAC%���s����_M)�Ǌ7؞���+���A
8X/�F
�d�r�"�^h�āƽnױ^�����Ǟ���ඓ��i]?@�b�� %�.7\|2ǖ�gG�4,�j_��'5���/�^^�h�`6҂�	KH^�ӌ%�~Tj�z�~0�e,���	M���W�.�.�pn��.&�dőF
��NV^lD�f]���M!�}�:7�M�q*�\M.-#�G�	�XD>�Ȏ����8�Dp�!_�s̄����A����yǓ��ګرS��SC��kM�R����Ȋ8�Lu��T�Z[�L���v*��|LR���$i��ME�%ٖ���@��Oh_�� �N�b cv%���I�R�6�[�s�i'�7��o]�&qi>iL���f[������ 丒����e�K�|�QDU_%	EW�Μ�9��W���w������J������͔�O!;���:7��w����̐p��*@�p��3�|� Yj/���(���3쥝z�|V�~�`��ڲ��a��(J+�f^M}�A���m�����R��f@����%c@�Qh���h���`�*�g�!��4�°R�U���s�W�Q��W`��~%&s^6@����8���Q�'G�'�@��ߞ2U#����������+���:L������cND'�#ڠ���Az��5��d�ɜ~�4y���.�5M����,_Up�)��HB� �W(�q�.Y�6+ɵ��|��:}!ۘ˘���C�>ş�n��搠�r�f���D����t�Q �?��B5YD�s�3���&d5:����W^}��:�����0���^,{�0{�%��8������R���*�=�^��6g����*�ܫ&���2�W���3��$�I�t��)l�ya�T8��=�]����"Y?"�V�L��	oMt��2��~���K'ݠf�ٴ�q��X�ak��ڗ�z�C�~�7z�B��m�Q`����b΀,���?����]�N�-��ƙ�&�+B�P�}%x�8�-��3X���¡v���n�
�����q Nf���mX6���������Tl1s��\��Y�L���~��1���g������o)�ʚ�8�x��D��W�Ш����U���D�ͷN"��#`�k���
X[�0�J���1}'(?@O�u{߽��%�a%����^>a�/X-��m��r��tS�˓�����18�1�����&X$�M���>�^�l���)÷ϒ!3}����[�֤oM�8���%{B�{0W�3���-JV^�u�W�����(��a�#}�^x�p??��%�J����0����͢h�����c�[T�o���Z��n��Z/a�4o�*d�"ޡ�q��N� ��1]\/�%�M�� �_c�ȗ������HH��R��!�]�,�Qd��pLc������1�[5m5���Д��V@Y�>.����vԸ�J3(?G����I��U����:V����$I�bأ�dB����۵��`��E�¸�Pڃ��qy�C�/p�l[�aQ�6\V���뺧�0��6����E�?��Ը�F	F��~|�K�!��m!�W���[��wX+�rۥ��u~ �δ��h^s�K	���u�db�FJ=��«3�����*�.�3{kᚭ���K`��գ8��G�����ѷrhf1���wq������3ə�c��b����G���9�Q���α��C�lg�݋EN�n	��4���Z���b�e�ӊ�p��hȟ5�@s��?�Y�A8VQa4��T�"5�РY�*µ�J�s��E2��)�~���a�
c�)~Ns�����c�� 1���9���+t�};���+�
*�N�ɐ_z��/��6�ۜ;�ܕu�@T�='���0řf�!��˔�́E�