��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d!z��� �vD�����?�gIp7��P 8���%)=:ϣddǝj����.�����{�`o0A�~�L&�{����`��6e:���W��ӥ����5/M�^��+ϵ��^��%^�F�6*v�����u*���b��`d��-l�Ņݪ���UFNř���}��.j,�e�� D�ǉ�$�8�R+���}�)�ΰq,D>�$�-otJe}4a����J��j�`1(۳�w����E�DE=�],��A�cF��M/r�����g��S
O���P�.]�BhwF >ju�9h-��l���#��eo�������HaV�s�e~�Q�5
�����k��:2���5r���<��)N�����b�B���d���6:�Y��U��ќ���Ė>���KT`e۾��I�ive`�xF%K�ѓih��W+Ӊ���4�O�bL�!78ؗ
e�٦�N�����փ��Ltf�ש�����L*b|�}+�b3����
kVTH�?^�y$V��g/�̀���(��x��7,=�4�$�S~�ͦ����q��G����I�"qo=����E�\�����
��/�g���9Aȉ���(zg�c�� ��Xy��`��28%�WBR�ρuL���F&6��Y�05����k`�	R����ޛ�]i|�g��ڐD�J��T���b>��[Tb��y;�-�dθTH�>R�3�l2@�BN}fa����1�
�BZ�95� B��WjeW�b;_1��M	����m��L[[�v���@�Ԇ�	!;�Z$�`�)�6v����g.���hDI������ѷ=HN�lӍ�`�rB)�؀g�L�� �Z�~��H����KIj�zUHjC��=��x�"�g�|D���fL��"���ʶ(��O_^x�2���ޓI��U� :� ��k�w�Wg!�� ��^�����z:#������%T�8�����K��r{rD�N��w���x�q!x��HԶy$ ����Nq��>_�,j~ݍ��󜂱�4�*�AAKl�u{�t�Nő�D�$�j{�gjߓ�?;�nt�%�~!Z��#�V�0WN
	��"��#[^�@7����\9�lA �^U�L������<����ˤ>�E�C�F"�8� n����D��W�.�� ����2����?fT�?�Ӊ��q ��Z�T{�Mu+��y쎶�e�)�e<��NK�'���#�&�ru�*Ru���� t��-X��A��/�N�d�bs�'pt9]��@��r�x�۵
�-y8��Z_�(5��ڣ�v8�����:�8z|��6�5ɘbgy��>ƶ$
�/�aP�[��lUw����,���#&��͗h�$66�N�ĕ��@��[�py2��ɣ�=SZ�D�=)��l���^*���%�YJ��i��#o�s׸�24�.Z�4��*���c5��8:G��f������'i�hǠ\x9�� �q���K������Qi �en�U�(�Ab�
6c�o)v�3=S�7\�T��!�|���oOU�k!^~Q�-y��Ì?�(��g�麗Fq��S�zQ(����).�J��Rh�=@�KQo��Ƣ���yQ5��7�.�B1w�B@l&�Fv�B�t4F��MvfE̮���q�"f�LХa���!]�4�rQ��n,����dv�M)�s�JRu��^Ҫ��S���h}\0�;������IN�r��L�t��=�����|�_���ň�.ydObDprV 2�㮤�6���'����b�MS%T�QN�hv���ޞ�����[g���f˪����S��exF�������:���6�\������>ocEYkz�ұ�䘞�e�9��9���u{ /�b�hN%,r�����ݺ,?O����;����d6�Z�d�I;�gw8m-2S���������W��o��VK�˅�Z=K{1�}�B�G��-��>���3�G����O��!}S%2�K�s��gg`�m�	j�Q1��`
�/p�Lb0av$���}�u��5|��)�,�&Z�5�%�̺H�ɗ��AS�Q�m�R���Vw�\����BjU?e"<�,i#g����+��Y=9�臨�L�F䃱t�]`,�K®��$��� `����KgF��� u��pxO����E�f�֮���W6�mE���zvc
��Ń�#6����9�,G8�ߋ�Y������P�vG�+��#3,�Q�2zY6U<4�9'�p�I���)�{�e������\1�.�j]�a������]Ԇ�h���I���l(h>F'iyN��)g�YS��W�����8Ջ��F1���.Tx��#���m�e�;x/��]��$NQ$��I�@~���Ѣg7Ei5����5��<畭�m�Kn�s��4�<�6�;M�/5";b�'��f��#�JV�x;NdA���Nmn"c3A��M�w�~n�y�9֟`G�Y)�F��w�aգr���y�Y�|.%a�zU)�B�a>�ý%������o��hM����ٙP���P�C�15 :��+��[��r�M�y��ͧ��;F�;&���A��A�<�ڸ���+���U�m�A��Mȹ�T}A|���ʖ�^\-"GN�6}��J�TǮ�
�Ў4O� *a޶J9
ƻK+���JD|e�A�ξN�� �-��7S+��U{	�x2oŕ`7�ׂ�:k".�T�#���˓�.D\��F�4�����C,+�\C:���ۧ�.�,�MMڑ*���"t�EL��&�v��B��~�YG�'�D�cG_��9�۸��/&��R�3/W���XkwhC�辻�2��'��� �	$څO�:\ܥ�5?mm�>w��
��b�威~D�v?�K2.���ԗ�e��uM�9����ֺ�������I�f��s����j�������<�r�Y��낌q���#:�ߨ�=��a��A΃�U�Δ��&�%$�.�����od��hӚXs@P��/���3_�$����
-L��e��ǊW����2�R��14�V�O�C��&d8:����&黼�,Is6I'"
�@�	n%i���H}�	Ďk<Az_|������ ��BMIx�^k�a��}�������I��%��C���g���i�^�4*cZ�����$C\C�+���Ӊ��a��#Tw�����ˊ�ڎ�w���ו���ʔe�|I�<�����t�a�3O��=������z�!��r��Q[��Ql�pz}sw�Qny߼5��Pu?v11[�������Ȼ{���F�nu�L̪ /(o�݄5׌���r�^�K��)_�� (��Rv�H���>O�[���p~��9�������fO����Y�� zsJum���<�ɑ�M��؜&t�&Z	�]x>��ɣ�Bm)���ǔ	�w�R{k%"�"81＠�gM^L�*�MQ3W$����g���ޙ�� � J���Yp6���x@VȞ��|O�|�E*�qO�~j��r�Z�I{:���V��$ԧ �N�Y�6Oe���P���G%�_��wp�}�7�*ٍ��P�;�t�g���ԙ;�}��	���x@��ȃ{�Z�^^�4��WJp��W�	#'+�k��������T�h��t��
K�)En]6g����.�F���i ��ǆ����ne��/�D��{lKN';(�z��I��r�[�S�,=��{��ܽ�
%1�P�a2N?U��5Wy���@2�$�8�*}=xhƤ�	�j)N	���pAzq��1
�UR����Ű��@ ������<LN�k}ы��k���U<�K�)ҵ�|N��4��uː�;q���v�#P�q���\�X}+�	�(�s�<W'����"Wx@Ē�o䢰�����H`��r����]�Q:��z�=W�i!�� ���:�d���DA���]����X����*��.��6pZv�O�Pb�+E�l���?MpF!ִ����S;{���u`����;�,C��m��q�!�Y���E�!DZ�}�9?�g�U�!̥`A���p?=����7����_o�OL��lq��Kk��Ű�������'{z�s�Ȃ�����˶��G����2z]�Z�D����fM�q�C!���nb�#`6J
q�F�gU�C3��'�s�����
z�������~|��OJq�u�Fo�;%�����<>X�/[�2�n08c��5�n��"|'�Ҫ��T��Zzh��J�]��]�N�<4���	�V���?����ڎ�͈��%��Hj)�) �hc�:�8�W�
�
��+��;�Z�O ��}�}-�A)*E������Y�Hw̖��L%���������A�+z5�gu�>17ur�.�;��3������5Y�G���l��ɒ��xb�E�e5���s�2(�j��!�L�8G��%��h��^ߍ
�s�+��y��(j�����|5���� �y\��q���r��ݪP�����L����v�?��U�k�&o�w�툏���]�绊��uK�q��+��t"�h	��̈́t���{��3%��|%�36� �y�]�4��D�K)�An�q�.KDe�O��%�@��k�k�U+�7��i�2�\[�('�"�� �N�5��[����x��[�����)��r�+�{�-5�2-����$�#�7|�-��vk�bC
�.���Fb��d#�v1~xoYkM�]
�� �'Z@nd��|p�ʧ��f��>��t�N�5S��4�ɿ(C7w��\�����dɍJ?'�J�|��7�;C@f�9���_ai|����H.�o�"��|4oU�vv� c�HX��<d�6����*��u�w�j�[����*�Z��Ӧ�C��%.+��7��c�\�?0�.���:z���6j�����BD����4�o�(W
���K��Y}3pa���=���65�m�K�X��C;��B �Q�"�:IA� U>�3��x�*f��� ��ɤE�Q��ͫ�\i^�~Z�Y�k�c}��k�J$��B<>!*Gcf�]^��z�I+�3�s!���]��ӧ�O�2�Ld����%��MB0��Ÿ�3_����ǃy����t68y�n����̓4Y��s����.�Q� ޱ<А�}�4W-�c�}K��U����9-�����4�����Q>���jk2�[T�ⶭa�9	-	U���&�k�������~����j��ܴi�%u�X�xo{� �&_���Wҫun�Ck��~ł_�7S�p.;V�%���س�?�1�m��A8�F�5y��