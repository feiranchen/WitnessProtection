��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�;�d�D�ƹ�ŋ+^կmh��V�#0�D��D�d��l"��|��̓�q��k�/_K���Mqt����>M2ӯʨ�O4ڕ�T|�b�rS"Γ�u_n;%HI��)nn��ىt����!����z�5��ak���\���H�be��
�!@	�0���Pf����[%yJJ<�ݞ�h1R�;,��=�5���������up�v0a������)�G���[r�x#��HI���O,ي���f�~|'>�h��w�����WS2��͙ϳ�:Y�\wQP�\���~�sL���Z��������,�ѹ�d�-z�X{���_e��F���W��s�ߒ�*�U �
Q��Q$2�2�~s~�a��ː}�NjK�b�3��ߋ�ԟ��a�������!U@�����\�ʃ9Jr�� q؆u�X�D�f�o� �<J�I0��~�g�pe��#�ٜ�׏���x��S����B�3&��[/�i�K6�W��\��fP� d�X�����S�n�w��ɗ���G}��� ���o�"�k؟$�o��%�:]"�I�C]h}*{L�[! AeX���L�&n۱�K����fK��B��-.�	��QI�^I^���8�vB������E�MQ�H�Qu�0Z�`�Z`�K���L�"� Db[ŵf�&���md��F���eg< ı6��C�H,���������2J���V�!ײ�2�	t������l1V�>�@�0A�z?Q���$����DS��YR	R�軉<�A>}�gH�-�Ѽ΄� ���^T��	D�)
6"�`�6�zej�`��5O!����$�M�f+���d�s��Z3��Q8�2��`��D��K���9��J�ɼ�lV���Q��\��Kz&�2��ȅ寡5R gɆ)E!d�#�r�Jv�v�v�tEz��և@��:i(w��*sV$3�t��2��NyC*�n`�FM�%�WLU>M���'���D�&�e@F�%j�ĦN�j����/)9�E6��'hk��6В�\�Jb��t�䡎b�^ą�q�ɘd]a�q���˽ۄ���i�_��ܴa"�9j�
䊲�2�e	&D2]��C��=����(؏�Ň-���]�T� bSk��^#��rv�J�AOVn;�J(��(��@�SJa�ǌ�%��m�K�3�Z3��n�X�zL\2�f�N��G�8�{����@�ͩr��"��>���=cS#k�|:���áo�s�&���2�1��E���(ˣ�x���ȝ���Ӵ�'�	�r�Λ忈��s���D
+:q#�!��l����Y��P��jg��ic�S�T��S�t=����tA4 ~:���)4��h��c��\�9W)����1�-_Ś^�A}f^� ���d�9��ӃD<��`�|��߰3	f�%l@��+wf�e�(��"N4sn�I�o�Qk =�. �z��%�H���≯��ɨ���bf��rB��N-)����6�zQ�:b�Kz��2c�Ү�����_��$1|	G��Ȥ����V�.Ҕ	��I#K!�s����}�P-���0�L������b?��}5����^�=��<��rOW6��*����;Z1%t���!h9D�a�}�!��%t�{:4	o���3]7j���]=ZzK����Tu� \B�.3@B�S�����.B �Q���0a�=��A_;g1"���ٍ�s u�T>�4C��[�7\����'�ھ^�&j��8�o�V%������PE��H�c��S]���HLVGj�?���d������-��~��S�	@�4���m2v�s<Y�ͮ��bkO�� �I�q��X�j6�����޴8�DF^�2S���G[�a�^�5�!�x)��m�Bﴮ������� =��d�#���*%�3i�!5J��gz�{@���$��1��-l�����լv����
z�@޼�K �	.����Y�xƇ�am'��G	�e����$}�+��^��k!�\�F���iWhĦd�D��U1���6��~V=�z.���0����uH���T8*`���(U2�%�6��S�`V���ڍf�h��2�������]\� aQ(f�^wj��>�N��e����[.z�.SZOJ�Q��>��,�+dBg*��Z�V� x��il$�܇��N��%�K�K����KP2���6l�@J�=,��֡H��k�si�W�K~4�<hIlКkvy�?8W]��������(3����W��Z���dC�$��֏*Y���ᜊE0�n}�%��ؤX����KY�vRʣ�ǔ�L��O��|�^)mM�%�a="6ƌt�*�P���	U/¹�P��MdR�Ln?4��܍_,�<�p�w����,��)�M| [�%�F�q�i���ӧL�?�g���y���Qi�H���tݺ>�y3ͫ�|K��F���O���
aPPrd�Q0��l$��+��w�Ճ�T�o����Y��@G�Ɖ��$]ڣQ��t�0�p��&����%X�c�4*�x�]*{6��E�J��R݌�"�c��e�94�ێ`���GU�,�06J����*z�����¯g`�r��&8E���y!3\ܞ��]3����U���f�rx�F,C�O���3T���1�ż�C�=��r�̅�6g�c�!9n�i]�^��Qժ�s���UMJE�/"�[��A�}t`*Զf�Է�����
�[�IB�ݏC�l����]�?u��,#5d� ��#h��\�U5����j_T1�����e(�L�$������P��BE����;غJ��3B*@&����F��]�X�h��a�Po�������M��2�h�k)Z���V�x%w��p
}syI�Ĝέ��:��i�tT��D���L6S�)�<k%�;P�����3����V)N~Xc�����iBަ�����A����?_��y��>�<�gB����D�����|�o�o�xL���~Fƅ��3�$E���=P(c� Yw~?Q�׎ޕ�dzk�D=��a#��י/0��^����R��&"�鰁%{ށu$,-+�oË}��.8��{�2,�"T���PW�C��Cx�V�:+�� ԋ���5��-��?k�{h���8�#8�A9,��M�J�v&����X�'Q����0!�W���[�sC�6s�)�nƈm�9���t�p��P����_u,j^}u��~�M�(�����^�7���^����.-�T^aK��h��%[cH�7E$�p�Z�N��G[��<DV��H�Ut�����'����(mY��aN��Fe:����j<G�@�$p�!���XJ,�F)7�fA����l��{��Z3�ef��1�ۖrCu����?`~X����B%������5�	^����	��E���P����X\�K��V��0/#]��Th���e� z���0yf�byj����Ż�y��P]��s 0��-��=-�ђ6�_�(� �6ٟ�/��(+�㧛_/�#����\��{L�������K\�@�.BM�0䩵��|��1�\�"��Aç�,��X�����w���Fm�䤱���;��u���.��Dы��	j��5�m5z�'�W -��T
���v�=/I��e����)�L0�ͷA�>o��p��ckG:N��i�T~�#�%F��?�n�~���>S@3j�"��,�z�G��[
������d���e�d����� j�-l�怖�a�j#}fF�]*W�ql������DS�Ų��[!�����t�.�*���ˍ�6t�9�6,=:�񘶢Ff��NΜ�Q�9�Cܥ�Qu9h��+���;SHօM�����x5鈱�C�K穙G4�>�]Z0=�����<0s@�/��-|���i�/y��v�RM-�F���Vŧ�1��}
f�����N�Q�g�j�(/�<��P-'mo�e���Ӯ�1��kf�K��8�d7)I�p�o_��@����S#֒���˨��	�ES����	Y�.�������N�-H3b��>u�$�RS�wU�N��j
xk���6A������.���W��D���)g���w�#ʬK As�"�VνzK3ڦS���:2�5g�+��f�$ʼ�Ԇ 'R=��r�-	Dcw3l#*/���OR�0Bxl�~���/��Pt6����I+z�y��w���o \��Jb1ybx%�8�V?�dJ��wfM�"��v@�Ԥ�6r��9�rj)�$	���GhZ��V��ӈ=��8��c�u�/i���K�ĹG�p݆��kB��S��o�Y]&���b^�� jVB?Ae��A�M3(榉��*�t��VdLbh�x��2�B_<�0�n����Qm,?�I�,m�ׇ�+t;|��."����s����h����
�S�*LEkN��r�=���!!lߔ�I*kB>qF}���I;���L0K���FvL����F2�����|?�Uf�$d�wX�{c�\-�O�n����Y�uo;�vivV��`��}��/7J���K�E��aK\
Ƅ$�d�m��&^"0)��ʽ�|˦x���y#H�TI���	�KH/gP���H��]{$+�~���4� $����m�}a{�=�t�?�-���ϑ�逌�-_4��AWYR�
 �\�~zK�w
�L/7(�7��9/��$}�?�Y�+��^Q���	h��m������+n���(OՐq@%����Le�t�n����@!YV Z�^¾F����9�������`�/cP�I��6�"@��R�>�(_<5P�����:�^�ـ�3�MId ��|Iۯ%Ư	Ԕ~��c��T���� �.��'�l�b�oW���a6?x�0"����o)�w�	����9F�4��.����F��5�/��i��#nGߧ��W<X��ڠ[)c�6�x�C�� �qN�I��gmޫ��W:k��r/T׀��6��Ѓ���������M��R������C���4�0����aH��"�t�'ѫܔ�y��a�/n��1���p��x���1�Wr:����v�(�8�u2�G]��懌�y:�AA�73־h�L�/6�9�Fm�*����ݜ�:���=!H5��浵ֻ���2.����(��[�=)��9ȁ۷�%��]�i;���ƫ���:$�-�t(i̙���%��e˦�|�m3ź9L�"�!r�/dk���}�'�I��%�hǽ���2UHy��E�&qf�O?��0��L%�dk
����[ST���͠�>0�{t1j]���>2�R[ڈ�1ʗ����=8�%�eO�����6|��;F���]U�ܪJ�ȭ��K_���2�����֪yEx�t�ա�� ��8�O���jLG	�[u�1u��գ��eR�5xŜ΄Vc-L�$(i]T� ҩW1j@c�	*ܑ�`��v�!�[����<�Kc��Z8a"�S�x����4�B��`�;�N����^i��w�`�\�k�`���	�j5��?^[נ���%�z�T���~~�;�,�8j�Z�ECa̼bL�����@�uXEl$� �{H�}ʸ�i�k�a��V��ӓu^�*�rsU?0*�y
x���	ț��x��ƫ�r�1#����yǂ��e�[n�$i|���$:���5vL�0_e	^|�C���]�+`žu��f4��u2�ړŘL$\��=������C�a��7W?�CQ�XD��ݟP�̞��{��C�ɉ>1���Dn8�L>w��)�$� V��o'���A3|�y;Ed�&VE�Cs	�6eK�K��2��Q�Q�ypDڊ�9jb�@���	(���v:���lg{
CX@���Oc��>"|�s�J�A�>���٬���D�����/�Yڑ�������&�!�G��"e��E�L8
6�����H�X��oh�z�7'����`�Z���1�|�y�/l>�"������M��؉��w:�o �G�I�r{D�9[�ՠ�a a�inwf���N���`�d��P7y��&��l9��`$�>U(��`��N���n��o���Sl�-��Ê��Q���${��s�_��t)��v`X"��6�:D��7�q�<��\��u�6��>�����w�0��Q��)����[��7�±+I�
��� . f�)��&@�}������.Yp1��B* t��8�|�)Bz���C�Oi_�,����M��ۊ��	#y'a� J�P��Yɐ�?���z�oH�DM�h�6�6�)���q�����g��n�L,f(+�%�g��2�
����c'9��ڦi�����CvG�>bX�ɚ�Q筕�.�9P��:l��5=~1�m����2c���%�|,b�7��o��m�f����[�´�WB�Y2�J�?�O�@v0ס�R�N��9u:����՛�#��Q��G���+��4ؕ��B��z�N��0vCS���$(n[�G�
��d<���w�tL"�h�~L�x��R���� z��<m�
����`�ۉ��NR�D��8�ߊd��t{���:)4�{ԷK`��#up��L��ᑙ��!c�� �t�x����N��ձ_-`i��.f��XǼn�$����	s؅B��r��,]��w�n��N��]JN�@b���@:�����Q����\n���XT�T�h�JZ�TD.Z����Z徰Ȃ3���V~9/a/YK\�����1�u'3���d	��^߆�3뺌ցom�d�O�<�\�!OS���f�����Ԡ��ᨓ�қo�Pr�<6p>T+�����
����_���n!6�@�3�"��a�dh�U"�L�T��)u��cO��l�6���e��
���1tX��	.5���\N�ټP�Z�h�>1c� ���4�ƃ�`T��������a��\	Z�~�^��9b̜`��Y�J����@��(_�e,����.8����[��g��^DI��F(���s5��	�n2=��i~b�݆�*�/cu<ݷ��J) VPyG���wIfk���i,���
#�?aԐyK�k%O,�=D��"r=?��XHf�Ck�8A�l��]�Lx��ޡQF�禤}��v@T�+�ǣ���|�LkM���κ�>Y����\�@�g>��'�/	bd�#��������wK�ߔ¡#ū�˰��!��0�,�':�D����p��K)iM;/�є5�2kT+?k��u*" �\�?H��;Pqg�3.���L��Ƞ��h���(��zn
���,�{H.�Dי�i5
L����=�*��.��#�_�w�t��9A̸r/�n ��	��xZ=g.���>FK�ST���$��
����6V�"o��h����d?�1N�C����:N�x2q��D�m�Z����g�N�KM���G�iU��&yv�����:./,��ȧKk@�� "�:o�Ь����G!��'���/@������:�~�Q�ܤ����Z}�ΰd��)��KL�s��;���fs��q�[���Y4�Dn3aAP�)U��7ղ>9&Qj��x��*��7� e׌��
�ń� �c�����n\����5ż'�]�w4�6�ႅK���o"�c/|'h�Y�����C��8A�(�Ec��d��xV�"	�m�	7��1�����GQ��9?�:�/>$�mؕ�%H'E���Ǎ4
��	{�2�(oa��kD�dh>n��`�>��j�7��Wk��[�HS@ {*	[��7��1E u�9��^GRW`��kqd+�}���9�����'�ұ;=��n�"8L=�?�4?:����fa�P�u���q����7hw���{��w�_���9��o��t�1��{�`�C^��*�����Ä�lUn�/̠ !X�υe֑���tx䒑m�RG���9}����ͬ��p�Q��"	=�*����Q��r���d��~��&i��ýu���cD��y�~Tv��¯��g�o����'��!&Ք�a�Y7m�m�ؐ_��QJ7s@���+O��ƹ]YB��m?7�*{���Z)�a��cܮ�#b#݅��ŠݯIyw{%~��z<g�w����{��渷p�b�}d�BY�XU[BZ�"��Gd��f�$]7I�+,���}��G�JQj�=�u�`@��{- 2�����C��K���ܠlm����SEd���z�Ed�m)��3I��*��DNaH"c����IN�����Ph��0�4N�̯����'ۏ(���hޤi�S�)2t�(�>�ݩ���Π�����2R�����:���+�=�W���͟�B.&�`Ӊ9e�R�%2|�y )A��ș��S1İ�q\���0�Z�]hbR��B��Kn��m�� ?n����(��}QK�6��j�g�8�S�W��|�>T�W��AA�A�Й���6G�5.�x��T�C4	Rnf+�_v�p��Ɠ��>ɰδ!I�Z�J�}��ԇl�����;�s��4C�#Y�"�{\HT����b=+��%������Z���-P~EA̡��%�*{��~()п���.y�8X��i,�k/L(�cy�P��J�3z
x��m�=��lXl�Z�ǖ�a(1���!�������<�+M��-a�2R|���M������/H���(����9|��Գ<t8�	Cr.����`|ƾ����e>HC�P�wV�^:�3����ʦ֯�X�ۘ�a�P�� ���$`��YcǆgQ<��x��G���OW��k|�2oL@���n�8v�_ �Wʵ�h7!��T�a�rcM�G*�	÷�׈ H�3 ����h�J�ye �/HW�4ŏ�nq��k4J�_��hY��3����.ڃާ7�9Vz�N��x�a=��,��"𳛳\ε)<�i���x/��������M�NY��0J�ѓ��Q�,�+���Ѯ	_����PI�N$0�'4'�uLf��p���-p�h�^ۡL��$�?��Y�#���� U�#8�'26랑��VDر����>����6�C�	�V��LW�I�NG�Ϳ-�x��eΌ�4�<e�~���m�$^ X�	��J��R�p)}�j0�T�_@r�L���
��W{kF����K	`��*��;��E�M[��u}�&�ZT��
�����Gt&�z�Iy�qiF@bɠ��zO�Ɯ��|�VE�)	]Iu �'d���]��7�x���#ߓ��?�@[�s�6�S�`�w�s,��*���n�J
*n���< ��3���X�$D`FV�䠾�UG�#ؒHD1Mة�ya��ň�,�H���S�j��qSs�@�!���>p��z�������t�)�}j*�Bu7���F��9�6��1x�Ԏ��0���� Y���C�05�]�)EN%�Yn-7��~���F�%�`��0��x'������~�u��]"o퀉)oH#Kz|H��M��"���:��R�W�~��V�Y)|��Ig�N�?��ׯ��Qz��*ǘ�I
}�z�t	���e��W��%l�+���h�͚�)Z�����f_�[̊S��SRK]�H�5^.Z)�T<��g�2ࡼPxT#��<�@Q:+��l�'�<!p��KU�	�з{~�hsU�o�O�pF~g�^le�ul���������,��H�q�@��4��+��6��=�F�z�r�I��hݳ�B�%�'̄�쌗�1Xh=�c#��2��W�&d�H�p�zdtC�\�1+��_���%Pll Ԟ��%����E��!nv1���
����0� �N@X�|�G�R�,�=r�2tU�uǆ��U�?h��k���"�����w�7�k3*��B��zK�(R����P5�4xݗ���u���2qv)�kZ+��CW�UL�T�[� �Gl�ǭ}�{O	N�<ȶ�'	�I��H�p!������Sw7��7���g5a������l�_Q��
�^!���n/�ֱ�����ڨ�X%F&[���9�h]��]�d�_~�B�7�Xҕ�K`Cu�O�?��W[t���_�yVW���k��<�E���^c�Ʒ�/M^�i�BK�kΉ�.�N��>��G�H�$�_��C?V�iU?���USXut5����-�ñV�]϶�<�=���w6��m��9��[���|��'��d�@"KU1��bM*�'i{�Z�����ܺ4�7��=��r�����o���?©���By����Y6Ue��]w�y�	��i|�׷GJ8����g(����ߨ��[��m��<��D���%\��������)�@~�᡿�._�`n�ݝB�X�p$�P��7�,���q{R�k�4�]?�p�|�f�S��g�v��X<�&�>���`�+s��9t����}���AK*n ���F�\��g� c�� "2�.�m�N0Fy���-	&��5'\/ު0��7�̪�o= 	���\&:�r���n� *��.��Gl���:X�?�uAI?M�n%�y�gll�
���?<Ub�@�|��g2b�QW�CP>�﷞��&.�����j���#��WL�5�B�	i�3�w�]	���/DԦtBL�){Z��� s����/+��é��n�a��X*�/j~�(2��&%Xpoyc�y�֋1�=�!��~����^�C6/�&<�zŒ���ĴW�[�E�X���/��IG&L%B��=8�pD~d�����)\�n�u��Y׊+���{��H[_FT�ʅ�ƁQ�~�-�ۛm+����*��j�E�Ǖ@��ؿ�e~WI���`'�S8g���<�ĭ���B-{ ����+ɮd��4�#?gH�=t���Å#L~k�^ZӲ䵏���9�=��.��ÿF/��Φ@���$uNC|Y����gծ��*�W�_�!խc��s�d��龆b��s�%g<�L�1<�2����՗3�?�(�U�, )�.R0UP%d�Xs��~�F/�4�Q��P}��H4<9���Λ�MG���D�m�8�����fL�!�\��QH�خ�����l��翭���g�x�HJ�F��3"�O��B:]��^8�j5�p�����ꗊ[��xm��c� �gL�W�U����R�`�G06pk��ì|;�`=�v�!�a���Yָ޳�����3�4�BQ��R]ѮK7�W���✟���;��Ҳ@����;��D.')�V��Yg� m'��Vj�YZƆ@
�Ec��N����M���-�$��0�{��5�D�#��'D)a ^A����:��d(�,���UZ���K�����<d�T�|�z��}5���1���4[�rd6��DYA�[�^���+�%ç]7����\��tL�uG�/l�{�_�Xfh�Iē�s���ƽ�Q�a�q���#:��2Ơ��D��Pղ�����n�C�R�;�,.��R�$Dg���AnT�ܬ�-!P��(*��� �Tjķ�6'�/��*�F�h� �Z %����y�`�X�yN�?����)���9H;�H�mz�O���w��~�\����$9Mlf���8��F p�����{S?���?n���3�!�0��3�H-�1�_ɮZ�h��$��X��	>��f�9�W=@���%���7H9?�[�V�Pr�`�3�$�ZΌ���E���i�g\0�B���B���\o�߷���o�V5��q�B{${=�`y1�o,�:�^��b1J�ah"�K�F1�Ѿ"��0p�M ���bj�sf�_짩���s�m�y�6���?}��']T�w�W�I!b
~��G�w�K�ꕑ�I����x<���F�j[��u�.�L}-�X�S����v�:S�������ӅxnJ�P���⒲I�G;��
��K�H����ͪ��%
�|pq�>�G��hF%��������[�܆�C=lH�,�l~���ˢ9F�z3�P��d�(�&/��@vftȠ�Q��R,ϔ} ;�8(n�e��ט��ma�$k�Я5��S��{s�^,��
��H����o�Z䞍��^f]�1��i}��J��"���]br���ALw�)鯧��y�T��,,,��] ��н 4'CF�U)J�����b4ʘq����ttIz���Ӎr̊�l��yz2�I�#Ǒ@Wx�e�������Cp��������J���"��ee]"�-
��)�a�ӧ@���m�Xü:RV�uzN��!�0�7�7��\$M$�UVf��
n�g�c3y3���~���g�QQd:	���f��幑���ʗ�nŢ,�����#�z'\'ԯ@}��`��C���������DA�b&�ј�l5|_�Oh�l��wYq+����q�q�'R�.W0��~�x$�!c���]KW����y��?�)�]~!��Z�Y������x���Wځ�?��D=)���٢�ƙ�(ss��4��E�F��_�@H���?$ĸ�X�ZHuf���pV����V�5y������=f��hj�P+�{.*"W���#f�r�6u*����c���F)����ڵ{$���u���*	UdP�XO��F�B�GQ��:�-�z����}_o��E�2O�'�R�%Ƌ�6��	�Ьf/�`!T0OF��Dc��	��6��/��$r��O��-��+_�i�o��XU��9��@ZN��>�F?�
�vę#��㖝O���ב�ީ���Q�.m,u>zm<S?&�i[ȗ���d�Y/�.���R��Qd�\ &�
��Ԡ�c���p�9��g��u��cY+G��`[76��* �I/Y�HRX+5����<o �u ���&/&�!XF��B��c��Я*$��N�[F