��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�Xn��8���ӱ�̷׊v#�p�<�@-�'���0���GD�`�F;�#x��i�!Δ�_zDf=�T�P��^8��ҍ ?=e���?���aN�� ��c���~�!ܮ�+ʳ ��.�#��b�1|��P��}T��]Df�+��͗��gW���ѕ�c��o����ͭWq�W`��A��w�?�S~ ��ޞI�?F3��h��(" ��1U7ѸH1.��6�Y\M�vU]��dN���j4�R�6;#�qy�u���o��4�~�]�?�+k��ڙ�L� �ͽ���c�8��k�Y[��/%6(2�Ȼ��$[�g���Ļ�'��:��uh��ʌ�jc7�����<Vz�5N>ʉ�:غ�'���R6]q��'>h5�d]���vn�7*^:��YW�HPZ�q:<p�FA���d���#�n�C����4ؕ����zI}>���L���S��*�(Y��=ҭ?����ַ�#Y�=�6=�K��iI�8x6iU]<�T}1����E�rM��|�0�7���Kl5�����L��Ԯ9%,�� SJ�a�6�޾��\��G�C9�K�������K�����:�hl�_?�	E��fZ��3y���O�N��S���/u��hpi��f���U��r":D-D3*݃�6;�%�2N�K��6���ڽ�pv(��z�,���/9����˻o�FknX���o�_�2�>|ҡ:��e���>|���]��?!�u��eظe]W|����́l�WHA��8bK#Q#��9�T�Χ ��bl���پ�0��xf� ޝ��h�v�
��DՏ�{w��;jK�����k�{��~�Ƥb�;D��ՑF�*F���^������#$Ԋ�0�Fҏr7;�� Aj�� #�t�K�����[e��N�}���/;����@��gU�kq�˲D��$���إēND���k╦�bp��8sY���&Ɓ0{'�!�'�E�m(ޑ�T��^��5����^��66���Ji�|̮��C���� |:�BWZ)^VT�b��t�n��%���y�:���+�0��mފ���.YVAv�f�e���c]��yp&p���:�7�q��k���-1~���l�1�����%Doٿ#���YvV'>�����>-�#�sP�"LP4�� m�:m3�c�Ձ͂�$o[�k6w4.6��� ���6B�䗑�Z�޹օ�f����G�p��4���.z�.cЊ����:�;־��M��u��h[��S�c��=[op�2�^c('�=����ȍ��/U-�Q��3����������'�2���-4l�����M��16�+�x�'��T���n��`6��&z����(���+m
u(��㫐��/F�V�w��b
L���+ư����EA�=5��DOlܕM��p4�,G_�3�-�:�0�CQ�&�=yGGue�0Q�9;��D
��xF������*C~W���8��	⚞-4۹R7�X�e��������������(@ψH�%���h�ހe^� ��y�:�3�v�r������Z\5��ɞ�~8�Y�K�%s���vjd8��{���U��vsTn��JmM.ܿ�0��^K����p��\�=��e�*��f$tV���c����
2�W�h�>܄���`g����!@?x��S	�����V���eu�x\�jS-�e���iH �� z��Er$����h���1\���/�����4ur-�����+�Dq���8:�Y��<�eQǣ1���Q��\!IL�ʣ�`��Ċ�E�H�=�&=�K��A�W�� �����C����TȂLg��ܡS�I_H�&�}1�$(���˭D}�{��k�d)�����	Q_#?ب{M��FȻ��D5ۋ���ο��D
���8����lt��(Gm_�Yt]��n-6:"�)�����N�˥G��4#S�+�H칼*c�l�H�0��f�r725a>4�o���W�D���'f�)�Ct@�VѪ?� ���Y�UΥU���d�b�#�v�Ӟ�d<3�d>�b��{���%�	��"K���CjD��- d�o�w���+{S�����#���n�
����>�N�G�Q>�.�K��(<Ev�V�����HAք�1d�|��a�>
2����GĮXʫa��Kr���H��,��}i0	4G����8qV�U?e�̨欨�\S(���V�a�M���h��kTmz3H	c�1�jR7f�+���Pש���s�Z��5�
,�w��i���?� �m���VE��_�WW%���O&N��R���&���Ε�>�Z3^��3�,��ƻ����sB�N�����D��q�)B���nj܃�ö�JC!rq���
� ��^���+����I}
���2�fSnoa1�	)0�S��f��i�K�.��$2�f l��$�d�HO`+��bOH��*���96�;��ĉ��ů
n[����I={�$O�6��rQ	��� :0Q���:S�HH�ۅǕ���F��٭�.�������%o!���	w�e{�K��t��0�-�VY�tl��86g�WeY��������k�zm�D!���@e�	�]
��p+��o]o`-x�~B���!3�{�Pk������I�'�3L�s�T��zٟ�)WGZx"G��5�� QR�N0�Vf�v�����ة�_]й̚������c4�ǌZ&�-ݜ7wgoA��e�1?�&����T�Z٪�Wx|	J��z��k�?q�E����4����0������g�,8�)�8Ѩ�	�T�����}O�M^�ˉ�=b[<�?��O�N�ݢ*ϭkM��d� `��g����m�6�7Z�E�!��}��E&�����0�ȕ`MK �.���ٜd�]��\��pZn#kΝ���|i��Խe��U�^1��jX%���G�\bB˾�U��kɜ�+ɹ���,�}8��rb<L�L���/`�3!c�c�� W�T�<#��Ɨ����&+lt����tS�2��ò��X ���E}AL����'���V���w��a��c��6�K>�ax<d��Gig��g"Bd9�&���iʉ�#(�3�,��1x%�m�Y-�ш�P���Nh�p��ն[e5s�.n�4;p�7�"���l=��٦�`��^r��-�(���޵���ώqBF�g#F\�{&�gJ��H^l�dA�̏���p�ʨ���d��B�C�M-�j\E:P�&�q�<� @�.eh�/��B�&�� hb��qt3����s�jTR�1��`���50C8̔g�����T�]�"*��k��.5�����u��A�J[ꚱ幬	k�si�+��ʐ�.h�/N��]��W>���(S� ]I��q|q�>k6�QC��4�eD5#�n䪃%���qj�R�m/���)��o�����-��J���e*5<c���1�N|D�~��B[��t��J2�/���E�M6)�x��V���|���Ѳ������bݢ�}/�o�g�h3��Ca�P/�3$�����X=��Et��U�n_|�Z����'\�)e�B��
	�3�I�ԓDb��������z����72�7"&�_�,�C�tܭ��gk�E����9)K\�(\�ձq��\��t	����U���C�ɵY;�4aQ�����J��������,��[�P�m+'����3�w$><��G͐�T\0}PЇ̪�D�k�>/��}L�D��E'�3�����	���x�o��Ń�l;���V2�W�=���z�̙��o��>-.���p,H=�yoW��VZ�=4 _�|�q"J�W�i�8���h�*:L���G	�X��e���':���<�R}��d�7O��|5�_$+�-���gA)��v�/)лp؝��P�He�r�
A&dw���0�'��Gy�x�>�}?�����Z��	�o}�}�|���s��Zx�����F�R�-�!&�� #��;�����t�T���1pLy3y�&۶c���]n'���/R$ht��1�v]����RG�~���{4��K�S���6�*����Ȫ�͈J͖:#���[�|� ���o0��K!w�4$�!	TӢ���sҍDr�D�r�	,İw.���7\}�X�ёJ��\mP=;��	)P̭��8Z��L<���P���e���^ޅ�'���Q��P�^������O�?'�vIk꡴�m'�-��Y7�kS�e��u�̀��7jW�⥱Kem2s$A'Ӱi^|^��h#�%�yҞ=�Q!�A��Jd/�t�盜�����(�j�<ʯ�Z����kgV3�:�Z���,��Q��*:V��>"�b�S��Cb�%L��aj5<��36�cM�HK�+_�l��e��g������0�f�Р�l����#�V�R�P�ye	ď��l+��"`��|���KƉ�<�H�>�a�E#�e��۠��0�1����^-����F!ي%̛�)Z�g��"�.�n��V���ȎJ~���H��c%^��ۚ,�9O
�c�~9�N�6�nI�9�����#�?Ng�&�J��W,�w�q	IHSU�$'�B��Dč,I���M����>��"��Lל�_J}�0ۘ�7)T/|:��W� A�;��38���T�����X�v��d쫤���^DɎӁ�V���K���x�����"I���^Sօ���4V~����>�E}�_"����\�ȋ��s*�ZE'�� �>��n�dY����ʗ� m�C4�)�W�'f��=�՚�Bۿ��y�CX��߿>�� �xԳբJ��|�o�C����J���ת=jf�s+�[����S������8��Z�y���$P�A���༘po�~��9���0e���ojXTT��NVf��+π[{Z��J=#�FiyzXJg��b��Ņ���~F�Ɇ��X˛�	�4��&A�&&X�]Nl�fv��j�.����c��6�2ޝ���Ǿ�	�S@�g	Y�27����r���� **-�
�#T�F�Ӳ��2ؖ��QU?��F:b$ȷ3�{�p����%�uy�x~� �V]������^c�2�ϲS�ꊱ���W�
E
+��<&B�Hi$�b͹4m�����8�X�~ћ
�eF��$��ؔ�P��ĸj�M����Y�y�OE�]zIo'϶������g��㔏FP䍵=�����Po��!�?;h�A2}kb�k�'�"��|̒}���f��I/ܡ� �������� y���������4�" �+����9�G�[���E��֥�zD{���h&"(��~��T�bm�aL��K��;�r�Ĵr�9���*U�����)_��K�I�qI�&�S��ׯUj�,�ǔ3�=�v	,[\�\�ݘh]��e����c�D�(I]�9�� �?�Oz�YF�?�RQ|򦚟�X(��0�-ȁz�x���>�ٽk싣��gw\�n���%?��|B��+�Kp�.m�?����6|��+f+,�1�4�񐓠(9�"ɂ�����:0t��u����1��-QY�qو+w�3w�mU�y��f/A�W��D��bZ�������'��F;��o	��
c-r��g����r�z��l���lZ�n�!U����ŕJ \RJ6.�0��u��7T����8�⼓�d�Y<��xwy���/��m���� ʙ8{�C�W�V���~�����j��>cI�#[~�\��x���/����N�w�Pyf��E�'����uο�!m�µ�˼�a�"6����9y�C@4@(�(�Kd��[���]xS���	��#T����?ٴC���[���6%"�'A��F�)�O.����g��uz*g�����=$��z|������9
�Ra�)Y�q���j�L��VG�밲q@w��[{|�l9�wߜLDwEK�ۇ�7޽�g���|!���(�p}��H��a���e����/�:��i*� `�U���
��m��y��|�9Ҕ�������#�G�3�腐5ʊ���M5��[]�_�w�?���_#��5tf���$,�{i6�o�	��=��0��j3�rF���P�[8��%���ς��`�m�ܽ^�\�5��'Č�5.i�U��y��:xZNgn�����%����jQ�E�d(�~Nj���)�
�G5_�N����{K��~S����D�|A�[u.������}����|������*����[����F��oO���cZ�~au"	��U>��B�]J�Df���	ޫ���)�w[ÕF���,lr<���������e5�FV�"6R�i�	y���,g�����=�o"C��s���'�yM��j��A\؉���2��5�!�(o�!�?K�E��c��t%�����ߘ�\����e<(��Zvp3���}����`��A�d���m�sk(��y��Ү�\(ͧO�w��Y�G;n�*{Z'���(�G��M�<:'��P�r��)������Q[鞷��(VV��}�5�#GΗh�cm*�E��z��.��c�)wL�$*$��k��:�'͚F�*��2�8�G4��F����p,s����,�����[V��K�M��a�\�g�zO��i�L���r����Ǒ''
�C��smc��X���Ed�Q;�iJR�[�n�O��^;�����ao[�1��gyJښ1eZ�ָ� Z�����vɒ�6\e� �]R���U|�]�ŝ>u	�-��/�Lh�ab)%�l�^<�Ҽ$�IzR	����Ԕ��aB�QC���&>
nLf���V�w\���Ϭ�uҐ�I�}�Z����?5��|N�y�
~Jm��B�:����s�j���^�!H!�2i~����!�$>l4��"|6��b+ȇ~�5�T��"���WKh&����,����;
��
�P�R*ޫ�� ��^r�i�o8�i���ؓ8[
���%LŢ��a#��v[��?�[+������B'�:��|&�! ���d�K�2a��|5�N'T�?uT+@*37�@��N�˒����	#��t?�+w��S$Xb9�J ����E�D=v�l1� ��m�{�=/U��g�%��>�f�Ô6X�(��Q���L��'�B�c��)¹
=�9gç����;�8uꃖ}U_��uT�Q�2��eK�Bs�'��G�6���XI�������#j_� ��sQ��'����<�j^���h��O���CVL�$�)t���K�iw�ls$���hj�/�ˡ���c�,B�Oh����#M���8��>�e��!���b_�B`��.Laz	W�ι�e�w�,�a�C
l�;��4������N��s���%��i5��v���%�9ѕK�#�  ���u_��pF�5	4���w�*����-Q��c7�N��ba�,����#��.��\u�rb�r9d<��'m���� ���9�*-�-�>tj�����e�q��m��v Ȁ��:o���r�oQ(ъ��>(�R�7�zBE�|P*���"IZ�;�dU���A8�-m���h�"�GoWEP��/������I=�BV\/��[������W�xw�`	ٳ*r�h��U��&��U�i_�c��!�3���܃��s-��1�xf��M��p���jY}Vt���ı�~����6=-F>�ZeZ��8�����z��<�9H8���Q�l�ԽK����h�?����]�7{y����%k�":�	�ID�Ɉ�2:�8� lߌ�ω2'.i�UB�/`ݵ8=/P���J�f/|Y6�������>�r}�Q�} ����Ӷk�����tx�.��Q��Y�S��F�
k;Ԗg��������Ea21^c<t��f�ꆄ�	~�p)�t�&��ށ��E�û=�U��D�9���2z�>)h'&l/k��.+X:�ǫe�,)Κ�������g�d�?�r�۷�d�#۱��*od"P����귚ri��ѱ욘�hY��n��:�aL�]��G��{ۮ.f���� �I���j)�:)O�
0��@�^uz��QZz,�� ��i�sVA�Ƹ^P%��TsYk7�ߩ�z��M�5�f$��-Kj���aJ�;qq��Y�0kz�G+�N���j@���iW$PŐ&t��p��'	b�����<�̷|S�s�����O��-��ц6�yf�h>j�����GV~����p��\��
E � 8I�=qi�\��Oi�v����B�5+�URY���ܚݿ�H�I���Ч�VMTT7��0�[(�>-�ݙ�Q��\5B�ozfAm�"��IHc�����T��MJ>`��=�S�"�9��/�Kj��f6�'�?͐�:��hp'S�]��A��4$4e~�㌣�cJ����hp�,��Ɣӭ8�&�ML1y��8.���
F_@/����:FM����]CX�/��s�'îL���==D�z����\:�"�A�:�3��B�^����}Jt�'�qr�@$5~4L�,�=�̊sE�NS��˒o���L����"�T�0����M{�߈��O/���Z� P^���!����M�e�O�9�IEòr��O��?��ZZC �ۄ��?E����;���M����@N�P�^�\ ����_Cb�y�۲�2w�cv�b�$���*P<����1M�/�咨i�u�ou	$3*�B�� �W5ǰ�
���Vw���j���BAJ�D�Pe���ն��0�2g:h��Bzǵ%~�+��[�+Lj�0�֜�39AHHu�:���諪$++�nR�`�	*�oX�[#���Ǐ�]W󯾇�(���bM�[(A�!��ЩJ���	]g{�B�^E�!�$4��ے�E���;��A�T,��1k主�>�W�w ���h���#�A�d�|,.e>��:�cDZ�v���6V�1M-��G�!��|,m�_���M<xV���Ĺ�OrU8m��c����n8A�f�8<�(��n˻�ƊbA�.�h�/����˫)�c"�}w�B��#닲���3�YL��6�c4����R�e���
�?CI��Ce�%�&5+n�1���S�#�Z�����_=w�'���5�z�S�t�9��l^����&Wf���{g(�B}h���>��CI�x�(���oE<,�)ɚ�Ņf@8��AT�U/�7�cE.�J��z6�'Q8�������Hz!׼��I�>��q��N5'��3�������%�F��"3`�K �)z?\L^`�1��9e��K�.�֟�����&���s�I����%̖½��|��\S�<v�מQ��ş�<G��%R^q�fԩs/ ��`���}�jP�'���&��q͞J�HM�B��/\�u�3� 7>�	܄���a�Nꕈn�ҥa9�P��py�hEo�i�>�?������H�b����n��=&�T��dK��i~Z�TK��F��ron�KE�wbX\��Z/X�ۓ:���p�7I3"�ka�kw?�?R�:��_]泸�]_Q�08�h��q��6�n���IІǠ�J�����7Xn���Z�+��6����"�;�P��T �vTz�/��(7�8-�H�L���t�
<��l�^��m�Ɠ"0�f��u�XV�:���86#c��.U>
?۱#^4䦍��%+����F�7������&cU��z����q��KY�]G�c�#ʠ؊w���`��x�3��i�I�{��d!���|���V���{e�t�T��*�V:��#N���J�~[ɐ��������"O@6�Ÿ�5�l��I��II��!i�I5��_�.�]�ݜpp�sR�Z�xs }����9�yͼ2���l�N;��o+�z5�&nB�Oz���g��[_4�h����_����T�.�8�������^���Ť��{>���6PR�:c�i��Vksz�8��A���h�������p"PT@��I�X�RH-|-���/��>���CϜ����M�j�7��#�r��C-��G�o0����<.��Ue����Q�����o@v3d�2���ŋʦl	lؚC�d/[IK�>���+�,V�V竤��Y����q��IKS�1�R�Y*�=dM%2k���څ�i>�<G�a�]�Q�����1�d�&�l8S���Ԓ�(t���*T>��}��.ޜ��L������ã��U-�(姚�N���*������S�7luIK�0�%Z��/{����+X'��k'�^�^Ob�!��m�-ZYN�K�2�gV!����b1�&bѷAC5�	�\O6W�J����u�s}����"�d	�+��ax}rF�-�k :�����Z�K;�wD��lm����fp��m-ec�x��������T)��j�P�� "C]9���$�S�<��|,ɑy�n�W=���Bc����6$2��c�׽=��2ea%��@�N������7�;/NL����R�&&h�������nޚr��x2

@��p]�j��8D��~���q;�Ƀ\]ħ�obA|��h1��<,�y���U��N� �d�1���<�=#��Gg���V��{�1૳�����M^�P~���̧��@�u=<�Ј*u���C/l�{Hy����V��?�f�2��pD�*z��y�n�B�{��	"Lr�^One#g[h��g˰i�8!�$�����ʋn�TV�⪵X����<�u���G&X-.��g�g 캠j-<��F}:��^g�Z��dTZF&�8�~�����i
9c�u�|hﶂU"�y���{�o��F�B%����!�w�k�ą#��>�7���<�{�R_����՛Jj<�|�����8O~k2H[��q!�s��{��9k��ۮ��/]WY����\o�Īb��m�|�m@�)��	��'m_���K������G&��1�}�qh����_�;c��@^OLm]]��Et��촺���P�< o&��I[��wn?u-��{��Z�#������]B
�=�EV$��(����0p�-.�7������1��@[$��6j�F��z���WIYV�@�)��%����r3����L�yM��w�#f�J���RT�K�[!pAv5a7���km��������3Z��o_��^0�1�=�\B���4�����R��;��Mm<෧-��xp2����k�w�!��-�'3�C}���/K^ZG��B_cV��[�#6���PY8T��iHo�V���!�Tbalf��w�0@2A�Mj��5�� �'ՠ*g+L���{���{�8���(m�������N�@}�[o���d��𕝓}8r��4�M�X.O��c�v�&�%X	W�{�����+�y�����2�x^�x�5�o1V�)�x��M�y�+MA����J-���]�v �q�Jtİ�C�רF
�#���fA���m��,�ȕij'\3�	��<��僯V9.����0��ɞ�V�!#���~׌�Ɂ�{AgAF�|Ʀ���ȩ����V���ګel��R��5�FA]�K �jA��S���y'Tu}!��Ԣ�Z0�@�$Q*5�3������^{�5�E�f���o|`*<?�cz@�J��v ��t��Q����,���3~X�,�z�¶p��7����[;�G��z$Cj��;g�"eJ>Sǒ��e��Uȳ�M0�j�n�ah��T��Y�l9!zK�n�K|J��*�^P���'Ԟ�RXS�P�ݑ^`R�m�&ve�n4[��d]A�xk��Vh����=��4~������L�"l U�s�>��1�iI�������o�e���U(�B����@�����.�D���V��9�&R�lS�JP �����G�6�k �W�Yj�@c!0{�#]4*|49�n�2
�nà5B�"�%�\�W�}R%ttZ酾����W��V&�� ��[��5-��Z�Ң��嗌�'�k�j��/�{�Z��v)��:�ehL�4Z,�� ���(�*oe��ǃ�X��h��mr�V�Hp��SV�o��$$H#KK�����W<Fj$~�{k��S�S��Z��D�)3/Yh��i�K@��A���/v��JtNG����>P�m�@���ۈՓ޶ �^g������b�D	>OI�����"V[��٭���ڃs��Z�PC���<��X�e֝�_Я�v����o 96^ff�x��UI��`��+_|�7��h��)�t4SaC�C��RO>����_KWn&��������֡�-H�Ny��Ɂ���sy���Ax1W������0^~J�mB<�z3�]����j� O���z�eo�����Rd����þ��"��>���/�uv�w��L�%��9]Ka����������1�T>�_��SZj��#lyJ� ]Q�0���E_:�+�-���{���J�Ѭ{)��rϽ�}���x��3�gÃ����4�1�C���o��0��F�2�n��9?kk.��������j���*��u��	���K���=����C���;KH$V��OctEdNb��^O��t�����=�(��_�-����n��]-D��%d�w���Rd��$f�6�2C����*g�A�C�e���������B�3����	��yF-9��u����U�4uN9��d���z�NYS��W	Z�V��dj&�Tdl���((G�Uu��?Ta�b����{��C0/5�4�C��݉>E��r���]8#����B#Pk�r�|�Z��.���6�Zss�
���3q��.�V�G�~����X�gNV�Ǩ.7Ȩ�-^��9q�� Ť3�G�1�wckmW��؛r)�?_ig�st�n�ZdH�<
v�h�%D�
㕼��L�S�,��!o1���iM���@��P���+��Z�lJ V]'75������7���`��.=1�Gx��0��Z���%�J
̯�2_�no��&zŖf��H��F�KԔ��Nq��A�w�Y���;	�I𢆴īio_3��0�
;�Ȼu�C&�־&�V0�$q�T+��qѮ[e�`nw���[�L#��)! B�
r�h�q��1Լ�����"r�(��=U �D�^w�R�X���W��߉t^������O�������4�5��qѬ焏i0"�
~mb���v��h����[��U�j%u��b�}";�5��\�K����;���R�0���գ�W���3���K��9�U�@�5�E+��8ϩ93df���k"������7��,������gl;�8�Pa}J68�{�{�X	V,���[����VvVa���S��Z��u�
�'=rq:w}bi:��E����oNї���r ��O40�����������V���Ęi�<潁��Ϙ�g��S*�3zLcV�t�7׼�vD�W_�_��á8�JZ3�r�L�l�������	k&,�%��ܭΖBS�.�Bv8� c\v}��&�Kw�������Xo,�_R�nR9^��L���r�Fe$±��L�7-Ɔ���nm��B�ގ������)�MuU���{�oI�`�_xw)���|�V.s��e���V� +�6�K���p�7w�D�(1f�ss���tZis�(Vy�)��(~N@j����\5��Nf��Y������,gB{�k�p�%���&OK�I���p���V�H�8��i �Ў�������[)�=�:;�T��Xc��	��P�������$�K�������a ):CX��0m��F�#�� t�,o�=T.�(�Y�Pu�e���L���5���q,�����7���-�$��#�Q"�E� ��ԕv+��jF��b9|9�{	���V�t#�OK�<�%�&�2�[o"uTh���û�#e�m|MN��������\���<��V������o�"u�}���^l_��0��Y8.�4�A[1�;�&�������E<�#��:[�}эY�E��J;$����.�,6���)��'�� "�ڀ�Col�3�7J{��q���xP���#��/}�e�3m�p�e��jE=T�tÞqj��]�	��}�1�b��~���Em{zqS�G!ȳW5�"�D���u�)��5����4�m^�F����`i��T3%~���>%Rc�3��L|����d��Q�K��F�(�z��F�».6�!�}a�rQ?�xM*#���h���?�`?��1�i�K7��_�;O��/�(|�9g+���rb��gt���&=�w��O��l�-�Do1�wf�*<	�ah���}S�Z��!$˿�����h�!�T��C�]����\��6���d6$܈iyR��u<�x�N�T���[�����gI����E�B�^YA��wlw�����b2G4�3��v��̕x���F���8ƫ߬��_t#��X�PJ&��Ϩ
ߎ�� Hb���N�7K�n~G�VV۱	�Rx4����ݡ��9(-�O��coW#.�b�� b� ��f^Pk�~��S��AGS,���1�\�(��ܡ�H�$�~2�~��e���W\��<�ƌ���z�l����rh�
��tg�/ۉ�go�[��>jh5\Zě�m�>Q�9.{N���E_Pić�����:��_�	���c����f����w�Ҽ����\Y�l�{D1m����~'���'���S���0-��3m�O��1=��4�0Z�"$�Y���aw6<<�)�4v�)
�%�x�#h��Q�g�W�����:T��`V*l�OE����/t��^-�><����}4]XD%�X���>�Vj5�r��k]���,�߭�@�PAU�⪹��kG�-�2����Lv���KSZ��w�Zo%h� �>��K�L�9ÚC� yo�z���u+
����Km!�A�r�(/��< ����0_��.�\�f޲�G���IN���v��}�&2�W��{�1�q��> ^:	(��Tu�C�<��s�q2�*.u0(��pZ��&~�{I�+E�mcf5Ο��WFwlc�X̎#�H�<�������� {|���}Ջw�����?�s�n���3��`���#�gK�(��KY��Ǎ]�ҁ�֩1�ه�'����f���(t]��E��Bs��]t�wz	-�����FM�j������8���=`�@�U���4��	^ʦ�tɣf��I2��U�蹪Ⱥ��&��v�6�B��s���S�����S�:fq�ћ|�8;lG S�C-�r���U^�R�GX���r;�/Ɏ���Э�p��d#�jo7���M�����u<B8��|0�6�Xɼ��ș3��q�yr%�vr�Kz�׊� �Aa�z{}�Bݩcx>���p�߷�E�lJ��|~����7H���3�~�!�K]���ЎE뚧�dc}�����Vc�� |2�����������8��Ş���j�Nt����P�6�qċi�j ��r5��Ő׵@��1��E�h*f3o2��� �Մ7%]�R$:���MG_����X���?CM7jSlUV��������#�����~��=���gKi�A��Ҭ�?X��Ao&�wI��Y�$ɾj�y/���Ϛ��uݿ�H�ܨ{�/Ɔ82�$-��Jk�)���w�#ö��Rn׷-����iN���H�3�s#��x�|u�q�I�U.8������}S���` ����Zv"N@ڤ��
�hՕ����� q�8��F��{X$��qqdґ���|��b�?7�� �BX�C��I0s�w
�1��ڀ���uNq����\u��ÌϹ&����ҋQb�[�
��?W�_�}�up/�vL�V�c�NW���/cP�ϩ����\R�i�2g���k�#'��V>��G����)C܇�Ӛ�"�����I>�(���4��)J�c��)b�i�Rب}+(+)O�¦R>m�i�Z߱��u��ʋ[����;�QCBe��Cs�t�EЏ�E��۰�K�\|L�څ�Nr>l�Hɮ�	M�^�0fr�P�yR�ȲH#�؈�°�돜LG�W*�U\.~Ԥ��}C:�Cc���Z���~8XL���C9����,�@0��
x�C3�[��X�bP���T�M5^��a��B,�sA��A˂���h�M^���(���FF���77���
*P�Mble�Z����	���TU
e� �wZ]h*63K�0d\T�:oq�fY�n�hdD?��pJT�7� PRA1���`���/��V'5Խ�
�|&�
%�oM(�}��ש��)�>z�r�m��e�"'É�l� ts�2���%2 ��&��H�ti,�s�%�/j-�m#[��!��GeP���B�>��W���v/��Nɑ��>sTi�I�Ѯ�@H���K����S�>n���f��v2�C�nR%Ҏ����B7f`�K�ZF�36����.�丨lp+�x�%���4^�����x~�,�ڱ�5k_��.GF��;��6�w���P�	$�1Y��.���¥���b�<%��6n��������8�<TY�=_���
 GӨ���xLnx���Sd":�}�X�$ِ5��7�1�vt�?�]x�a���Ye����פm?���Y3v��̳�4�ɪ��a�b�8yD�4����Y�}&ˌ*�a����:Gq��\���Rn��)L^��Y�0h�]xjLz>���n{'V� 8wV|=��͐��k�ГF��aSj���R��b�SJn������7���^j����p�h��i)Iٹb�	��ek�p_˝�O�F������}�[�x�t����j���)����XGRz���E�dW�c鈅'�3�z��3/����	�h�r�˂�1G�=/1��G^5��ᱤ��r���m�����m�?d�œv~��������6�aD���{���!��W��-�?|��{i�/~
���8¶�=rNk�\볡�l��C�i��Z��!Q�z���C*b��Uԏ�'vn��Ę|
'��_������:A����ɘQ'���,�Z��v��c=h�e#;,��ɮޤ������ix.�}I��*�=�����诇j�W�g�ϥ�.U����2pE9�����z9��61�>��&f<7ٰ%�>�}�a�}��^
~��N��v��;u!= H�\s���� ��:bϜ��"��RET0(nO�5[�<�YU�ֺ�MBM>?��P-@��~��8�S^�Q%��̣� �0cl���>���0�ּ��Z{�Jl�L��Y-�˙���t�ܢu�r�\c��L��%
������.^gX눱�љ�x��pD�;�E*1p,`�_����f1'�4P�H>eS�$u/7͡Ҿ���A�q6���^6'"c,muÇ�P��+@8���y����9X�#��b�A�Vͤ���ŧ?6e؊��|���ؼ���S>�@B�.�d-�rDsL8�vj@�ꠜ����r���(~���b� �u�/�d\hD���j��{E��ѹȢ� _n�0�h
ejx�^���a��L)L���8Tⶠ�� �z�v%��p�g��PV̛©C�{9�B! ��#!�B0A�5�ь��+ �.͵�P�yzC	.zdp�@.��ө��T �s�en/2�=[��q�#b�A�������f�ʣ:�91g���%�ݜ���^IW4M&���E'�R�v�����z�4ߨ"�N�տ���/ق�'�F�M׫�����7U2qO�� *ԍ#�:��Ţ8c��vٞ�`>U�-��|����H{,���rL������#dO�	�F#��r.09�'3�Ȑ��lk��l����i�wv�k�%Zq5�h.�\	�J.�wς�}�����b��S�9wM�=3mW��s�>�>�G��]X_9$�x	| ���D��/iF���_�>�8jo*E]�@'��gMd��&玾YUͨˋ��(1�e�CّoN��
�l]E�>1�lN��Δ�y|"����o�k�Ȗ��p��p'y�mv��2|D�"�ƃzqXN���.;P<�'E,��{kX�Բ�tֵ�6���c�"����ڃ�M��������s�]���
�M�V
�_/DjU��2��mJ��%��5A��{�w�ʲ��0a��s�=\U� �)�Z��e�V,�G9gMC$]j�d+3��i^}P�{�CIZU���6M��p��ݬ�,%���bŧN>��G���cK�0���6���Vi�e+B:2��I�Vd�l�C� ��:���3���n`[�B8Ĭ5K�ٚq�,�{Y���80 ��@y���=7�G��O��}�ݕ�)lQ����˧������=]�0/1�MWe�����5�6F� Y]t5�Z�!�+0�	�y��>�\l���"�P�s���n��T����}3<�z�N�Yo�*�l�Ԏ����!�	L`�xo�y����Y�r�p o��ڽ�nG�<�Wa��D�#�v8j0�T��RQk�b�
��qd���0:}��u���<��c:5Yi�evՙ��1]Y>����`���R_�ɉ%mw,�(��
��*�E�HDm��&��cIIs�+��L%Zfδ)B<ex#�In<�$������h�0s#='`���Ažr�%
\΂��L *�e���w���[�%?\�S÷d~��oP����Ͻ��|*b��X�r"��p�3U�L&�j6ׇ�cBBV;)�G9a�|�+�N,���)~�](M����]	\�S^ �k�쥿m�&�ϯ&����vvG�1�[Ph�[��#�WEq�K���y��t2�&`�~���;N"��>�4��R������3�Q����|ٌɛ^�ث8��`X���bM�� "K���F<�y�U�1!����.m}��4!es�~�Zp�]�Z�r�ޗW�i�Ɋ1
j�4��J�8�4�����r�9�V4Wcw�����:=��q�4I$텹���S�ƚ?�|�.i�Ցkt��c���ѳ�_ ��.nc9�-�N2U��\��#���i��S�ǋ5�tV91���b��@�`M�G��emU���mUj������v;�i�hx�9Nz�@������U��+�H�����������������Y#�=�J�2���N�	$tV-
U J��lש�=�}���T�ũH_�KJ4?�C-����62^nc��;l�����,XƑdQ1|��^&�j���nTql�>b�9a�0��y�]ro,�Q��a�	��}xxI��N�a�M��4d'��K|���b#�'S�^��΁_>���Pkw��2V�����>Azz�Þ�}Qz��b��*PshG�ι�gL�X�!$�����!��^9�{����a�}ST�I���g���u-�
���lԀ����~'8��*4�o>
��h�G`}���Jl��]���?�Ϛ5h��Yc�Pc���O��LK�O�@8�҅�l8D� �cH9�:���s�[��q��;�2N���NE�$7�mb�G߃*�KΚt%2�r*�z��DvL����0�A\ʵL����~s��$I��I�x00?�7��F�k"~{�w���`��.�A�h8�h�pc?a���X�K�25i֑���(8��	�����F�Z_Ό�:s/��E�NȬ�O����פ��+�'�w�Ȼ�s�*��5�O��%Z��>N�@Ҫ�+K����n6qӟ��b<��R�� �Z����� a�R����{6���#��c	E|��5�3��j��$Y�L�n
�vAb�?�A��1�J�S��و-�!QX���\�#������qp�~�Ɓ=�6�D�o�x%����T���ɂ�6�v7��������,x׎�!d����'�U̂�ɢі�\M�w����h�� `{!ܜȟk�=����'J�.���y/.�'!��:F�c���E�5���|e�c|XXLGN�]Sj]ARX���,���u��4
��l٤p՚[�Lq���^��2�6�&C)9 1��~gR�0�23'S�4��N�G0�ggԑ�)l�ӎ"�lb%mʥ�ט�{.�X��,6����F�Vj�,. ��@��՗������<+Q�׳�S���+����F�yi%+��2&��0�M���k�Q��/y������V��*X	�韎�g�ж���������/N�%2ؙ�z��߳�5��<��El;Q��O��-�;Ik��XS4߬/oh�b��B]��Y�1���7)���k�;���5:�h߶qD:N�?3�q�����!��s	9�Bqu���l�	XWB��.�J.��l ���Ȃ�f,�r���l.t{��p��s°�Ǖ,�\ѥuK<��N��z0�v�q~�v<�qv�n���$��9�í� ��,�r��^^�l ��Y6�ߺE��{��� ��Ʒ���`��Qe�?�⁋�^	�"ꔵcm���J�7
NPq��Hߵ����H'�fB����� �J���C,���5 �\|n��I��݀թdhȂCX�~N��o�0(GH��PwH����,�旌����<TIQ�ы����3�k|\\�,ۤ[!���~~p�F�k��>a��_3s�߀z{n�m�~Z0Wn�X
�T��V��֮:|�o;����Z)B�Hr��<vhEKgٸ7�~�S�-���[,C�zLB7��n�}�9���H�%D��R�fզ�D궽�k�8)Uo� �xɩPAG/�{�#|�#jd���w{�,�8��Uon����"Ɓ�zy�.�\��jz�W��M	�t�����*&=�9��A��ZE&�Nh�ښS����r���V<uh��f��]�#��<��.s�nB�|���5b�����5�_*mF[�lET��2�ݶl�/� >¸�̏�P�3�d�
�&�Z��3@-	pMXqm���b2'��7��B���T��%�H"�X����UTg�p�>���-����d�l3L��.�~�)���W��EN[�K�ѼD
]�C�ݓ����|�Y�g�;�5Y�klR�lC��xD��,I+).i)ϗCu��o��3����[���*:g�w� ���Io�̎r��a��<��#�7.�[�6Udy@恣��A��-�˥+�҈@`[��������d?�x�>K�l��jT���1" ��%�`�p�|��\j�����Nl� 0|%ƃ���(3�9'Y�d���j�`R�Oi�8y�_ELy���S	�̨�����iZ�A	��*0{Ϧz��e�)���;�k�ZR���{��JP? �o�����u�;~��g��-?ٜ>2r�E�=9q )g(�W�N;��	/���t��VW��ڐ�e����kg�O�>I匢{C����W�wJ�T�����|��oa:��6r�&c�5���[t�XBUQ���&�����k%���i  �Aڳm�Ĝ)�=$ߑ���\H�`���C������0ٱ�5@���JEOS�_lrZw?C0���uÓ�x=7W<��F�m �ԬR�<p!4^k��f��z[Mzۤdc�T�*V%}��V�v��Mq�}+����|[p�)b1_��s�'d�%#>��%��&��}��G��
������\c�^�w�B�	�8=	s�sS��b)Kq#^?��pN�`D۵O�������
JZ��M�wLn��r�x�S��-XߺȖ�.�\*�R�I�W��V�`�?N�@o!5�2Sh��,��zAl�: ɸd��r<�o�)o�KH�#�ڿ��3��Y,)�aC�|���g�#L]
�^g�3W\�mjg��_���^���\�A�z
Z뇛{��m��D�^�R[;� P}���ZM�������|�5�����d���KVs�P�V���� �����d�����������t�5�o\V�	�P`��yd��݊X�\�7榯�0l�=��>Q?��)�8�)(>���ܔ�Ŷ���V����"t����h�13Kj4R3��O��Ct�KIdv����MZ3��{�6�3 Q5;� S�K��6/��)�?��ȑ��UfIR|�,��W� ?>t��5�T���i [���d#���s�u���W�7 �� �ӎ�̨�OMk�����{':B�;�������d 3��� 6K�Wj��d}�|;;�b=��8U��s\C��^āMU����Ru��uni�~�;���;a?1R�������)e�So� S3�J��y�Z��%�2d�]N��������Y<��H@� ��3��E�6B�RX�E9���`A
,fA�;T4�R�������RB��y�ϰr��
�s��c���˥x�u"��}�D�'Xu��M��({Gs��� Q�i�:��H�S+�`���(Ԯ��m��\��^ÌS�L=��'��Qm��ۤ���PI	�In#~�!�^"'��P`��c�R�K1�G����?�ҵ�y���5k��@|#X�0~����`xFHR[�Fg�=5���'�܃� ��G���h���U�D'�[w�(4%�
���[��QM��o8����z�`j�u|M��-s۱vG|4�Izz6ϳ(��,
И�zיB��l����h�L5�� ��5D�Q���[����nT�`�ۚ��J��s�Q;�. p�&�p�.����	1�H5��FI�g1ИD�(�0��k�WT����BP""=���l� ����;S��6�6R1�-��\���u�@������q�����)��y����� �铮i����ԧ'����`9 �v�5#R_�ko�!,���%�%�Ș�p�$����
`l[Ҹ`66MNn+D;e	��X�[P&�G�SB½��r�p���2� �3�3TƁF���`kC�2��ĺG��w���O�Us.��8蝣�<��H��D(��Tx�
~� 4r���o�^���l��H��d-�b�S5��qn�D.�?0������������إ_g)4l4��*���,@��f�3o�U;y�0����~Nɂ3��v7�F�W*�٧�U�u������2�6b�;qw0�&0t���ǀ��MK̩�BsW�e���'����k�عm�����fdLkx;��3�㬌`��Q�B�R��/0�`ڍ�������(��_�|]���S�k��
���L�cV>�T��b��DN��N~�Y��q���*U?	a[�ޒ2rW������POx,�W�����)�aCk@�f�d��� )I��.�z��M���;��U��ol9Z��<t^������Y�`�,/�(��Xfrn��F�1�o}}��_�<k�j�V-�y���(�6��!RI�
SY�;S^Eu<'Qk���u�afA��,?46��i�A�n�l��q�=$C{�$[�ɵ���w[�ZW��}�}bt]�ʹn|���J�L���|���B�����R{���"ˠ���0!Y8X��7n[��OH�� 95:sDf�ŝ��:����]�c3�����&w�,�v�a0V����YB��^��GCv�g1t�dsO��?>�$��<�pl�$g��(�"�v���׍��j�k���3TY��2PRʪ���c>n`�s�DEr��}r���� ���f�Yu�C��[���0@�4NS�e���a��Ľ՗K�й?���o��'G��-��L����ȻWݬ�&��4pߵ� ��ɘQ�bC��OO��Pf1��E&�K����1�']�%M��(�a�U�j��{�����2��������F�����$;����iI��1J�!K�����5�V�0�.'x¥�����FNBVKY��A������X���?ǌ(�,�[6A�U�)��:�K���`�*��'��1(K���b���Y�烧mS���{�4�! 5a�4]�m�����«�W���d��{���e~����h�[kU�D�l���)�Aץ�]{�1����S�py��2�6�r5�# *9Y�e)�J��Yce�KY]i�h=�[�!��&��\ Qt�A�Cz��Z�L^�֝�\�טVU��9Z��P�1J�K-��O0��Kq�ʅ;�y���[���V2Ϧ�N��4���4@h.��uzE{�R}ք�
���<!:f�
�#��nf7&}'�3�b�N�Ast������w2;���ey��(���+�N;пM��T][Շ���4A��f熁.b���R�%ǋ�[��p��� ��1D�-"JK�Os��{'�'sNQM�e(�.$�6��ִ`ocxeO�m1�1�d��>�.E�A���bKo���v�'sf��;}���~�xT�'0��⁤��݅}�G��`�&�@j���l&�"��'���X	|��1�����ah��ٓ&$S-�N{wkk q��r]�Z�M��`m�w`کa|aB�هĽ�Ӳ_����Sܬ�D�~F�X���"K~MdU���񓆔��RȠN�i!���c�����g�x`�tU�r�)q����h1�1ØiAy#����8�P7�w�t��7�",���Arʙ��P��,�!x�!m��*-lH���I��ό~�2��5sy�o�s��!��:�2��Ue��D ɂ� �ø�x�������n!�3봏R��Z�S!�E�D�3�,pK��I�P�8�I�٤I?ҟs�{r����Ŭ7�ڎd'�T�d&t?h�i �p*o?���d��ѱ֒_�V$w�xN��BΝ��Cz+.Hf�\]�F,wN`<`�8^�V�. ��)e��aդ@�Z��������R:̳l	�v��,el� �V���0���¡�7����e�w!�y�j�6i�9��y9�މ�Q��扖���#9ب6�'���+�;Ȏ/]�g-�X�����y,��L)~a,#�x�u�cPtH��>�C2"�����2��u^I�?]��z��wG�c(W��wu�W��5����(�!��T���<v��^gCN@�Ѐ���Ƀp �~`�,�#� �!@_��$�+�&`�J��|�T_'�mK-,p��k�L���
ꯇ���
o���D��P����nyOK�1c7C�$	�e4��q���F��ܸ�"Q��y4{͑��Vs�n�(�c�$��ݏ_ɲ��p���s�%m�z����]��4�]{P>G����z��͗�,%�#@j��@a�ܴ�n>����7?��y��-�o$y]1-]gC���);ۓ9M�M�O��_�5~�fZ�7ʾߟ}ɣփs@)|_)+oK�g���V+��m��)/�oPi�u�z4�e�����n{�
�S��b ��MNtVy*����ĺ� $�otuM5La���r:�m[�����Y.J 2�L��S
����,�ф�����7�B������,!6)φK��
��Z|��	�n�xIڻk�G2�4M(����%Y�]�o@˷�;3`�LrL̔�}k~�= ���W��c��r���eHJ~#�@)�!ؓ�HF%jQ�s�]�N�ݰ��x���CU�J��]b��)}�hnIq�KC�=��E���-��c�
����f	���*��'m�M��"�W�:��ƅm>�����\�^�����5UYk��H�`���x�Ҿ�������*H�ep-���C���#֏�XyH,\�D��ܥ>m��� ��ܐD����G&׈������/҇})����􇾚�)�.�aD�Mr��Ȯ�%�K��@��.<kl����^x��ã(�X�w,��əȇS���.�KDS�t�U����'��AՑ�"�yY*)&�fNP0�*��U<�]�u�A�^Tr�#Ƕ�Gs�~�h?;6�� }����lk��0d}��H�ha��ǰ,��e�N�P\Y�#y���ٞު�J��JSmV�B��2/�R��yK\3I%r��L��oX3$r1����-����bg��Lۨ���4˨1Hm�������;)��7���t�Q�?�=�!�,��b� �9�$�C��ޖi,u};�>����Iy3��D.gڀx8XM�)V�xd���;�b B�q�N�(�,�5$� ��Qȶ�:QZt�D3X��ge�2���s���쇱/B��l�q��'B?�L%�8�����
�.9ZC��\q��ʖ-V�?&����k7��V��7�9��z���F�ZKq�]2�F�=�m�߲"��@���� 6OB���N{�`�}8e`y�R��/�>CJ�X�'
�H�vB�[��P7�`�jj��\��O�#�z{E5I���<��8܂"�� �;����nS��Sx��a�"�j���8M�i��ø��1�D�UcQ@?n�X����(���at�'�����MT�i��$_��CN����f�A�S�]m7��򌧗�˃��jέ��}��#�a{�����Af�1�?�#�f���i��A~P���v���~X����6��E9 a��Ŀ�M�b�ˎL���G��lҶ�<��G����du�q����6�Lh$��	��ԏ{?�Y%�I����S��2��ϝ<7����e(c3�U�a��� �z]�$��7�L�ag���C�sIGC"�8%���"��$U<��{,$~CR�?R>����\{�m�Bx��#�7m6��k�qAw��x��rXEw�?NĿ{�8�Y((pR��.?yd#i��;�U/OV0Zi�X���e�NMB�)_��(K�)��r띅÷���"zW��FB��&X��������ź�T�i>~/	�OA��B��.����c��Q���χ���mb~��%�������3��h��;0�|�K&�	9{���#��c���'��;������-������V��KѢ\)��Ss��H��x��0�[�mω�Y�ᑽ�_/���6:����L��}r����t��э�=���~Y8S aymR����#���ڠNnԸ��G�b���;��a
Gr�dF%A�?�R&4ޟLGF��Ә��x�,>V��k�C�(uqY؛t���`U���];4��`]|�
�Lq���-�T�~I���V���2�|"�L�s_�\y�{���h���SE^r�'����˦9v��ZzV���4"�K�s;������&����'����
�WW�$��o�?�/�������>`�y��Y8���\`�n�-����ꔋ��oiЯ����Q�-?��;I� <M#���k�.���',&
q��d�o�¡|Q(?���C��mc�]�ۧ���'C����G�B��H $�{OMI
$���a$u5��.�\�`-4p��IGcS���r�=C��P��_��!�V�o�ȩ�x��� ��x9h+`��6�-u���V7�b�����.�y�?c��b����P��%�A��@#��&@�O��ż�C��[8S��ى�\�ڵ4�xu4��`�:����-O53�yCd�ۨ�wG�$��9�z���;�1���l!h[�Ý��}��1��d("h��Z 0eXƌ]�P�e�y�z�Icr�gST�zg���
�POd�w���	�O�u�J�XloJ�X:�}1S�r���k+mGt�v�����3�c�mH�6s�ަ�����_D9�"��
GF���4A�w.�����ްLQ�!��Sw�j�z�6�6�۶�g��X֢]U��7��LZ�$ta�$u}�^�w?a 5�~G5�Z�_��K�H���hL���v�(~sG���c�p�h��7S��:j�Uy{�?�Tk�r�1�"A���3V8K]��Һ��3�Qg+���_MH_������n.�]��
�#.��Cτj�N��*�d�}Jݕ�{?P=N�-@1�+c�+���+/�����.�#�B|텯�jU�Jrٹ��2���Z���V
S�ʒ���Z���CWJ'˂w���6���쑛#wM�� ���!)d4����e�����%�Ī��&��^w�=��
L���8�
��
�i��h"Vi?G-Atm����A�y¸h�C�F�k���*fz!���2�o�K���ѻ����n>r�s����� ��py\�����`C�f�9R��!�{�MŌL�f�XC�i�<5�q�ʣ����/�J��ي��Ukl�K/�c k*��XQ,a��}G;��p��M!�k�0�3�d�mscn�}�����S��ɸ-��}���[?ܝE��0�i;�&�3D��*��ÆͶx`Z��=-��h����Ϯ+��D�7iu����"�
�P��ҍ�D��@w���<�;z9ܹ����I��\Ft�̻���QCq�pm�#�7p�hn���:�)�t��Ƭ�.��N�:[�Zإ,"S���G�J����/у9ڱ	��Z�. �>uB��Xl?n2Y������E�z�<B�1�M���[�L�@��)a� %M��$ʤeSb��S��r����Z�C�.���	�+�����ӗ�Ds�%�Zǀ�Eb����K��A���E9$D!�P@y����M�LV56D��T��5��mL��8<M�@}�!t�m�OM�n�j8�)�>��_ʗN��4���>��(k�k���?y�1�f�BI
����Ǝc�Cg�#�hㅩ��o�,ZXO���|�]b��-'q���&���_��߷�X�c���p�qn�k�w�:eӰ�My^H�<M�c�|�s<��\�S)�1�W�����{M��c��R?��3�|�V��*��&g���J�}:#����
E"��2O5�%k�+5+��M�C�J����~�w�#?\fbq:r'Ș�z�>V���Z\�ڪa �7��8b��i�j�Ӑ�#cD�'%��u�4{ٟe=�8O�$J��\9�U>�@�Ã���᨝��2�du���:��e!��tr�E���҅�"�I�(vqڋ*"�A��6�T���0��͘{7�v<��&Ir�@d��A�LN��kZ��ז$YNi�Ȗ�x�V&,0J�qV�Lo.�k���xe��Ȗ�ND8�w��l�b�͘��	�R,��l�a����7��j�#L_����[lQ*�$�}�	��x2��-��/�#�V��+u?
�<M��:H욽�]����.�4�O����	�x�������
=�@��$M�\��>KÎ�T�#u:��c%�¯�S"&��$�hJ�J�	�-ߍ{x�����E�C":8�<�q���s2?�ќ�J�(30�<؏�b5
�|H�un:^���Z;���1��P`�GD���Quƶ�=Bv�rܫ����ˁ�Ǔ��o��7�s�dف ʺ �8=�$6O�ZF)��D�q�4��S
��@�6�vO��+ۻk!���0|�J�׃-�|���sץ�%u[���+D�0��!��FXh���E�XU��!��G�_/Q�.K�J�h\�A$�M�r�����7;�$(0f�t�p#�n�K1�\�&��!���Ǧ�M�2 d�1��rGC}����O@�sF�����=���n�)�xr�sn�&v�ˀi��*#s��N��}��{��D�cBǗGc7r0�j{���wk�vWF�"�~�7.�d:b�
x�Ơ���E�ĝ���b6���B��lq��Fj`4��]o�]�k����=�of���P��h"��3f�-]/�p��^ Ͼa�j�T����Ɲ�����ǂ���3�UA����|�:1���3l&�\�Q����Ǜ�qw<ß&��}*�����%1ƑHsU�}J�k�
�V\J����Ɋ� � ��4��i����@5og�Ǡ�f���HB~��#���ό#fZ�8l��j�p������N�;���K�b��:�����b���̰�8��ŗp8ް���?��N��8_�G�D�����m����D=�q���wU����N��/���S��#�sh��G���w:V퓲^Zx����< l��xq;��Zu�\q3+q+hv[�x��K!��o���D9�>A�y]��x&��k������mT���b��yżZ6as����X�ZBg�k�N$ ���>��@�J��(�D�(‪P��'	C����ox_��������F�[w��~o�K�M`��95�m�0��R�[�M���������8��6��-3��̼������`J��uB��p�+�*W3?��
d���"��,`ٌ9�o�A���+� B\/���|�� �X��*�B��2�$S���+e��ȋq�&A��5��y?"p�q[�fㇵ�9&����.�]*�9Hh�4L���@1�J����2͚}�#�CI�w��{v\!ew-�f]pkM��3nE�r��8��=iE���ت���X#g�u{f�I&�|yzc��3\ T�!������@��
�"�,�D���b�猼�r��s��k�F�p��(�^��DE���,�����Tät�̐'���8��M��<jj�KB�#}��>z�̕6�GAY!,�S���K�"��B��Δ���f-��7
S�=s���&��Tw}vR�^DxCk�qı�!�i�P9��[�m� R�8�#]��۠��R�O��`v{H�`�ٮѢhLz�od�����9�Y؉C;��q�j{���Z�;�_��T:-�n�[��r�[���&mL*�I4��1k
��[͑�'_�3�/�v稾s���)��u;Z��WɺRMɔ:N�� ���T%ss����^$��M�*��+���aj̓��ں�a&7<���q��w����r�;�V]���N��G23EX�י�*U�=�m�u\=^�YS��rE��A�m13��zRE�|֮"�'�ǡB� D�1�8��ݍؼ�~�1�Z�`��#(��#X"A�#�����v9�y�i�.S�$�=�Vǁ�8n�D%��T^b��A��=��N���l�0�w�	�
1j�F�W,dT��#�KR�&(Ա HC��C"[ �0a���fi	��)�(�1O�⫞��SOm� V��2��kk.ENͼ�v�ͿY������O)>�,w�3�/y���gV1�2WCB�����|�݁�	�jD>�m�i�#(�*NcRpY.+E'���H�u�t�+�)�}g'l�W?#۬L���ȇ�4���fWFH2A�n�~-���׉u`)���P�́��폆����[ɋ\��C�0�V*]Z���A�i:;������	
E�י����Q���O��@ݝ{�PbN�ۼ��\f�U�!��*L��1',�NP��qp��c�̵{f��8����Na�A�;s</��}�����? i��%���3v�7�^��J]��J��^�s��VK� [���"�b�&l�/E�����^yf��^Y�8D��16`ŽS�Ϫu��/��'�Kb��U��@���F?<�c(��d��� �b��,�u�#�O�BȰp*6
�F��&3����F~b�[{���^��{���#T��-]�ObF��Μv�"�����
ѵ"s ��b��~��2"1�t$�z�]�Q����'�	\��ܰͥCh/N14��Ϻ����jiN�������1!� U�0�c̋&��"#��&Y�q��͐���3�x�N��'J�:'��/wE�0�4��1�9m "r$��E\�:���A��/i�n)�D�B���=�����yU��銏�cb�]����0|�-�tLGrm1��7ﳯ�u�mWF�{62�V�ob�w�@^�M%//�S3�R�,�Wd�^_-L-��s���o�q,�v�З�q}o�Sx�a�|�q�2���9w��y�'z��h�a��!�	�/O��Inտ�'S���I��E]���Fh�NǋǶ��������Q"�X�uY[�h��[��`��x߀��/խ�]�G1��`�\a��·uL5��W�*�l1����l�#�%�z�W>���UtQ����^��c����ʶL�=�+2��">��:ZX�I�����O�4��S�V��
LE��J����oy��+gڭ9��-�_#�;�乔힞-��4˦����3��5�r�Կｮj��Nu��Sm=�T�0�Ț�m��@�w8��!�MHQ�5�;"tH���S��T_Vhz���?��_��}��L�{YR�%����jtч	�� M1����&a��ts/I�dəJS�c�VY�aE��������Qx�섮�6��n5�,Sz�q�c�';*MNT{q#�"�j+���o�s	�i���/��[%l`�������൒3�����A���n��0��-]���\�OLϓ��ϣg,�l3��_��m�d/�4�=��M@x
��/^8b�ā�㖺 0b���#Rnz+;�si@���:�Ɵd�����ׂx��n�8K+��X^`�fx�Q;�ܼ��f�AUnV\�1�~�j�5f&���#c/$�h��`�ʥ��iк2m���z�+@y�kQJ�܃m���*Ar�"���6��,v ��x.�n��W���4{�f�@��|�˵M�t���D��:{ �%��d�_��*��v(l����T0�?��qeM\�@��pͬ�x��c��.���*\�G���l˜�97�c��OO�?Z�1���=�.ʊa�
��2*ܕ���R��h햻f��J�g����Tt(�6W�b&|e4�`�-��;r�WҶ��U��Ru\
j�یq��Hj�]s�����@�L�Nd���xH��q-0�}\�Z�j������v��.�]���������W{b��}��Z����!�`X?Fס��T��jJ%��g�]Ѣ�lg�Q�
E�>X��rWp����e��,q��ؓ�ޭI�H�]��Ǐ��趮nNyo>GE�G�Mx���kLܔK��Y]����P�����:��A��Rb|^����S�׿.[.ۆh
�r�-x֜h�����	�c���ԛR��Ő9K�s&h��rጣ�]����ͽ:v�9�='�,�q��Ř+���U�p�,�W�-��R�ܗ��EL���_&92��Cu�o�5��pf�t�8x)��2���lf����ZUX>��R�H����#�+�^^h��-O,��1{�+Gfp̘�
�W'��HG�'���^,Ot��F��!͉�S�\C�X������x=sw�WK;��3�Xm�#��d#���Ȫ'��'��S��A;��mY�`�-�����>��ZY�h,Jp��#���ܺ#'��y2h�o*┍��T\#���0g�_���B�5s3���A�;��hj�gk
����D��ǫ�U[0㖐o������`'!�:7�4�'�
�H�dJ*ZǛ��<Dx���S��Y��pJ �E�m~���C���].L����0f��K�_ kc$�z镦��hMɜy�hM U��n�h��/�T%������+' �'rb�4��R��k�]K�7���s����E�Ԅ/XU��!�jF�6x��w��>k�r�ӈ2�C�T�/��d��l���h-S�mM�6s/��j��N���}��p�-_�p�v��c��b'[9�0%=p���o��
�3����	Q��R��n]<���Ի)M65*�A�H#���+ �?���F�U��b�sy�֬�(%16z�>5�9�)s�j��c�q����|���6Z�}��T��W�n��ȋdS��+]A����<%h
�G�~���R�*�	�/h" X ER�#	�����苈�t�LY�L�]��)��c"�uR}jqV9�F��)G&��69���䙎M8Fi7E���@e�$3Dr)���ڟ�ƀ�9L���9���u(��W�# _�B����nv:�X��X��޿�?zf���E.tCA�"��"P��s���sP\=ˊO�,�ƺT�ڃ%�`r~$23Ip�/S1;.����8+n�n �!��Sv���g�9w�ЎS�z'��E���am%R��P(�lP��e���A�<�����@O�"�ahU�ĆC.�}�"��<9?�oK����x���Mm��.#z�+�|vc�ײ&��`h��h̒�}�����xZ<{qdJ��H������)	hǷo{�:���_�BlC���ңT֌��`�%��)F�o~i\�g�3ۭ�Կ�}$��j:B�og�u����r/_]�#n����E���8O�DFX��E��FP����;K��k�0H�65�;��gKW�?9��znro͵���P�X����n��m���3iTvoG+��W6������Z�`�5#� ��#��%���)w㵍�r.F��+0�=�D���u�0�b�$���N.&j�?i��}"Vڴ�9� �7V
tq%���aU�9N׻Y�
q"q8@���b����;�2N�;��շ7t4E-�G���q���;�6��\:A���e|C�C,��c�X��7E,�������1��Ik�mc�F����lj�)5��Ͱ�fΦ&�Ň+��K�
$�lO�/��I���)QH�x�?0W��Tb&��T�0A����*��_(�Ю�u�{9:6��<ҝ�v�LA8���p���$Q`v���'�s�3�Z�-�G���1���=�N,�E��]��8E�:�m1I�����9�%B:�
�&�o��e	|����~��lֺ���\p����Ku�"#����m^!F��IF� vF&
 ��6��;!'=~� �5I�r#Vf}%̤�ȗ<<"t��ĘL�[�7���~6��������q�9;��r���o�;�Fb�	��C$'x䢛��S˹�}w8��U7����5�[VR�E���������M?��r�Ѓ��1�����6��j�>��^#��~f�c�g�J�ٴ֒�y�n�̦���/v���TΑ�M } �֠唑�]�tO�|�<����������)�Jz�����\,����Sc�u9��y|���G����J�,{b����PM&��LR�<1��S[��0`�8�9�U4��h�½Ǡ��D �\�aV#�n��Xe)DluE0Hߐ8�Aߡ#��3>����DW^���u�x�����Тe��rژ.:um��:6Wx~�g��_���a^��l�ݦ��|	�*9_�s����S�I��,j5�[u&�'�~`y�d��ٽ�|�!tr��Z�Ӆ�'-�\|NȒ��)���fz3�ЏK޽C�7�?5l�:��=�Z�?$@�M�t>�6�*����D�	����Hnj�Г��=Ð��w��Nu������yQ����꼡�d���� $�eMe���>K!�����O�*��@��a�e�E M���Q:(y+��E�
�t<��,���ə�
�4��]q8k�f�W�F��U7̛,!��s~p�<N`A�:vḪ�k�`N��|�1�tĈ-�Gʳ�/�6 �z�"��Ƨ^Z��Ý9Y�UM;���/�9W���mӪ�f7�w�]�G�<��\ZeV��X�ܔ�z#i.Y!�8��<��P��n�1� ��jڇ�N�U���D6
�rK�ѡ��'u�	u��g���4����$�!� c�P�@�\���=?: ���E���#L6(q���~S�'�Aw����}m�	pf�D���>mc7��U��a�ZPB�����J;W�vq���<��f�ٌ�\�P�/����yӴ���&m__���h�p�4���������p
�������0h�ITw3�&���(#B@$#�ݔ/��r�ű�M\S���@Ka
8���N�~�.
Ean�֠��K��?���^�b�'i�GX-�RuJz�df�@���0�I~����_3��;ԉр�HQ�8�(�(m$�ak�R�f�����+I�hQ���$��7S���:%�R#�����Z�hR���<����8�r��x�|s�&#^r��$N��d�;�s˺B�#(f�h��}cv���g�I*�}?'J�7��ѐv�콖�L:� 2nŃ���f��P꥝����٢љu�0��w���M
������|�tA�I�+�qqq�һ)�R9�X���=>�Ve�W4��^�/6@�q99'���y�IIl�F�N���Dj�4'��}�d!�����8��}*$*0�����#X�*�[�d(��� -�1���Bvg�e��aYK�2�ٟKBy��	�Z����Ŀ�'q����7��Qi{2H��w�B���!sl��৹�#�c��E�TR���ٱփ)������1�T1g���l�@���OB�<�&�q,~^�����d�����d�+|" �bpf�>�Iur��L��c��2!�p�Y:N���3�>(�:7��Z��韷�	�B�m���dP۠��S�u��@C"����k���҃�x[`��7Qr��G��ݤ��y����ͻ��[!;��m���-+��Ġ�h#���F`v=����V��@�����L��gX,(#N��R��ءz��M�doϴ
w:0V��� � {��O�'eq��	�b^H<p
�N���I�@�L!k_�ڃ�]��BrP�v��Ё��8)��1O� �>��rm�c�LrrF/�
96`�cUi������T.��~{����yf0Tu]��A�d�NJO����F�Z�5�{#ｘ:/F��q
Y�o��ls��i�X���^-�sߋ�a���0��P��담\�V���E�	g7{#$^�j�"Q?�9'M��(�Ȋq�6m�8غ����4��/���K؝�?ss /r�[�8�ύk��\�Z2�Ga�9"X!��������h��_�"p�~���s�g86E�>��9�ɕD���Z9���� Bw;����-�"î�
t�@�l�sZ�y�Qh�YC7������Lq�y��󝘄��`��~��9�;�w��Բ3t7<�#���?�R��~�b]kT`����mmn$����J��T|g�̭�;u{�R|��"(�Þ��!���h�|Zn�,�'dk��{��h0DΜ�4"�W�;�{}J�r�ü�A�5 �`��]��@��/���%�E�b�aě"��78�����e@�=�D����ڲ�K`%(�R�b��aq�y���Q�Xꗽy]H��XƝ������jg�*������)q��qRȻDo��d�W|EWQ1<~�q���,�.�ҿ�����6�9纙�~o�8_��s�]u�<_4k
P{�%;
��`��)��Ut�y�_�B\is�v�iY�
/�_��\VTi;�z�"��C��>������ҭyYk�6/
]��9#ј��2��?uY�5��^+�q��/=�'����8�H�m菡��=�T�a��Kl���;�'��#��o�F���f�&��R"=��1����Z�~��upv��D�]���Y���tZ�O
`a[TM\��<�,�"\��]V���[c���
�{�>�eN�xW���"+�0�Y��a�u�Y�E,U��Ӂ-��^����X���Z�"��Hv�S�xJ���.��$���n�Γv~M���Q��_T;Z�'(h*���V�tb&$(���˘Z�wꁐ�tP�w���8P���*{&~��E��������Ϡ�e8#_��$�������6/�@Gv�cz�U,�n+S����\�+�ֈ�b��?��&L�n�̠U`����#6D��Uݮ�A�wļ��_����)�Z��	 䶜��϶����6Obw�v̾)��5�M����ߵ] ������]0D<Q�'��"�,�'fmR����S\�Ks_����T�4牼����`1]������k��ܫ8��i3����D�
�G�7%`����,��X�R���-��!3xʂnܭkl�p\&I�-R���6���t��QU��R�"���ap��J����2Mz)���J}B�[��\W�ڥ��>-�w�H���tH����/?���4�i+���_��K��fz[(�Y�}�z_}�=,�?�0�M����n\;X��0��z\��_��U���s�M�3m��F�z�a~�!��}��	��'�t_���EA��a�4y���[��Q�FkK�]�j�,#G7>�6H;0���R���_�c>�%�P������vʗ�ޕ���Ö�;�4e�s�Xg�'�J������|���7v�z�l	9@oܬ����#��#?��k��B���ƛ^~��~�rg9��uX	���{�[Pʾ��Xh����d�>����M�a�<+h�#�{2�%5�>´9%t鉡LFW�ˑ���Q)4t(v�'��f�ݵK���M flo�n��F0��> /q��u��5~_�`(����$�md=���gK�~�	�A�X��w�QV���d!�rS�τ�vZ	�r���{B�}Ř�S�����?!㞻�<��
Pٕ����0C�6R����Ox�Yz�/V�>y��.�����9�%Y���@[2庻�5��iz��d��%�_� ��������ǯ�8fc�h��/7�Q�����$4���\�X)�����LĬ44�
'���׆/�R�ዋ:={X)&�t�+�8�K{8<E{L���cn����1@����6C0�&��V�J������r��c7ܴs�%1��/��_�I�|{>[:�07[pK�nל3�}���q�.ZŅ.��}>(~^Ԯ�}Q3f�r�Lv&=C$ot|Ju/�3ٓ_���ҖUr��5D��A3wg��[՚9l��t3��Yk��ȏ���x�1g��zռ���)��pn-r�H�|=�Ͱ0�;�s�=pk�a�� [��3������)��i�ʵw�\�D�b
E�hz���`@>�-H����<~���u7�
����q՟sت����vE��j
�k9La��j���<_�ӂ�M5F�em��%A=m��S`���O?�aq��C���^����E`�
����A׶/k{ ���'i�+;�F�t"���2�ii�PCO���_y�E{)��n��̾�>��i7,�Nq!���l�?�CL�ɰUg���c��q������֓�>��NEm{���L*�w�ۑ�u'̩�$�#Z�r�#W�^"֋��o ����}�PwB��[^x����'����Ô.�����q?E.��g�u�S$9�������k�����pʣ�v8�dt��Kg��xq �̆s� �	�� ��bP�V���6. �Ј�"p9�"Z�����J����� �>�Nj��j�ٚ�=��w=.���N��Z�<5j�́��2~^Q�`.��b'�z��OX��ۘK�7��Esi㪱�u��ژ��F��;�����Y`AW���P� TF��aA��K��*�
ڥa�gFx�Z���%��5t�u�&x3�
��h���,߷
2>�I�|��!��x�X��s����}~�M��Z^��.���;m��7���S�J#Y���l�yI2s�����ج�w!�S�˲_<蝛�~�l6�K�Qq�dvL����Ї�"���MXj�v��<L ?D���:�:�M��_��Zӄ�2 ]����ւ�7��C|���\�.\�� ´�i�N��I��n�Y���C�@�%@�>�+��]���XZ����ʢEy6�fE���"�:-�y��0WfP>�!W��g����H8O�h���
�*#��5����ч9�v�8}��7`����V-��U-E�N�jÇҟy�*U��]�5Zt�W��T�KE4:���b���$D*1�H��/&����KX��G���HQ{ϊ�b���������Y��B!�;�䊯�?u��J(q&Ϯ�����Ah�բ&��JIx �b7j O����Ut��pZ�����$'��%!���;�r���W�s��S����� g.Ā�(7��G�(�[KVq�9�(�1��f;y'2&^	۫��͛p$�֙�ܞޗ�|���§��Z�~x]����G���r���Yi�b|"���z��],�Bm����?��*��)ر��v�ek8&Q���Ԛ.~���b5�`Al_������@����\���)�tʹ��yaL� �vJ+�0��:��m2��}5j��.Z��Q��ZM�, s��7�q�
�&	EE��2̓7�"�4B��P�_B�ϒ��]�����H�^����.��s�oG����(J��D�E�=tA�lD.�JZ�i��}����1��0�+����`{�P �����ER��/�~��f����	�hkҬ{�EҮ�L�BW2���c�Q0-��]�̷��R1�>1CI�˭��r�RIO��w,�*e��v����=���tR+ �]bہ�l��'l�e^�lj��I������s���<��ڗ�M�L�x�-�.wi�?��mM��\ϯ����JK��3=���Q��F�G4�fiL��Ukv�}_cHr�]jS�����U.B�Q��v��v��(Q�,�cΫۿ���j5��������	Wc��C����w��	�$���I�́Az��c/�>�s��o��+���e3����O1�w@��w��������ة%/o�!蛍P{^y	GFAĻ߰��&����iY��ɻ�,)��,�m0�4i�(��z���6��JL-�7���=�lf�>ы�<��i�qT�5�lu-1K�%@��v��O��;����/K�)L8o���AX�U��Sj#̜�b� ��X>o�
z�a�t��ӹ���1I�~ߝ�f����ƌ*��z0�����שF"��������=H�d������~��[�8��l
yz������S�bYr4�j��QES��#�Z	��3{�f�ԁU����R���j��?[:1��ɇ�M��w*�࿾�В����		~��ࣦ+V'�:R44WU�tUt�����V��x縖��B��>�_e�X+�մ�eE�-���'�;<�������x��W9���o$K;�:Vs�W���}'����Y�˷��\�!��kl]���E�cK>���b�fH��E�ڼ��F�@�bJ�5��l���%D��3�?�	I��\���5����KO��Pl_mn;	Q[V�:�_�eM���0W1t���O�҉��|c�_*��-�+�_��쩗љ4�)���y�ޑv���/R�5��h�ɭ������'���e�1_�3W Gs����~P%��w�~4cߥvk�e-�{��+��>��E�	�?E���A'�%% '��e�Az��S����h9D䪒����$�Rە�܍�96�C�8�Ākɩp���殈G&�����Đ`���iٸ��o�9�+!�\W�>�O�$[W�F��:�9mW����� �`�c����g�ԉco�a��ʂa����v�V`�H~3�h�)nk�D�h�[�`�"g�j^	V�%C�Lf���ב�����{�;�f�{���Z�%<_�AknqI�U�g#�Qy|�F�{%٪���p���:�V�����{f�'���B0siXV�	R-0�v���T&jZ(6S�_7�`s��69N!|Xw�>&C��^�ê�� U����	��~������h�A�A#���!\R)S�y��a�[Xx���=����/32i�k�7 �(�H��z�c8��"��c��ؿ򥵆��qK�pv��*L���k�V�0�7n�"�**�=�B������^J�fA-W��ϓ4�^<����GuSUk��-w�Ö˸=w�i�UEA
��v0�
QC3G!�F�@�����R�\>�Wn�.�|M�����
ѧ��M���i��k��+�@�����1�/F3Ye�*��d���J����=�V�2�0�H����N��E-���䬢��[N��3p]Px{�!R�lA���]WV�ƒ�kc��;BɤJc�>9���{b��6ͤ��׌�Y�\��'�~B�I�.�Y-*(ȷ���{��a�FFً������,!���'�Li܀�0jǮ��yq2Zt�f1T�Jf�}�tX��͇k��p��3��u�e+_XG�Q�GS.�w�?w|⏳�T7ǈ�;�
<�gY#H�a�T*N���2�[A���xh��.�Ǳ_��ۻ�k@�]�c���bR~������X�$JAߺS�Hh�,Ӹ���Y��F�?���Bv{�q���LY;#��}��;�����ٔ/\�����4"��Fb��9t*�k�*�	��ߢ�瘐�����	q���G��
b[|T�X��מ�ĕ���`<%L��S&s=�ꄙ �ٵu,b�/h69����&�t%pD���N,_�����O�[9$�]�at��)� �Ȧ������s̫�ƒV�N��}���B�{�8H)K�{"l���reG����!<#�b�ϭ���ߵE���,ڠ���%K��'"9W�+��p@����qvY��I�P��$�]���9����jJT��9����	���#��}� ���4wY j����l7K�9,����Tj��F��iT����('b�)B��1f�$8��{pm��>	�� �T�9>���(	��`MH���f�����y�-/7<줇#�-�G@���d�S��J���@��`ޔ�� Bq?���*�7^��q_y`$��&��ܿЪzc��a���/5g��fO���5���$3��^�:��4�+��[i�/�H���R���tc��y��TaP��ҍ"���o�`	���̔3/=Ra��J0y'����u���WAMļd��cb�d�N�7.�E����h�"U���p���N���������m�'�w��qj�V%!=a����+�W=��?�?+"WV�%h�]ю�l%^G�C�rr��?�|ʔ�/�>�Q?�!�,/wk���d��J1�S�H�e�U�<Jg��`Lp�qTCϐ��D�}���c6al���!y^O��+������T=�ǒ��
���&݁��򿯮�Z̠(m3͟��=�x��]�V�N����ộ�F��Q$˥�B���!hN�ke�~
J��Nzzݿ�B��xI�~K������ДfB�T�)�M5�y��P����������mh�?���椳��`,�������Nh.k��)�����[���|[w�ca�U��;J��tFm=�I�ոp.�0���0��3��Ȱ,�t���$y(�i����=9%�fdM�SZ�
mF�,Ns̓x2-)�=�1�Խ��zao�x42䮥I�g���S��+�C�?���<�8e<���R0Sk3u����aTfGWPB�8�mG�<��kH���y�Q�U�u �}j�;�v��ņ)�(��Y!؜���'̔Ok�b��Y{���o},?�O�k��OT�����tX54x�Q�3+g}����V�c/FcΪ�ʥ��V���J��}�#��cl���z�mbD�k{��^��b��܇���l>4�I]g�*�1/�)��W�#��W�o_��"����^\��뗂��,yy�Gu�7��M���:[P�:#����V�ڢ��POQ��
h\G�=!����=}	���I�lx��x��M
G~���h���Q>վ���Z��~��� !����{����U��=�#���'$S�̳$��p�1c=q��ڦ]!� ���%����6��.}�������
�r����BF���6�w؏@�]G�O"�;���Zm�
�'���-7Y�$
��Qrȡ���Q<��O�`��u@Fǭ�����S�2�DB
+��HD�ڭ7Ki�5@L�(5k��[���*���E�z��_cV��Y�9W-���L�-,O	c��<��� :�s҃��u�4�2�-L�^hI�q��\'Ǫ^����а�2rZ�p��w�u���!�x�/���r>D���h#=m�HҜm/U\+�q!��F"D�:�F�H��&g~�0�'�h5���Q9��50���1/
��ͨ>�T� �c�C����%���V˟c~��$dg������	�����o�NC.�%=6mk`���0I�۟��������	B�+c�[܋�A!�������.�ҿzG#q���Ι�s
�~��>�Ԥo!������76k��)S،�PΩp��:��� <բ����>
�h�@5���Ϟ�9<�A���T~%,f�Z�Ǵ��Iď�A%���T�C����Ї�w��؊�"L��|L��6��з�w}��c���ј��?I��6x��#_�����el�����Z����?_X�Ld]3A�N<o���9����ȟ��Pk+3a�f�n�\�L�<[��1��G���ri.>wJO���@z\-��Bt4_���fj�O�Z����B�R���w�$��Y�L� �%g�E�`��.,u�� K}�Xvu���B�!;�����]1ݤMO9b6�ΔRq~]j�x�-�벼��	�W!�].g��	�T�a��:27a����9���c-a�E�W��M�繉�r�6���5�G�j��愁���A�[��K<��c�y�����"hiFظ�g��X]T.J��.B���9aL�g�@���=�	&���:X���sQV
�gO��U]�g S���.���� v�c�i)�J��M�O�~�W�^���Zn�8�����c`�kT������}�EQ�!�5i�������<��
����J~�*FMBD�ا:0�1��0��c(X�!J�������]��e0�kD ��'���>O��2-{�[�����I�:e#���H�,tHbVY� �D��C�HʪE���� �]Cm�����4:q��0�x�@h��@ܖ�D�� !���d��;��p�J���`Vt�J�	업o��}�kb[�όa�[��|͗ \�����U<"�8�xh����b
�:��J�Kϼm"��t�����~H���d��2Y@�ds�gam�1T-k+"�؂bߨ�������<�	�I� }�b��[T}ɷi�B8?C���껴f/�������!|r���\,)'���ȩ����܃)��W�����V¿�ϸk��>8�C�{��7�*5�Tx�$s�g��Ү����'d���?�nhx�u�����^ش��J2��n����q-M������7օ�/9�m�
��Ma��	�S���fH���;
`:#�9_�}�έBK���j5��J*h��p�]�7��IvM���͕�4n����P0W�7?�5��b��ǋ@�o��_�'Ȫ�K3duIrXa���)zx�V��H'�k�H/�MW����U����m� �b=RD�*%I�`3�
���_E�+��[�%l�[Ml�_��ۅ��y8߱��S����{��z���pkW%��.-����]�H������dNw����{p��1`
��R�抐�ߊu��ȗ�G�q�Z�o(��2��."�Jd��z��	p.#��G�"�#��bUʗ%��'���:��/?�xMpўY憥��w�.�
M�gZ�h���6�` MW�]T�'���*��5�����"}D�<����t����*K� Vծ�����U�x;�)+ʌC]�?�.`�}lN΋��9ͬ卞����l9�^R�Q%g	sR,�ya�k�1v�>�� XR�2�+AXmχ�>�>Tj��[$Ufnժ���
Il�铝`�\�����5�;k�p%��0�۸��g����Ɩ_�7m�ھ��\5_��jc�tQ����6��g���ԩb�;��"�-@���Yn=���1��B�.���~���O]_!Z��4ue�mf�����gzu��X��Z)��]��d#��˸UvP��U��Ƀ9��#�!�d�65���#��!`�J�]_X��gX��~(̓�����%�Buy���05���2_����$2����KƢ&�dG8�U�M�B����$APߕ��1" M�Z��4���=�s쇑�����Heْi��f��鴑���Y3qT�of��BM��#�P�g��Nb�KtB���m�/�N����� '�!S�x1z�I����Ň/��h�.�e|�A�$d�
Z��fG��Q-�7b)ZV�u1r3j�B
�U��E��zr����A��m��u�b����\��|O�*�3��UCz>}�q��;o�'r�Ϋ]_B�F�q�D�wS��|ٻ���P�9|�N���m���9.y�`vQL'R��0GS�WO��H(6V�C����r��Z�q0L�S���N�Z���'5֒F����8�YO��'6�~20$� n?,̚m�o��,� �6�с<�����@�gzL��uxS�|@��^h�Ɨ��(}*N������{3�* �Qk>��LW�&7K�P<����	�r)k-2�	�#��l�f�}�;}}е�����N	߶�8�^�L ��$�?�����\.�cC�f��B�2��[�ϛc`��+O�V�l�4�le��
}�~ε쁚T�r���nei�3\H��O����I�I�K�e�Ȭbw<(H��z��$�D�ҟC`�aܮ3"'3/R�+p⪄-\�{��#Օ%�0^ى�!�Xz�V{�]��ڑ�D���cGxoDV^��ظ�0U�e�@��r-����¸Q���1�-�.�wXIz����-v�Ggr&/Z��wϏT��+K��GU�����L��]�U���ڔ.��o/ZD�ҷ�����Ơf1f���w5�o�!M���zgL�.���N��uK�������+��
xi.���몟��w·��LL�&�L�s���<X�����fX��v�}w>��<	[�H�R�]JvleT�,��NL��	�[-:�o��j�s)�����\������F�����Sl��=��^�b��!B�\�9R����j�u��Fp�Q#~�4����\������)��'���?1��lVƂ�3-�,I�G(%����8_w�v{S�F&h�>�Er����_>��%�����IG�U�[�OC �qϷ��e��8s�`B�d2��-<j���d��%�RB5�ﴕ�=
;D�+L���&7��`��:�V&��xHՀJ*�C»�a�U��R}˲ǂ3��4�ܥ�#gm�<F2[_��ȿ#�	$�q�"#*+�H����Cq�� EW� ~{�b5z��?4��̼̅G#U�}��
�8��CI#\��o�T�!]�˲�~|����KHWY}t���`�8��p1�0�:��xa�D/uj/Z������/2`o�T߯?������y�o&E��ZP[,�4rr<x��ea���#3� ��h2��Twk����}I�?:��g&}���A�OH��R�]��5�7d��N�DSHz��F��+����[M��}����������s�]�LM3�(�X�:�Vp?A����q�KwT&L���z�I%%�Fԩ�!��qt%��f�Ja���ڂi�?�u5� ���s�CҞ��ΪF�CK�� o���יP"���Cn��=^�r�<X�ܭ�ԡ�����)�O&k�8�yBﮗ��77p����:����
�1�����/�ӎ��+rs����<�!F�#g�j(BZ�0~�avRi,�Ʊ�KKd ��m��Ѳ� ؈U�fdۡ7�*��Ul��Kҽ�=�	��;aI�80��Ty����;�����6WU�or��5�}�D� �k	���3�f�ܚ�L��ꭓ6��Bh<Y0�u����IU-��T��rb{!��ŭVIu�$}?�����d��>A�ڪje��d�4�|U�Ǣ��3�ۘ���$T\A�ժ�p'R�*�D_�L�!YO)��_1�
P�$�쇕���kv�p������kz4c���~�O�Ũ7~�������5�K��d(Da>%
rQ΄*p��v=�)d���&��O�=��r���;[�W�)�4�[)�4)���9�iʦ�^D�I���r��g��K�_��wO�M/V�������Ⓟ s�8�^����Z��/�J�_Eqo������/Q�b��m�(�aV�Ĥ'��;4t¨˒�^(�D��)�_�M��˩����Ӻ�>��+�
��8}>N+5s�y�M��7�{���I��Kz��#דΥS>YmM1c�` ??r�b�Ɛ�0OW٥eS���G�,�C���p��A������������]����xcf>] )���]SZ�	"��s��5���-���C98h�e}W�^�dD��;�����fI<~���2�J�_�����������������9�����kW\��؃��8~�ؼ�5,�`B<[�Ư"��S�v����߅tǧ��96�4b�1i��.��P��ܽ�q݉������F��Գ�_	��7�v�hY�BQ���#9����sV1���K�-�Rz�p��������~��Daŀ��F`��^U�pO[^a,�vYSDù�����^5���9��w��_�w�_B�$"�E��S0�/�C;��#fp�4-�0`dѓ����}G�����ڥ�aOhX�7�1����X+b_�mZ8[�;�)��񽯮���O��Y���tB����΁*ʬ{m�#[ۅ�:|
��:t]!0�����n�]`]��_�� :��GE7X�He�! KY}V�[h��_������5'v��W5`xf~ћ�슍4͍�<V�x�xH��eQ	@⦠<OE
=e���XM�{0�G�A��fv21�a��-Kr�B@�nJ�'���G�J7�z[�ѫ�*d7]��.
���-���,�ѥ�/x@erb�d&��s�Xm�����f�a6�w�Ԣ���u��3�g~��I�1ܖB�N���P�I_&����qެ�a�qٝ���B��cm�P�#Lu�P*�F!�XT0��-�b&�Cʶe�2��.j�ꮒ�#�#cƬ߈h)�طA�UpԁR�Tr�Y8	b6Jө)�B��!�QX��S#�zo?��;�k�"�.��x-�>�s�)z��VB�M8�#8�N����>Hw�I}a�ʊ�[z�N�f(�vH�HF*ߺ�઎6|WE�5C]��.X#'�y8�$K U���[��fk{����䱊�4Ѫ�"�,�Օ������nG�8$"؁��r��=��#@؞j�t���.C����g�N�J��=ۃF�2�B]�D9b	�����Xp����+I[�C.�ꦽ�?�{$��R��m-�E�L��}�[i��o�O�-�GZ�����&��x�ۄ��i���B����]qObz��%�Y��f��t1e�,����1 Q��D���,�~�q.%���ӄ uR����ќ�]��Yb���G/o���Mmw̬'CN0�Z�|O�+eq�� .����x;I���W���]�Z��d��`�ut�ƽ5u �}�d�2��/#�)��"PQ��y���*��u1�K���r��Ž�鸳�V���A�*��Ќ���#9s�K�����	��J���Do$5��gvD�[*�H��M֚�A# e�n���R��>� 5�ST梏�a�c��]�d~m0mbJ]�q>���o���J���h4�8��_IVDQ����k��7�_^ĥ{o�AwY���H���o�Zy��ʿ�����WCQ��	���fA#�Կeގ�wHm�z�c��6?�[.{v���V�Y�,1��U�$�i�{68j�i�w�������T��-щB5�Ϳ�xV	�4xx̞L.�\A5��jMf5O$�`w��S��'������	���ϰ�%R�GO��LN�?�Q.;�s]����g����Q�1���x�����)�B7(xu[*��e�=
��������R/���~��a�9��)O�P�濶lp����3L���O3\�~�&�ݸg�e�$���h��<�(���[ln�/����wֻ���l�D���{
m9��4���h.��H���$����"e]�%�:i"��EQ��}|s�H�e�췟`Ő�5k���j��c�j�˿GB���N@)FJGL�0�F�>��������&O�71�%��T��L���H[���aʞ_�x�O�Ḻ��zϥy��/���l�%�rʟ��)@PU�E�I���(2��V����KF�5���~�)����8b\�99�P�u�v���T��M����J�r�?��rE�\?�����/�i�c���IK`��~
 �m\(��k�Z��Z@�O�C(@�!E�0�	E�6�N�9��_&��C���}l�T"��z�5�ZM�i�y`�\����a�W΄��O�_B�ԫ2�1(�^�zSNTo�i��3�
����+h2�a�뵒�U�BT��b�r��~I(�Ձ���(�x�6�Ӕ������ڪ��0�Z2�E�� ��w�������|�P���?��,�����g��(��/�:(��x.�k�3����z��A|��F���3{<jo0E~0�L�46�����@nrx��Vp~-�f7�V����Ob�Rr:S�Ŀ��ߞaо6�Ҳ
x�����q�4�r���1�o$��2p��O�g��F.����"�؋@L�&s��:ѓw�f����Ȉ)�gp(��\'�)y(��Fx��R9w\�� /��3
̭bڏW�F��@&��y	D�Q`�y�!��א��i�u�lb�&A]f�n������_
o�W��� ��{����R𳮵����S+��a

/֒#��� �?-���8�C��LWw�R\CzPJ��O�F�s�/A*[�,���"̸�ǳ��=G2z�H�h����i|�?�ghV/����١�xx���5(�(���V�ruhd +s��zML⳱��(H��ד�MN�e��L���
��F���\D��*��=-0�5��]��ƽg����h���ὛV1��/dξs�5�|������n�� AM�]��@f�Y8���l����k��Ҕ��]6��8N�a���+}��N9m��d�㊹�:�O�Bf�`�Yّ�C�ĠVh0nm�|����;�\ZK,�X8%/��}�������ޠ�j��z)���P����<����}������~����`��_j��o3	��5i���d2�M��pRw*�}��v��⍜o,iuk��s�tR��|J!��8{-v�3���9�f�-����OS���Eő�}-�XVt��J�w��R�h���qݘ��A�i�q!_��ԉo��H�����޺@;�}e:.��ȑ�k�����ux	u2S�f�K�
���V���RoG��8�����y��enaK+��D���%�]ƻ�*�X��C7l��l��(x�|����NW�2QW�Ӥ)�%���l������'q���#QSl�e`���74��<���3���#���KAӓ`�Ԋ�������x���4���W��φ7�0D�Ϻݮe�
	Bj�x¯]���;�
� +�S=Y	3�*��~�����Q٫j�������g#��l��������_9F�:ZA� �ƍ��cI7�|��}�	��`j&?Y���xk�A`��3̫D�����k1���RI�U�"�#�����Q��2�a�\ă�@!�Y���!��B���
Y�)kY��y�	�s�+|ye_XB�!Wj"|���R�V���]'���y򏄕�ń�X�K��Fн�`���hK��3s���䛓W�D��p'>0p���Bm��tq[�Je+���Y	`1X�I]7X��7fݗJ�F��ã0��m�'x�5��g�9c��6����@5x�Ɏ{u��b����e0.��ۂT`N�q��]xnt���z�%����_�<ﲃ���d#�'�ja�uNƙ[ub(��;�g�,�G�$��u����m6���i*]����d�4	���v��;�HU�����J<im�]U��b��{�_= ;�deh�U�%	 ���p�w+m���V�����7�-��_2��%��h�v��2`�dd��_��f<�F�f������{u�,�|A��U�7L�<Iy�b��B�t���&K�2%�ەER� PL�P���s�P���v��(U�C{�|���u��[Vi$F�El����y��,B�[@b-��Np��*���t��H�_��vYj��'�.ɕ2 \�z��B ����R!��*�<ӻY�L����Pd�o[�6�j��&�y
?�-�R��Y���O�j*�5ę��!��l�A�,�0iO�4u$�Z<:�`���=���4c e	)��l�M��(ǚ ѫ�Ǭ��kɏ�\a��Ѓs(Q�cІ�B�T�1�K��%ˆ�ER���U~R���4�Y�J��B���Ǭh��ˑ@��E���]G�4�gVQ�L�ݔ1��Ch"Ш7/��vg���w��fr��8�mo}bY�.Ղ�;-��'9�Ҵ]�a,R��q���������_sC2ƱzP���D�=�S�剨r��ѿ&�V���:�7�T'h��aȄ��lW��$�w������c�g=���u�,U  ��BFGX�sX���![�����	�V�z����e[����V	T�� ��������i2Um�Co`[���D�w:O��qG��W]�%gn��b�(�/�]�2ۮ���#� n���I������1�vM�5�9�|���Ç]Z�Y�С�J�nػje��� ��3şe])#F���-����Ľʵ��(`�0�߆��!\@dt����خ ��Y�Tё�T�t�r�3~O<$hzH�O�:/hH~��D���A�:�B�z�,$��h���)����Er8�^B�j%�M>�˒��������A�c�
C�(Hal@����Ga3ê�.�pEG�7^tL�Xv���FJ��x\��A�#�>q%%��]�\Y/�\�`I��i�����R|���+�$�G�7�Ғk�ЦK����q���3~k1���F�!؀�6�y�C*�$��!	������q#t�1Ֆ1E�P9$t���Ҳf�c�A�?~�w|}Dd������"�'����Vڷ��ɷ����q�}xצJ�Qc�b��;߉)�6T^�!eU���
�Bj+�h�݀�
d�X��w�I�.�)8=�GF����!�N ���c��� P@��|�<x�`��E�s�ǹ㬟�/�z��n�,nJ)z6�t��D��ڜ�+ac	%��h�jpEi��$���A{+[�J���6ѷ��@�%��1�[�7!v�5��/f��A6��h�^7[�3K�bV��w�:'ު<6tO0�%g�e2'{�.���}%.}�y�*�w�֦�F;@g�!�d���(��h�h��	���h/�4�D�O�1м�������/:<��~(� ���P(:�M�nbBm3y<Rh���US����/3�<�@�Y2N�X���&������A���Z�j��XU����֑�'�X��8�J�Bhb��^��F$̌6g�]�����,~�BQ]� LM5���%C�Ɏ����K%M&��U���(��-�F��i�#o��aw�8�V��ZLX�ͼm�IՑ��d{�&�9JcI�
Ni*g�M+,�f�Ǉ�X��C�O� A���[�D�@�i�$U���B8����Sq���,�47*:����&8���:���_�L2��ǦdC��^��4}:�C�~]�E!�
��R�F ="�j`�+�d�t:��������1���	�������f�7OM�|	����u���G�'|g��u��NVCɭ���zXud��̀w���!aU�_h����
l�$*��4��X��5��f/14��ӽ/{�7�D�jh���#7f�(i�����a�6�7��ei���  ���TLQt�����7z4]�/B^�@*G�M���Qc���kt��{p�:�i2Q��9{73)D�ڵ45Zý�tP��i��/'�R��(,b���V���񹱍 �	1�AHMM<]f�_;j폞��[9l�7����(�d�fe��0�M�L�����r�́�8H��7gG?A�pTk�Q��2;��hS�{��rꫪ4��3�T)�R����`]�N������-���@������76�;)�`����;� ����a�����t��\�I���`܇?�hg�[u�W
"_k��ud�:����|NB�sj+�����;����f�O�M]�X�q׆a6%ԙ��L�M~�D*�~�z?��l�a��\�ېr�a;�}!��m��<׌gfSd��!j�׆	Y.)Es�U`�(�D���W���%�떧���HĐR��!;rM{���#�g`�s�%���&���`���a�Y��d��>AVo��5E�,MP���8f�{\2���&]� �D�̈/ȆMRH]�~�A��x�*p�y�����G��C�5p"{���zsԩ�F�!�\�xY��
3M+�c�<���k��QEaI3
�)�}�nh�{�Z��a��C`˩��?�}Pi���x��Id~oe����BcL��� 9�NW�?�����$[�Ђ�j��%?.7�#A_.���/�kշ�0(����FhmzOjI�۷��k6��Ǉm�w�� ǜ�[F=�g|�%G��E��uO�S]`Z��$������'�z��tL���+�rs%�1�J�u�I
I�sd�L��HN�*�����ԎY=����Zz��n]=�uM�Е����0^˔a>kc���|�%���MY8�C��?L㻏,�A��J�m=�z�,V/G�E�Ȝ����cM��?�'T�tZ��I4��yŬ��_Oߝ��O=r���愤�0�����ai����~l���ySc�c<(���X���c����W�RN�3̡���P���g_r�k_|�!l9���pM(~���2'�����m��9��~T���ͩ����괢�f^��k'�(Y���}S�{�t�0Ǫ`;DD��b�� ��y���/���B���m)Ώf��P�;�d�Gk�S+�I�Ҧlq�Sq���i���-�VZ�w��{��O�Z'mE)�?Ր�~�s���t+��к�T߆����n���wfF��4�ݒڊ�/ɫ�i�û-�4_V`i�CNݺ.���,��
��f��kC_V¶�a�C��>G9y)�=��yl�:���^�����?��P�9(̧����4�ny�N��12S��Z٤�_���ϐ�����U/>D��;�m'kc�UJ���gV�z����#�5_��3�Ɣ��L>L�:��b��8uNR���K6���Q��]\�f'�a5�M�z,�	�N����$��<x\��}3rݳ\8|��ʩ9w�j��4��d/'�p���k�r�3.�M�,f�5�-���5�PQ ��8"�C����uiJ��J�S�	z݃K�`�)m�Xm�F��2S/d�9���S���δ���q�Q��P��.������9�R��;�*�����+��5��b5W��̬��.䭆�F�/�e�j��9D�P�� ��W��;�D�������H�������?u�b#|�VVEc�,�3u%���;9H!�t#lh`�B}~��(Ia�%j��(���AG�=T���/�)���{G��{#��7+�f��	8]2�3��7^�˱�1%�x|�I�ĝ �\K�uFxŀY��}��U�-��x���q�"@�`�"��%�F6A��`A%���I ����'�,���Й�&� �E��AI��	w���t�"�����3vt"��
��o�W��en���m��Af`\f�E��Z��C�?��]��{T�*B����\�2����Q�~��Wd�.���5C赚���v����Ԓ�/e]�f �w� kQ�u@ϚF�^�_�]k�ް��u�fb.Sr���6R9���%1~d��{�����M��z�ݗ3k�[ =�яޯ<e)Ǯ@��f945�+��=S}����*�g�y���=+;�ͱ�x�z됾$���'��"���_��"���x�YR���uV��D ��4?	��e���H>:bѧ2�� �9g��Η=\��c�o=��������ei�;c~č*��s�ruS�VP�.w5��Q҆)��O����ѺA��kֱ�9$�(�
ˎV?�!�6����7i�Ih�T�B��-)��;љ_���-��B<��2���ɻd�~�Y�a*�r���k�DWc�5�7:�`K�58v�J7��+}� �2JL����id+dRG+?�1�9�3���s+���f�e�9�Fk$���nu&F��j�. �걯z��[T�2іƇA�%�(��H�qҕ!rUΩ>���m�f+%%<����� �|G{`�������$�U?�;��������qZ��J�����9G�I�Y��1��hV��18�7�W/����+sWq��(<۔��Eͭ�3��GG���B��bklH�^��-&��_����I�
�P/v�Տ߄D�m�Ch����̇�D���T+�W�H:~�!��K�;�D+�
���1!<o aQ�M��>����#��mn-����bl��<�������U�VuE�ӧ�)� �\(T1���J��N����ã�ă�s�>m��O�`���q���tv���u�lW�ݱ��m�ϫ�Z<MMm�\ ��Jټ�B��6,�u9c9��7�à�g[wN����ʸX���&:���R]��-׬DoAɩQfW�WQ�n��{���fr͖�O�'���$�f��-��E�"q���O5;;��]gs|F1��P��GeL*�gfl��;j����+~2�}�`� �zP�q%j�]8�-�O���^M�}�D�L#v6�P�=G��iP����g�cB䱄#MzH�Mr��[�q�T��3���}`=���B�?K��>��i�	0��$�(��Pm#1��p=��\�����ͨ7�5����h+�5�F�Ie��)�]�b�� T�H�^\]7���o��;��l�r����!��������P	X�!^�҇i�.���8�,3�{�5*��w��ō�'!2+s��)��Ew*��2�|��5�\g_h*.�3� �[B>��G�,������*����r��2Q����LD>��|�Z2S�}R�3���]^�����A?z]n.Hفa�^���V�������!�������>�f���#����'�^�d�t
(���2*������@��0S]@���(t6�xq�@�����O�Q�0ڟd
7U�GxOX�+�N)�p�xݼ^�%�K��0J9zs��i�V�O��'�Qh긃��Ԁ~$L��k��Ĺ]��<KF�������xz���&@��������v<W������D�t~>���.�e~{���A�_��=%����>�~ȸ�`��!P]��YVf��gmZheIRE�YG�9��ဖ,���b	�ܣ����Ʉ4�A]��4@��	��Z��-���3����#UD�z�k����cC��[a��m,f�Ikڕ8�"��{%����xϔ�X*�����Q�]H�&���\$���a���Ԋ�P�܊��P]H�G��@4Њ\&aA�gHy-Z����<��Xg͋��¥��LZ����PR�ޢ���`�?:�����?6m�Vq���O��M���	㖱��i:�̹{-#���pwJ��y����!���K;�껠{�Lv�K�a/��\��Ŧ�VSM��`Oo�eq���S+mC�]^� �%�W�v�5P����--��V�������i-�:d�V!,d���G����Ox\����b��20�yNnj���a�n0H&>�`�٥j85<�1?5�E,�n��B�G�w��Q_������e�>��E�c8m?�_}�z��"t*�~��댌j�Z|� 47�ś��,�X�����fe�\��)��$R�=�G���C���D4�8Ո%be���L�mדd1���ٰ�}�y��M�<(�a��n/���3�.k�D�<&Id�p/�i.<Y����Rw-I�Z��D~��J�ߏ:�2R�?��Dn��j@P^���)�n�?�� j���F�\Ł^����"��Q�eoV��ʒЁ�z�� �H��C�Y�b�9�f���T�͛c1��Us�-j֮3���V���p����)*G�x����A�7�@tYJ_2�>��Dd ;��X|���Y�yCuK����_���\��r,&�C��7��s2k�Z��N���ǽ�rn�j�Ӡp=kl��A����r
�)�/kU�������l���%	O��"h�NZS}8��K%���q� �Oz1~*K��#�f���� ��0f�d�TovqԷ��~Ci�Ю��*���O7�}��w�Z�G����E|/��*�8���Xʪ�a��yb�+��b���̥j���15v	���e����F�rur�#~[�C��U��	T�V�O�X�XXF�q���q�1C>�i	��0B#~S����Gˑ�3�L��&vb&*�K}��?o_�eU7���,�iӝ7H�=g�Y.}W냧n������7�=����{�Oh���ܹ>/׹��K6lh]�����U�i�oX�uY9�9G�W2XZ�D�b���{+XSU��偛/��:i�00o��	#,Sǳ��P`���Ș��<6˭>]z��;��F2�)��r��Mu-f<8�Qz�K`���|:�j����F��涅�f+�u�QW|���ͪ����%�T���`+�H.G��=��Z��S���ꋢ���	j�,��곆#���0t�g�2�:��Q�b�UU(l̀���f�c4H�A��Ѱ�y;2 :�0w��-7�5�K��3s�1�Ny]���� �����B6��/�3��d��/���&:Q����!C!�\g��S,f��_`:3yb�Il��5�_�ˁ����"��'�X�E��Y�Im6��_�[� ���qeڼ�Y9�*nޟ�ж�5�4)=S��s��<���7\� ���2PT
^����0�o�ݠN��v�Ao�����V��ϴO�C�a��̺��MJ.t��
�gtF�5��>Hn��3��&��
��tY	�� '
����)9��ߪ��u�/=�+�@��'�ry_�	�nN��^;��P�j�oo��iJ˪���G�����Tp�M�]���_L]��o	��W0�^9��Y8��>U$�b�& ���ȂN8��jRؚ!B��҅�ɫL4`�������6ȧ��(a!�\��ZF$��um��d����,�(��^ �l��G U�W�=�f���g�I�X�	���Q��t�\~����}І�Z3ujm�(��d�Bu���w��^?��*����R�R��;�=U`�xއ���د�.r�|ދ|Ǒ�x����L�;�H���k�%��"��/*���&w��?�;Kؿ`�����J��(`2��>Km��:��p�O���|��)G^҆=�b�ԗ��u�Q~�ɥ8=~���Y�b)�� v�m\J�o����Ղ��L�B�w�U1�8�u-�[ <N�����z��54�=g_p�����7��%���Sd�|��0&X�X�����2rG���b��Cg#���Z{��{�9� �R�}| �M�`�(�Q�QsO���������B�H����vZղ%����U�+8���vq�]Y����jx�oF(V/z���kQ�B ���Uh�|�4S�N�?��dk��w���Q)�wyDZ�z�-��s�I|h:3�`%
�T{ ]��՚���w���[�ÿ3����=o86��E\�,�rж�ч��Dߞ>�� ��Q8ʿ,Tt0@�`�\S$�B7�h�A�6�û��Vw�qb4��Ճ���ZB�>I���Ѩybա��V�8�Is5��}u\���uر�|`1��"S��c묊$f��i=�U=�:�#y�\�	w�%�2)���nG��V�T��N�7��P:yg3��`��	�B�S𵲗჎/ovy������X!����t��Kz�Y~pE�
q� M�K���O��=lnɺȝ���b�����}�J��N���;���'��2�P�㠬�����ˊbM�g��g���c��y�����r��㳤r^<�o�~?;B��s�8U�딧�ԌG�B��*!B���H�
���tH�I.:����GQ|�~l���?؊JiO����?�� ���Y���a����O��t���+��a���pF��nGٖ�
�d�Tܨ�	x~7�rm��˿�R�(� \o	�4Y@ ���[���9��<�r���1k2~Zb��i�={ESL��f�=��7&c㲋����97_��^UMY������I�;�i�[�c�%��ܞ[~���Ј�~V���D��G���~�n~���L��ኍ|gH^���诺�g��Le�5����y]noͶݭi�*�ȭ�OE���w�lҲ��+�y�¯���E�Ǹ̹�SkQ�ú�VxG���$2j���*���oP4��G�f~��cK�D��X�>.Q!�۪h*AG@d�$�L/�(i�n�u]� ���8�3)����_x�|������_��1�-k&�C�Ƚ��#��Yu�$�>|�*z�x7�qӣLd}��w�s"B�dKRB��y�"��y{��Fm�r�BMK��Ì��%��M��k�j�3�����+����Q���	P7��H,�����GޢZ�-WG�d�#�r5H载��9[�pJ���m�Z-d��f�0G[�d�1�0��'M�#u�M��gى�|�L!���Lil�Ū7�i��Ŗ�1�Re(rA6$���`/��Vpxw�P�@oD��j�A��I������_�!�d�7���F�������hK�LOn�Hڵ^�V/��c� �}^�q�W=����E��nY��զ�VmƁ�d��r��v�r	���Kғ�wRK���g�A��'?������7l �T=+�г��x�Bw�κ��x���_ʮ�&u�E�&��l����_0�,$۟47?�]b��CX̑��_$h���L�J�"mp���+o�V�A�~��=���z?�oR�P��Y��i��*��½m����m���@��`��+ �����W?���%vY�~^���Ce��e�ƅ�xL�W��$���>�ڠ�޻��N�t�,�����qObyT�a4��t�3.�Kl]U��xK�� +Om^	�-i5t
�'u�����Q���Һ��̌4v�*d��^82Pb���pL�F�%W�f{��x@����U_���<���{8/I���-��LK���"44Ъ��k	k��}���5�x��f���w�u�|>�џ�L�iA�DXj/���·���lmGE��p�V'�n��/�K���T	F��s�h[����QC
����R�!.F(�o�e�|Q&0�	M�4к��S��b��E
�)Z� ��]����='~@s�t��M�O��� ģ#[��zN�AL_�ڕ�,yHvp���o�དྷ�ή[�x�@y������
�F|]s��W���!�bY�!s�&#�bUj��hy�!C,�J��!V�$�݂�0�����˹��A_ٯ�\9X�>v4`�:�+I<�Q����tQ��2��WH��CO3�f�����Lr$��Jdx�aI絢^&`�
�?%K׈��£;���j�7k.w���U� v��k��iQ@����$�L�3Gxv2ԙ
\�[?�9J�~)�4����+NR�bz�e���ַ�A�������D�H"{!a�&;i��q��1),�x{L�'�2�j)��9y�ձ��u��X�|]v�!��Ü�	:z��<������oE+�%0W>f�{����jV�1��~���H��XԂlo�,�u�wU��ȶ5Y~2 B���C�TX�9KU}��+eC��i5S��<N�(�K'�"�꙾�&�J�qL�.^"TAٿP\��r�/�����1ƭE,-�ax⌷��+�+ګ0/�$i���ʮ�Qa""�k�[@��Vg���rN:�%�T�D�!���M#R�`�QW����(��r>���٥M�A��z0�{���u�4�؅<j���~ �N*����
��͐��Q�1��K�o02�";B����6���{���✊{އ��=���p� ����V5˚����0�[_����CyU�St	w��3u �4�Q�p1����i�bƖ*v�����ԏ�M�E�}Lv|*v�{�W���5#z�d�KZ@n�BpQs��ߪ�W��vPl�<��&^4�LA�2ϥ��oN�Y�+����G��x��{�O��������%?�J�G:�Z����#c��U2�@�w47#�-VJ��F�x˄��g��iR<w>^H?�O\�����D�T!��/���K�!G��)�t��'��P6�� D��D`Q�����<�%�O(�[Y�ѩ�����p�G(���e/�������/����YZB��|?�^$ v+��u�2�l5*�h��_m�W��0���c�R�ey�q��
%�B(^�Ǜ �\^5}v�* �.�*��F�X�7�q��`��� f��j�r0��fY#��ie��#�V�}u�-u~�+֩�f�ʀ��ؒ_��wU\�~O�U+0�4�%�~k,���	��Q#��Q��݁+oG������=���xi�7SV�ZӢ���
K���G��L��NGOsq�?�U�1ϕj��c~g�ed,��
6�>d���0{@����N��\cz-��^�
�����j�=�1����HH�z՗u+��ԩg},��q�uP��Bi�]��0eڱ����_ƹ�)@���9'�����A�ߍprw���9A��z�bW8��lm[�yQ��;z�%���U�>���o��֠��v�2c�B���i�V2}е�Rs�m���UN�P,�����v�֏����l���n#�H����0;��?1^�gy:쟥Rrk��p��a��.\L!�Uc7B�
%������8��J�y��G�.�,w0����E�W���53.�iy��>5�V٭.�Z��{���n�-�<hm��
���ʋȎǶڕ�no+څ���� @oտ�M�N�]E|rmfi/c�H)���S�!$�_'f��X½A�x�&��(���y��0r�듧�+@%�78#���8~bĴM��P��|��jݐC������ޓW���ɪ�=U�(�v2$�Xg���������X\���Pj���ɕ� �~)���"|$�G�b9�����/�+�=�	����C��|?����J��Z���RD?$�y�d�G�P�V��@���aU7�sk��Y��~�	$��k���@Ss�s$ה�^�AB�T���c�5,�c3�΃Mƍ#
ы��fN�]��L�n��x�����ER%���_`�N��A��a�x=���R�j|�
�\J������=����&+*�i�H�2R�����f�H�ґ��?[�������Юp� �J���6����{��E�Z/e���H����������>w}�j�3��6�WRd'�FY��^/-����>fd�?P?�r84��k��!��G_i�G^���0C���Q�w���^�˄?ƍ��%
�|�;X���K�!��K��F]+`�Vl�=��e�ud��X@!�|���rb5���Q*Pw���f���IR?��&�T��ZCe�"���8�Kd��&���!Ll�Ao���T�
���J/������d�Z��h��~'^+�r@�ЁCK�.�".��U^��	Ԡd��'����K���Z�$�ma�S$,�׏�>Տ���r?b)x,�Т�w���L��3���I��/9I��C�x&E�F�n�~+
�692{(��E` &7�xH�乂�=�a%����F'S;u��g��|.y6�
ur��7��.���E������V^�� �����fM�5H9�E%*j�U>���DGn6~���t�l��~-��k����,�fTK�G��B�Lo�30�K&|W��j3��^��HY D�K�8v��x�P��A.�ANC�S��%4W�~����tT���Z��V��H�sw�;��>��n�R��.��\�	�*a/���ts�s�KA��H�b����L�a�̫N\cX�Vʫ��a�
g�c\X��]>s�pN���gcٌ�S�<W/v�Q�Rk�(�^]�+����.��sV̊)%QS��طq�/�/�����A!=����	��0C���G�-���C�)D"�#/��M:#��
:���կ[|���{M:��Z`wﹶ����z,?��z�2����ѫ��ox�O΅a-��t��]C�Aw�Y��ԗ�w���QK����������0n�hm�N��h��\�ra��XM ۏp͝���'7��g���������0���ރ�edo���6yXƼ7��%2)�P��	H�ޔ5h%��D��JP3���#�<���^�s�q#E�
�	,Oc�X���,Ծ
L�E 24S	9;\��d͖#�o�7�=��5��T���b�) ��:���ґK���-����4/dDͤ#R�]�G���k�A:��~���"�p��Ʒ�|��ݣPH��@p~�9�)!�	9���ܬ��T�IQv)�~G�`&�olB��5�­T��c�$K�kC+ g}"��`��4��G�`��2n��N\��� [n2�wl�p_ty�b�ؽ q��#���qqN8+�J�ؾ���X�4,��/aƛ����*8���"2bL�]�ė�Gdcg��y.�7�ظ�Ӡ�x���FM��U,$3|t��DYO��8�{�5��P|���_[�%Xw��I )1���\�R��s`�	���K�F�ٶy�s���PZ�^����^��1`y�	�c��)�%n^�C�$I܎@�Y�ײ?\�T~4�~���E��cg�/���+3Ѵ^��uz4�Zǐ��z_�n\�Qmi,v
��qǩ��9ޯ]H=��d�F]�X��~%���T	kL��tO��-B B��qbH���^����N��eP/تi{�eګW��G.��`�i5&�m�V�}�w��[3����*��L�:*��x�K��nI��CA�y$H�7U'�Ŗڈ�e��3E��S<����t��ΰ:���b��������4�T3���.���9�/*d�t?�c�������Ķ�tNc�vǪ��LM��n���xp�JyGD�$Zvar\��x+�݋�%�t�6!Jo��3�{�dE�&�8�X�1�lQE�%-�P����7������� ��)]�Ӣ����]�}3g�\��$TA��0�"���z��dr ���$����H��%ڀ� N-�"�)�B�"��{ėv֨�2�����[N�5��Z��2 ���L�w�U'CKY�w� 70�t�)�A�y��y&�4�J��ɬ���+_p��9�߉��8U:�Vsf��{�uP�"�`�3t9إ����/\r�)��$�
�XL��UW0��Y�8H�={>�Q��6��|2��0K��e��8+	�$7�	���s@u�� ��)e�5���mKEu0Zc5� 2�6�V���8Fz��,�`�XA&���I�v��π�P���z�� ���#�b�i"���yؙ5�>�����/	�.�7R��J���0jd�-=��c�5�q�%��.�5�B�[��������Y�#�/�iD;�%Fk���Y�D($({�v+�؞W���"$[��NhC��`o�i ���5����v`ӊ��ܥ��Cj��}�8�$X��� "�R*���11��:��ǒ陬�)-���M�(&r�Qx�G?��'��]��ڱ��y�:�X�^�V��P$��}-�F��i�X;u�j�w��S]6�0���-T1�I��E�}9lUv
�]�~pUN0j�����9����ぴ����vي��;tq�gm ^�u���r:('�,�k��|کy\n!�MǸ}f�'��h���<�	�o%bh�#�zk׍�"5����_S��S�!�[6l���S#+�/��4r ������t/��K8��M��g
mU�?*v���.=d�`�� �pP���o�����[�r�+�<k�ػ��ޮ�[w�z[�sS`�%�`����%֯���۷O�\��#u<!;,	���wPy��5�V�<I��g��V~�Y��y�&�>t<�8ѹ�(+��O�?�N/��(��4x�����-������d�����¥W^�GZ�����<1����|d~��rn���.�"�=\>���_��A��P�`a둪��5eG`&~��n��&щ�6�ӠHbb{C�Ь�Ę6[��4�{�z���M)��G\�g��,�ű8Vg%��u�L�]�vÃ����;�#J$-�̓�k!�*�{�mܨ ���^3
�r���<��iɢyߌq�N1����	�U�kM��h<���V�.Z. 3{.�ۿcH&��@B���15�&��Q=�3�u���/���Em���&�c�s��Et�S��b�#�ˍ�^О�9<���r�T�o�4�)�����4��K����ܢ������߳~O�p1y j��\��o����C?�|C1s�������҅rĞ��a5O��3���& �I�٭�l֥�\�TESEQ�^+>�_�\d�B�ވ����1cW� ��:�hPn#0������\������ 	W��q�~���o�I)�"	�>�z- �ͻN�]�Bs-e;t�����i=�Z����Ŀ��:\��B����9��=<#�7ou��ͪ�{�9��.X�+3o>D��P���6Ӧ?�������k�DC&JQ��)�,��ڠ��v������9���&�f�d���r������3 ��,�ȥ�3'T�s������v"���Z�Е�����A�?�ĽO
�K���> ��@�u�c%�a�v����4��$.�`�J�j��܃�,�T���ۛM�Z��?9��7�Er�Q\F�@�&$X��m�$�B�A�ӹ�|��h��C�W`��B��ba��l���}~�2N���gѵ���xa�%���x:��Щ� Ї��R%��q?���e�*d]̳i1z�<��ތDؠu�rf,�o���<�a6z�Ȅ�C[�?�Ro4�<k9�����|�T�K��W�r�R��9A�����w�Xn�>�� �r�.���<=������v�cK#���J�)'3�����o��ht�vy�Ne"��4�so�"�=���C��p�e@�R77��9֌7kA��1vY�"q��r v#yQ=�����4��H�
]&�_�牒h���C��b�y@^U�*�@>�9�I��,�G�6����F���8�vV�	q���=��0��NF�)�o�3��"�Ͼ��yy�ݏ��F/%ȩOf�O��\O?���j(�9F�K4.��z����!� �4�.��eg�?.��l�]#���Ģͬ�'��3��~Q�%�Ι1L���q�f��S�9��e&���tc�DM���Qp-��2����J3�>�.�>ȥL�D��if=A.������j!��yAsͭ��p�v�h>YN�3(�\ِ�af�}�4;��R��cq^M�_xd^�S�Ԋ@!	ڤ �'��������S�Jو�h��*�� ��g�_;�;qU���H�S3���+�(nY�Z�
�;d90-Қ+��ޥ�^��M�=6w֩��ֺ/0)
��SH#�e��l�@��B*0�>�+S�v�
ڝW���n�ˋH��Ikq9Ͽ:'t9�ӡ&�+����-���x}=�,`��KBbfY�9�E�
�hֹ��犞��i��x�wK$j} ��-�0�m@��ֆ)D��[l��C^�/�^G��&����>L��yJE2Y+�x�*@��y�b`����_*����l>a�i��`P� <�z���^��}���Aq��v���л~I}�į3A��җ�m@S�)�Y2��Su'���+nv������*k��gA[ٙ_j��Sא�����^���+�h�L�Vu_tA���{��rIe��FډEɈY	��,>�i�ތ��R�>� ���3o*��^?au��?�\���P��Y�j م��@D�5�*�e�������[��P�Ⱦ�Љ�\*%�#08#�h�U�E�K,�W�4 o��|*�nm�B�0�Ʒ�&g����͏9��w��<��_$/��bbD�Y�ޗ�	bYJ���á�	��s:�DۛD'.��C1z1�/��"H�ɞo��G����>`·_8J�>M!X��1���#'�����*i^��}���������4�A�&�g��>(��A �5s�jq����^�+o���|��μ�}��|\Kw_y�R9	?���`��pn/��u��vq�� ����*��.��7�8/���\����M8H����<,�0��k�%:Vǋ���1?!�B��H���?*k�$�8�%�28����A�?3'��j��OJ�I^JTY��������Yq>6b��y�3�K��xΟ���Hj�	��Mp��ڼ����(���(|��Fψr����!D�~��M8��z�u�e���9���1�����`# ��J 7|�mo��t�m!���B����<`�K�-�,qx�B��������h�H��r���:���YQB�~�)�h>tً�,���]��Ұ���e�޹笫@�%;kf�춴H��}���4,���b�n���?i���_��R8�)���<Y�f���ʑA�,���M�aM���a��O������ ,�!����&9	,�����bY" �H:@����xVQ�0y�����]NB>a����]h�;�tUq��i��ɇ������U��ɧ�l�YՖ����pg��_Qĭ-%Do���,�%��+Ϲ����zt�ԡY�[ܵm3e�~Ak��+d�E�W;c�SM���j�`ة��Dט�0B�%0[�����2}� [{(�ŤM��U.6E*Az|MAh�<j�^�Է�=���FB�ymZU���Z�H���,�B~kC�	�)����A��])�:�)�:Wk��ز���k#��y0Ԃ4��)"��E��ɼ�V�2I�g&U/�/�s�W�Kw�0��=�Y�&�jo��b}8�NvL�v�-��v)3���YS.?��V�5�563�#%�w� #��%X9�Sjlm�8A�;.� ��!s$yDI@�/��d�ZTt?�|oh�~�IG��v��DE�E6�"�JI�֜[�m���㙧����#��OR �-�4���]л	7+�c,����_ٳG�M��x�>BD��n˱�8	b	D>�C��	q~c#h��p�*m�M���gL�����>�";��P%�6!'�����ǉ�BJ>�Y%<���TY�Cr�]HP\�T�&���[��w';��JQ�NU>.�{�Bp��wDw�}i�䁠S��76���s�ۆ�����Jl����UboQt�\9��=�*�Z�!\I� Td�����2�f��V���N�0�=%�l����m�Xn�c}�t��h?�S��\��[S4�o*�!Y��cΡ���'#�L�	�a�`�8�M*�g!�n������b�Dtd	hM����m�w#$B#�}[a�\PJ�J��J��l�|�6"��Uс��ز���!I�C[���Qt�(��c��t���N�g�U8�t�~u�=��ة��x��;v�6 ��~��^x#���{ ����G��,Yn�ky��	Ġ�x_��̈́����j���w,"�]���&5߫��gl�ߥ�8PQ`w	C��퐷�h+���Kn�ۃ'��ĥ	�~�nMe�k�\!Y;۝PZ{x/�-n4�;�;����2��Ǌt�҉����\mBq*v��ݞ���6��I�w��'��tڹz���5���f@��%)ن�w�3 �\�9���';�	���b�$  ���L��d_��p*�Y�M��ҠC����i<�3P�8��\���.����rE�ff�1TTn��k����S���I�v��Oi�C1���_�������{"Z���Յ+
�o���0y7E'�_H ^ݔ� �W3�]>�E�|D����Ց��+C�	�IJ	�x���DN�����LK�M��wa ������6u�7硂h��( ���_�K)�5p�*yB��Nk��%%�[aƅ�[(����)�t���Ӗѐ7?����G`sw�wg�H�8k�E9�nn��$��0����	71��'v�]"��*��zH����r��@�T.Χ���K1\�g0�/r�bvH����k�h�?�賿`�΃5m{�=W��`�CZf���7����#;�e���v"��#�vlF@�BPtt�����A�? �E�Ba\	��٨�(Ϗ�{�$��ۨ��X��v~!�.k-y˖�T
�6���Ѝ��7��.�\[)s[y,b�AS�=��"f_�Mhɖ��&L�(�tԭl�&t��̂`}�ۢ�]�I�*�l%5d��h�Ko;�(����1���*Xyts�Iɞ&6���n��Ɠ�~��0�NPW%�a ܚ�̡e�X	�.X��,|��I$cj*��j�����՚�T��F��/����p�H*;<�+T5,0\7�$���qM$�e�JcgS�Ջ��X�L	��>�B�mw%0$f�1J+�Gar�� U`A$�6nt$;����2��;U�����D"B����/h�"��vI	C��}B�����e��FCK��<_�F�x��`5�]�r0��ꝋQh��J��q�o�Q}�~���5�jvH��V��w��Cޮo����п�U:��xz�L�L�Q�{=��e����}+!���8X*&�i5Xf�i�<X�Lx?3�dP�>`�v�U�y�N����3��/�MpT�D���?
�Y��0V�lN�W�y��Cn6y�T(�����]��%�k�?�GU�#�{!��u����[ȥ����ș������b� be� Xe*�K �$����k�NM�ygI@:@����� �u �m�o���[���3H�^ᖻ�B�JJ�u�@W�9"�t6��(N�2�v;)z��]�6��"C2�����B]T#m�A q<�L ��tG�1:Ѹ�sDYI����X��ǝ�t%�;�T'Ɖ�˘ W]4u8�{%a��^Ȟc�'lL�q��iex`� ��اk�'�킑%��yO�N�Bp��ސ�]�����U)� _��_C���X�K�q��`�fM�����K�j��Ck�ؔP��}Y��=I:ɞQ���y�V�0��u�a�x5��>�L�ӭΩ\a���|��>o߲Μ���e����G?���cJb.,��mMAř����:Z�[���7�*�"%8k_���6ݡ�H�t4�������,���u�=]y�E�*�a�q��iWߨ�p�k�d��v��`j��5��9�,|��%*��j���}\�؞��	�1�{���>P[�S�ޭXWXKM�  X�8���6Bbie���&�=:�kp�o'��r�u�D�t��w�}Rǚ�!n\),�r5T�1ըp�Xݺp�p�r��6Ⱐ�&��DpNk��[�Ꜹ�_C=��$��'F��fs����9�]b����m#���+	5��tWw�E��hhv+d2s-�C�t�fd"�z/t��DTՂ�1:%d���Za^�`=�Ň��)J���u�J�
��鲂N���'�r��4�BYkZ�W��8q�W�
����m��1�I؛jG1jM�h�cY���������l�G��䆈��G����o1%�����!�N��7��/'�n	~U�;W���(K���R�͗�z1r���o֘�.ȷ��n^o�Z����g��մ�	R�����C���v�+�jq곸R�+�.�Y�U0NP'�뀕��/�τA��jQ�mА%�`6�X�)��s.��0��b�4;"J�S�/��,�M��n���8�	�ɵ�C+���tY]|,��JzkB8C�Z|9;i�
s(�,���wy��^�v�(�B�4�+����Óُ!����iZ��3�ϲΠG���#��˘�{��u���&3w�ggb���G)�}M�yT	!pY,�}�U��+��<}c�$A��Ѥ�_���M�t������4��,�kT��o��=����\;��9˅y�
E�	Rs� *c�(�d�sXO��W�i
Y�N�c^[�-�Q���]D���6�1+O��"����6]��*�" ��.��buYam1%*C�pR���֒��� 5�9�� ���En58�_����ۣ^��>8W!V�SԈ4���F���l���S�W?|�1Hb�Vكه0Z�I��J79.�xá��^^n��|4��%�	Ġ]�=�m%����°g�g4a�����G���Ņ|�	0�U�p.�1~�T��nQ��ˊ�/�.u�jh�>(�FK�x�*���>p�Z��W��0���1-�j���֢�a)_��zº§��G�	�m��� ��� ��d�7Y�5�y �`�IRE_�/���Ƞ7���&�;���d�I��P���rX�؀S�4v���Zˡ��wZ$s���m����w4�L1o��c`���A�^�k����|j0�l�r��W8����"����Z1,	������.�X�:壯g���+k�;}��$RQ�.@���� ���(�)�xej�i��)�A<;8]�^|��9�:��pn��=�~�a����Y��K���q4��M[�BxCm�i������p����"]��������H٩�B_׉�mY��4`_T
�|<�o��A�Uń?@�&|�Dß�<%0�� Rt�k�>�����V�7'2�.�^�R�u���O��׋��S�0|'ϡ�߈����7�;��%"M���12����o4߹�����>:p6˗���p	��&��W�Y���hg�aF���ՅZ�W��yA��gL��[9O�������ܲ[{[��2�Y퍲(��K!W��x`����k����x)����oh��W��I��F�k���U����c�/QH�������5�J��&}�UQ�6w�T��t��wY��9ȅ��0,�l�!����6q(�Tw�i.�#��k	��݉j��)�hYEg��w�Ԝ�|o!�BuE*VS�`��t���ª3�\�e;n�8���,J}^���&��U_�m���̭��J���$f�
��$��w�nx�� f͕�ࢮU���b+0�_WJ���EU��~1%��7����xKd��O�6�f���|l%@{�B������`Wʑ8�OX_#���-�ʉ1�(���;��������P���l��V�G���#,X�܌����� &}c�y���~��4�^�]�s�KH2��X����+qz��-lP0]\-}�F� 5~�)���Hk�.�v�|�9g&���]����y�~����{׋szfA��+k�?֧����I���F{��/%����(�\]�9�Ъ=���%��\�s?Ũ#2��cEAO�.`z]$J#᨝�����$�������d2dm�k+	D�F� [��bW
U+ GHI;s��g�_��v��Z�ɬ��}�I���r0��'X���*�v6�ȪYZ����+#*�O��+��{��F��5��w;*����7��[����T<fT�x�C.�4-y#L�vO�����T��0Z��h�b�3R ��KnӪ
k�DX��杻Xi2��[R��6��s#����T&/�c\v�k y2��^��}f�����ʒ�FߎLX��6���~X̹��;J����gpH���~���wǰU;j^�R���t{88�o��ij�{��i�F'f,}��?m�I�ҵ����J܊h'�:iV����\ؔHA0S$y���l�LO!��iԸ���d��,���V����b�8��z�w��Uv|J1�x�͉�̕�����nXH*�r���_ǔ����1A��0������'��#���J�����U�az1	P�����ڻQ�����kM]�����M��Y�g��H�(�#�r'��l�׍����{�T�3�uCy�KZ��n�Ljv�e�д?�F2��~5߻_�ˊu@�i*�>,����#��
�X�n��̆ V�e���%�~�(�Ϛ'�Dd'�~Z#�\��TE��[,���D�Ko~�-��pMW@�q��ɥʋ�E=�}���c����g�(^��?��!±ю�ģ�fϖ6mPv΂�oG�������j�7���'X�z8�G�����idޘ�i��&�Ѹ[�A#6�y�V�Ul�����s�����Hq�v\U����N�u�8+,��Y����&:u�So`� 7�ȶv�:����_;�L�3���_�(�l�	�rL������p<��]#Yw߷�Lo��0u�2��6��������afE�:p��㵊���}��8Eʍ_��2�!ZN�n�<��]l�WI`o��F���{iĻ���f
*Gr��������D���AJ8�'��6�qA�*t;�l6_��wᥨ�`��Bk��Ք�9d��c8g��x��<<�Dpgx(�q`-cf����~�����F_��/"{�Q�\~.1��RR�z��kY-h�{��A�Dͼ�˂���x��Ⱦ�V%l�?^XϦ�k�l+�|�O�A��X}��m�w#���F�z�� ���zkJp��6���>����&���/*�D�F ����F��"`����Y�W����T!<k����� �C�%�b��va�e��r g�5��n�vը()�y~��<�� U8���o ���ӳ���On��;KfgK�; w�S�ֺ��iò��#�)�Ɉ�׸��T���Q#���Z7N���Du`�rC�+X9T�m/���'��i��n��)�:3uD![��0k�JSb�+B�5�ğ�Sv��} In@�h�W�=$qp�#����e��.]!�X0b(��������%���q1|;%�FWms�L��~}�hׅ䈤Sp��]ճo�Z�'(�1�z��C�x���9Z`������܀}���v(��7�&�#��
�ܫ�?��2�sC��ɨ�E�P\�r��/Ҹ�Q&̵�C��_��T��|VLq.�e��EY�^3�J�����钢p��F3n	XɘT:�:����: �eaЧ����n�'�oJ�Xcз`)�j؄)��"�|I�MH��C:�1�pX���ĸ�#e����|�Lv���l�1��ಜb��bsE���5��F��D������,�k�aA�fڪB� L��3��*����$j�0��S/�V>�dmi��7�M�i�?Ķ'St�J�ocWyk�_~Fk��^0�6wJY󥞻0����9���	�8����6:0ׂ���ҙ�q�?ϫ��C�K���R�C��r�
L�xŞR,��<��i[�����ڿ�ppp4�#�zpKq��Tg�6�!�3�iӾ��]��L*��[�(�˟x2w:Vvr�P3���jG�*|
R	f-{n	�p�2d!ܖx]=?��h_d��RUыc��ǔ��$fv�`n@�󕃂'�����T�Ӈ�(�+���~�c[����;�����P��L�۶�����|v�߻je����AEW�(���mF^��u%�rb�;Y+�{x��!;ZY�[?����=�dBi���+�n���s�0�N򘨨l���pO8'�Ӄj�?--.
�rO���)��s��0
[	G=���e,���s������%�k���-���	��Ƿ:����Ax@h�lV�K.���ӐZ��8s# �6�8�z�>��֔�u|{������H��o���;{��]ʭmrgB�f�G����J���^���8��I�HQ�]c���&a���������o^-R� 1�h��E��5�<M�p�o�����}^A�����GT�0�<!y�����C���^ݺd��ԂW7Rza�Qі#��Ҵ3��A���W!!�!��X���>&\���W[tt��t�i����x{�b����ךO����~l��d��� aN�qk4�A��k��0E�M[Y����o#��f��.�K�(A�P�m���Ck���b�@��
!"���Y�zx�f��]�Ɗ�Y\D����_����F��v���&��w-]+U�4A��c{�4�����&��b����~U2+:5�ēp�x� �EJ����P�4�"�ӨѨ���M���T����C���D�V�s��p!˭��鎚�`vE��R;)��3��[u	OV������k�����f3��䓯@!o�g7_��={3c��w�%� ��a�	�vc
lM��F�^��֐�n��t>�v}�Ђ�9�_��h���>�hh桻�u)�t)�q,
舚�A*��v���	8 �T䞝2�x$�`�=��6C�s��aE2ko9�'sI����:��]��[ma�����?mF�6*��{��m�(���*� �AI42�Z�u�ķ�xU��xW;��vi�UW"����)�o�LR�x@�(�}4���CX�`,*���'[�[�CL�x�Pv��n�h�J�84�e�	w2�� ��`���Ēm��l���͆�5W��D-S(��m��V�G������I�c�� �Nn�L	{v�%��4e�������DnkJR��	[lD�r\�![wo�|i��Ꝛ"�6Z�V.��*�܀9# ��xCFFW�D1��"b��rF�"[���|I����q�qs��k4�����ꄇ�w͞X���ZBR�RI�fzG�����/3�K9�c"0[����ۣ�c�᠂��۴7�N��������(�W�yL�b�B�)�7Au�S�.z-2�\Z~�۽
�.5��$ޝv�R��q�-�h� �b�|�5Iõ5�x����]�sQ�*�F�.�T�E�ს�<'�hh�mv-!G@4��+wM>�~��=�?%�r��Z�Ly�3*��hf���:.���j�VH�/�(%,�g)��9�=l�-���;�yc-�TIR���A}�9��D��v�$;�<ج�L�6����/_�W�v�˸�O-[��%��_�Ra4}��'dV�d%��D�p�5<�������1#f�f. �ΜJ�T� �� �I�����B�J�p��=������g����]�z������"r�,b5jj��{>;A�v�en�CԼ733Nҳb�V�_[�"�&M%����v����К͡g�w�Fe`>�<*DR��'�������>��Iz���pJ1���P=��!!��0�E���}�y�����ѱ���af%ɵ�TA�%V���[n��P"�y� �����J*����5�B�y����\�(l_39��)�<���DY�4EV=�ԫ���F"d9���4��.�pz�r�� ��y},�H�a�)�o�S5����9���z������w�	���	A���X�%��B"�<�-�:�ln��� ��Zۋ���B_
f�M(�K$�[�*��c���	����o��z�H&�S*0Jk�<t��1��7i&J������B6T&2�}����S�!E�/˒��n�n/T���x:5U�� �H��I{b%��1MRvܜpvR�8��fj�.� 1h�N'�:�3�[�~s��2��-*��FN%��jԝ��T�Y�W�
>�4�����������(m�ƺ���9���y�@<�i��\�U`^&@�~��[��c\K�$�R��KD��u���W;'*�$�V�~*�M���[�
�C	����J��[c��p�W�n�a�%�݄��J�	�B�1����I�Ó%u�d5�=`� F�:bN�(Fd�K���@/aϒɘ������]��Z���ˈm6�����@1�=����:vLȖ{8Nv)+����7�U�j]J��ͷV���y��\�BNb������Ro�=E���;r]K9R�Z�!�;��$�N��1d"S��O�I�Gj��PO���$�����g�p���{�|r��<����R���}k�\b�AZD0����jio�b\]�����U�<��MT�W���On�2^�ԸpS�M�����0�$�����@F�wS�KT��ݚ�l�P=u}<O���3��kr=��N���纆�P�o�<��G\�:��Sn��(πӐ٨���p����L
�V�����fs{�������I)��=�R��2�
T�Q�:N=�ϠR~$������S�K<�/�N��q}˛��1ɡ.L�k/I�)����9_��1a��qaE��m�(��#bc��nqWNIc B�L���D>.&f�s|_�ϔ]�(��I�E�������L�������Vn��ây�=j�p��mZ~ ��?&� Fr���_�vc�&��%���J}9 �T��m���.��4��ث����C��6�D��HC+�XDZE�b�G�(�������g�*2ZN4f�ெ��[U�J���8&�i-���|��`>zOϒP~���۶E$/�}���hY�bU�e�HwL=P�@�k�	�̕TD��H�m�~���� �}%�Mȥ��5Z)��c�0,�E��M���9�C�5������t,�W����q �뵛��rP�����4�|�W� �������z$PU�p��R�6x��O����]$-�d�=}�q�)�Z![ eYvd�����i�>����P��/���i�z�%�|?�z�l�`Qe�l��3���+����A0ᷬ��_��N�ɘv<��B��[��~;b�^�Qxo�x'�-y9"D&m����J6.$P�4^Ę'3HAo/+�[i;5޴} ���ߠ��/�����$�t�㖪a�7�FQbK������7"ݙ)'m~��sze��ۣ0*^��n��V/�.�)��:f��~��r��mB��q��ˀ��u�T��A(Ǌ����?5٨&���n�4'����p>��,���v��x����l�N����?V37n���r>_���*�� 9�J�xe�
R}�j5�ޮ#�܂$�=!:!E��k�����q�c�����g��̓����n�T��I�Pl<fjnFF8X�4���RY�$a�.��<S+���&����i��WW�<���U���ux_�L�-�U�s������V�p��8���L�)Ėנ �����e�+{��2�s< ��U�9����b�7�	���R]���j��<Ql��&+�� ��
Q�O��GE!���c2�Հ�i�GbW�~e��~`%�LR��'�`ԟ��aً��W���:Y�J+� ��A����T���(�/���c�~$����Ի�sط�Ty���qz(�z��vVtu����F��z�/orw6���.�Y"_¯N
s���+�.}���ҏ^�?0?��-�wd�#u�	tQ�X8�Qu�:;��嫴~����ƋrIۈ�������r��{��k�;�-�,Ė9X���:+rё���RE����pH���'�G��2 ��@AQ؊oŐC�������j� 6'j�&�v�ԥښ�eY�Lv
�ʺ��ԑ= �byN�
��}�\|v>{@�Q;�\̶GN�Q���5,��B�����	I������@��'^�Z����"���^�]�ˢ��|�I��J�91��dZ��S^�[��߼m8��Q��� 8&���ʱ�����Rꅡ�`q'h��x%��]���l�K�.Dk�;��SQهv�%�K�v{[��,���+"�S�I��<������rC�,�s\�f�^~�Jc�n?ZS"
��p4�k��ӽ	+��׼d���+��CS'z�P���a�����Nݪ��-O��e�U�����;uo�b�	���n=�(f>�j��e�m~e��?I@�Ϡ:Xc��mQD$��^e_�&��?^FŸ���8'�a�����a_
qEm.rr����^>.(���ݴ��m.���Mm9`�ڷš1�����Ȁ�_�,T�{���j_�Ȗ�_#Q��0k���E@p5J��9�f������VJEuR'��o� �a ��\ۑ��8�-oW�i_���ǥ��)�9B�q��,�xǶ�0�Ҏ���]��ː5��hYS��K�����7�9q�O�b��T�x�>=�C�/i�v+���qYA�6z�����S]ŁH²^/�� �Gp�����-s�zH��`XJVk����!���4 �:`�2I�xR'S<}T�"��&��#2�;�m�l�f�G\�����{�7'��)��Q�>��Z�B>� W=ؙWl]��Ӑ?/��<��%�@��z�E<A���[�3�x�ȁ�s�@cW��y��#M��N%�s�����a�6�]9�5tD��A�o1Ê��"��~[9�Q���W���zU�` �3��������\�9�5��y������c�U���FBpQ�v2��j�Y�Wy �p�/�+�^�ĳ���:_&}�V�J���"��0��b�&��������;]�!��{�aۇG�dK�X��Yn���q
���V����ܰ��p��h��[����bJDk%�Y Bc�SB2bҠ|e�����+�Ռ%�Wd#����x���� R,|A
5[�����^���J|�V(DL��q�8�e�Ў\^օCG�����/'�o\�Ս�9`��0J�W��>H>�ZT�#�W��FY�[a��7o@	#3ѻ<Q�'��}��E�Lu���ո�yG�J��:NQ"+�7X��3&r����W]��5�1��7[�/�~ ��޾B���P C%b�����f �Ǵ
��n���,��1Y�Ros�B#��`q&�^�['��Zo�&e�=�f�P@��UH��Y�𤵍.?�@i����=7i�Ѣ+h/�<@.v���M#`Lµ���P���)���m߾:e��ͺ���s��j�^���	���Y�U��=��u�|����Q�y�_������z��u@^#W4<᲻t�Zz.Yz���/��3����[�~�#�d��|���f�n_+�k{�&��vajF5R�+q�NM�m@�H�R�d
�;�����%f�5���h	����x�R��@�L�Q\ng��.��'ZI�Mn���lパ@�Z������6���o�A��b7���߼�wc�w�bk�ߚ����)�dں���qhU%�!��q?��K��
5��2k��L�a����p��y�Z=�m���Tx[˩Ux�85HĝH�_�.�rf��
!��õ~�kŷ]����b̆O�q)���'�h"��2X+����j�5&+��A��Dq8Ϫ��8W`?�!eT������2fFQ���Ȳw�Z�h$n��'�mUp��NmDv:�T�q-ɼ6�h��;�Ø��Si�w0�w�c��
��ِ�1�����/��N�2�q��U�B-#�!�RbG�'H� �_LF4�y>h�Ӷ~�!�(D�yL>���a���aӧ�G���I	����-��fe�+���X�@9�K+i�<�И�z)����f]ٔ��*�T#qz�b.-!���9#�G�/������"�ڼ$9�ߞ$��i�]&9ħ��4(��N�"M͘�w�`���#����J��~�}�nY<)�Y�Rj\N�Q���+���z�[�Ӥ���j���E/.Jg�m^�鷇�-S�os<��܆���$*'1K�����a��uؼ���`�p�~�I��fr�,"/B݃�'h��n{,^����C�Ł~�x2���p  �M֣D@T��	F�[E���څND�����k��Ww}�2�	�3�F"G�΍E�'�tx�^R�,u&o�%���N�Npo�O.��K��&�0�e�J�s�B�j���Vl_���R�T�ΑϨ��g!��wGh��)n V�n�=�~|h����G���w�
4c�E�5s�XϽ�*���.�d�v�4}F ��iذ�~ &P�l���6K�����T�t�c�y<�l�{�=���J���ƚ�D���f~��-�Qs"K��IL�����U��*a��O�VB��e~�|k1��R�U�dА@t?�  �y#)��L��k�X��^�	���a�p��M���s����� �ʌ��)����Ç﷬�� O�O