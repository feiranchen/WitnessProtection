��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�EH7n�[pOY@������n*���/�%Y���y��:Q
m�=�iy�W��_�!_�� �@������u9s�V��M��ˠ �4|��0�f�~o����}����z�������
�學�'�A~��.��h**��n�r</�$X%[�����rWIx��:���a.����m�O4B���k��zg�O��(��gԿ����;��F�N&S0rU� �؇�7���k��TM�hrW���M@�c�"���kR�!~/>q�Q�����Z���4m�zq�l{�bRa۶���]E�17^7	Χ_6��8r������BFq�-sTe��'v)�����#�ف6��n�m�ό	��v<UyF���Ay*�	�q�����o�w�k�]� ��У�� �h�Cu��qB</������Ӽ1͛��6�{����F��'?oB¦3^3l�����{s�x�l�}����\H?�h���>]ڀ�&��&�_#���[A�� G�`1��JGC���&�,=�_jYi�x_+�>�d��.�^���]Pk\�a�H;�'�J�9����%�Gޓ�NM�!;	��Y�*�H�~�EX�m�� 2��TI��V�V�!�փ� �$���վ��?R3x�*6**���M&7`^�x�	�!���~6��T�Q����,=n>Q_��H����|���@,���<�Ęv�\N���r�S}���6� ��� ��^2������Ol>m�J�S�1�^���]vc�)�fk��}�ӳ�[䪒��˧T�я��t��h�:9�67��X�Y@�l91�o3M�/�
iA�Y���{ݩ)`����9ӫ��h�J����ޙ���d��UJk3�<�I�n�����X�%?�������nZ(
?h*Aɗ}|3r�j���`#���=)3����uO��.pU��W�^�O��QGCrn����3��]7>�}G\�� ����g�e��F�m��y�$��9m#Ij�$�"���{C-�=��(� v�o��`��S�̎�b�iլcR$	^��W�'��
��B؜
s��*k�Q�0�73=b@N�`�ܻ-�,]����QO&Z�_����8��g�@z�8mu(��� ���=�E1<bw�����;�F*bS�%�&�{�'�uX�����=Ԫ�Q�n~�T
��X�n���1���,�yّ���Zf)�@x�V�͹y������bS�A���s��-�O�ZᠠP�{�#�I��Θڼ$G:sY�����z��7�8��;����=oza׫@R>� 2Ls����U�@l�����������a�I���s����g��-��?���M�xL 3�c��#`��"c7z���&e�{O�so�PT��t0�a*��L�D�wyu���W;��O��ib�7�������/��J���-";Y� �7�����\B��y_�9�\���������<��>+ ���+�l"uTuV����'�<(�C'�k��ms��ϭҰ˰40�����i�R��u6���3v'����ۺi;8�Z2�j�Uk^%�7;˜�w:٭�=��V�f���Ղn��:o]z�O����h���4㌸����Ͻ�E@^�wN��ꬷ5��K?�AKQ]_��+d��4�9�*�1 ��(��7�R�B�A�FI5�&VQ� ��f��>F�wg���ū0_
E3��y���S@�[��P��r���M�(�D�-��꙲#� !�e������^=�yy��>ےWzYܫ������9絗�(���d��$B4�n�S�'ڈ��"U:7��Ƙ)�@j�"M�̯����A�f�97l���OeB�p�lrR��J[qG���NF�q�����>�t"�oʹ�/��˞�ֿ3� �d�\]\I	֭��dղ�E�{����h��2rRm�W]*)��Ko�� �#���g	A��:�Y�/q��.�$$�8���W���W�88ǍŝkaS��
��zA�z:[v��oקܪ�]��ع��n��\j<K���=��O!`o����� �u��v��<Y/�b��e-�H��^��]?e��d������X���ȮP*v��m��tv�xя����������u����q��Ѵ� ��Qy�%!�O;�H��Э��m2()ed�t,غtp�@���0���Fk}R�����+AHzE*���ٝc��N�3�~炍��w�f�:scN	Π���I�<���W��*Z���)�a���tˣ&N,��?�z������jח��Q
�Էљ%n���+��α�=^a~J��g*?ӻ����X��`�3T �E��9]Z�x�*猁��f���~����Ң�3{��{�{�Y�oc)\K7=��v��q���%ޑ�w�DS\>z�|���2a�-�{.�hd�d��߽����ާ{7�����G� %ґ�糞:�j���ߠ>)���5	���Q	x	_�>d��G���eDwF8>-�������k�_~�^w�^҅&4�<H^$ɡ�rK�W�4��^������P*��g0�+�I��tIrX��a%G.@����;י����P�I�t}02 ��5	����M<�m�7���LΖ�{��Gu#����&��>%ٽ��N�~��F�zz�|~
��Tg܈4�� �4�"_\�Lx �)~iu�k����re4���m�vH)F�4�����L�nUG,���u�����"<ar!N2&���1x��ZJ���Ғ�KT�b��C�l� ��ie���S��&`�/X�6�aAHl�NŸ�3�G��Rd�(,o"X�J?�7$a���`�M"n����~�.����)T�q:OLXV��W��P�@�-#4eNg��y�Ǻ����������Q@�dg��jd�ҧ�hȥ���$3�v��Ѽ�r�Q���ZN�uI:�J�R���Aoᳶ�Bi�G&��뢷
��Z~O�EMtCq�Y�V��V-%��`�x�'ǅ���N貟&ܶ�n�ܟ/�"��vC��
j��j�B��"M�VG� %���J.����������Ⲿ�_�n��K�A�ź�A�8��(�K0B]N����|@$�P��8Կ7��\�(��Q�JEz�Qv�;"�0{�p�B&~/�k�Ee%�mT���.�x��|㔏t�
�q|����a���-����8G�h��n*��d����=�8�u�� ����R��qj����֫�%��g_L�B+Hzξ�ރ�
͵����4�H�pxP���@�[*Y���� ������wT�{q+�ʇfq��K�ɬ��d�r�]��B�l�]���43���E��?�E7
!�Ž�;���u��L,
�����Z��ʇL���\��J�Ikxd�Fr۝�>�hĐvz�Q0$�"C��2s3�\�݇���;D���Nu����w��j0�j �̕��.>���
?�R<�)M�x04;Yõ�C�(�&!ޔ�
D��/�TG��e�K: ֌媿y�x<��7r��x�����6�9��"�W1GX�"Ȕ|�ԍ	|�8O!�`���O>_�?M.�1L����,+���b������4%`x�JiO������',-o0���l��i�E��s�i�Q�]�u���b�e�!�:a�h�fuQ,�z�V��C7`)����9w���_5Ɔ[��q�;.�ъ�9Kuΰ��۳�����p���19��4t�r��ay�;��DJƕ�T�٠�Y�"P�R8/.���c���]�]z�ѽ�?v��^&7�g���v�r�t"*��FL��ՒO�!��2�m� <��tћW��^���-`�+���.֮&�J�5����Vd�H\�3��z��X�x�z���H7:���ll.&1�4۴�쟼��l�m���ş��h�qxH[1�����v5��������mH�Cr���5�OPI���	�׭����@#�x(uu��s��[(Nq��b^\���%.�ě՟xr@dq�����>7���hG%��A�ǿ	�CO�q�Dz祳H�Qۚ��9V��-����I^�n�_!��Ѡ@V�gc�פT�e��Bj��#%�uZRS�䬰w%U` ���Ԯ�=�Bꀇ��5^���ifS@������b R� ��I6Q�p��"��w��r:_C�~��,�j*~-��6�s�� �W�%�)'��;|X�`-G�q����H���p��G�˝�bb�@3��sW* �ي���M�a��uqʛ ���'��v�99!6pp���:��I���Y���K��v���<ljY���ÁJ�iI�$�(Q�(i%PjN��4��ՠꭐ
ﵯt� �.C	G8i�����'y�䋩7�P6�6M��[7D�����Q���w�	���ne�b!܃R�5ߞ?�[З��7��Bs�,�tx��D����ʓCBDo$6ڜ�h�V#&�eo�ɺK���{$aO�/>WkA��p��$�й�b�9Z~1�Q�U_	L|�n�޷�ٔ��'��(z�멌ڸ?�U�a�����ʞt�f.��퉔%J'��x�L$�U�l���K��ޒ)�W$���.`0}� L�-�VW�ջ�)�6�=
F�_�x��[se�F�:W�8�U�G���3���_�w/��`�⚀D��xA�W�!�8���x@So��k:b�6�9�q$Z5�]�C�s���K{�'��0�]�L?T����ca����{Sc�_�AN��|���	j C,@�A(`ao�4Ʒ]��+�)�bbh"B�&��n}e�ڽ|uw:K5/]��r�4�`�)q{?8�,�Qi)���C\U�m	� �G�L�y�ޖP�D�0��{�����f�����eȆbCxHu�8�X�喾�&	�>!���>�A�tх�uU#)ƹI�	����e�|q��v���_���d5�*�\���m��ƂQ�N$<�@r�+m���Ǣ�S�$B��g���{����G�>f�P��Ųq��~'Ö�ۖ5P�n��O���g���ltA��Ւ�q������A|�[�uH�s��?@��
�8��v��mΧ��@S�����3Q��SpǈN(N�ZpS�������茴�(�1�I7��D������{s���8��;uAb���wp��
6��n�́B>�}%�k�������e@$q�q�G^@C@]m�g�eTq�6L�n���`= MX��!��/��&��'+M]>�&��$ZyYy�h��=A�Ů/}Cs#����ڲ@�+,��>,c�$!Q�gto�fn���V0���'�L��^ɑ �٨^.m�j%[�G�N�/�QU*=p�O`0�p�WSΖ����n3c�I��5�f��|��X��(�Ql7���i���1I��S$�jч|[6�Y�C�wc������k�tq�ZC�����V*J�h�@A{3�H�q���=�wgƂ�lc���;�J��<�t�@X��R���	�TzKKlhp��V���vZ��}@]0A��^F��%���2��y�uf-|���`��\���o�J�E`4����Tg�q���(�Kz�7�#���O�$[��;���R���<��BEժ�txT	cXʶхk]ܮَk�8���Q�����R��;�s�$���]�4�kH.�9D���:V�6��s�9��8�j.o���H���E��!4�Fݟ��Nn�1$��h�~m?���&j�A8��ZzGw�x+��$�u�ќ~e�I	���`e�{n��FF��qȂ ���R��ء�$]�[���wJ۱�T�E8a�;Vf�"���Ji�ay�^�:�=mL��Y����-�����b�Q8M�M�/�����g3 ��g���f*fa�1}#�!�XZ
nyi����߉��h�=~�O��^f^��'�#u�1���x��P�=&��ܶ�5;��)��v�3������"4SI���}���C;ق��y��%��/"� �f�d;�.�gK�G"/��"5Z*U�l9�:(�x�P��'�VҔ��I3e2���p8(&�/�����^��-\��8�C��r�PG@B�<�ӈ�Ґ����y&I�"�hzp`��5a'�0�8�|9!C��5�L|!<T��'��O�d�j^���GqL~�f�	6���8�W�J�0 -
�0�5�ݜN	��WN"t���F澠��gH�qj