��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�O��?A~'�1�{/t���O�&���۾^y�w�%������$@E4��Z 2�AһYV@�b�&) S=�N����r�r��{诀7�d��s}��t�,��Dl)w��EK$�	뱫���.��ǝ]'�[�C��I²��7����>�vҜ_L�ARI�P�kX�a;*���c�p�ғ�O	�1�2yoD;��a�@�v��]�̲��u뙱�Y`�}����-�2�}K�p6ͅ>*�� v��b=����ELlߝ��O����V/W�j��Z�y��ʙwf�c���eQ1�{ԟVR9�H ��9�bq�]��X��_�R(
�k:d�
�{��������%�����<����_�[~�q���n�a����*#�]h�[�+O���\�>!>��^�".Y�;���Q7Γ�yq���\�z������; ̻v�-���|'��������g0��]�gFw��hn�"�WW�OPV���a�2�O�&ƃ�yq���nA�i�����I����n���!�X#�z�0��р�������\�IP�`��5��^Y��=�|O�E�k-"��f������wN��lm3�����9O�����I4���E��{J����0b�\W`R��Mdy��)��T���
Y���,�x� 'G%�SI����7�vW��'Ю�����h}[:�E�QD>7,/����89�s����E+(瓤�al��P��
\��	���Є�"��[1���~Nqе�x�L���z�x��y:i۸�*S����������3/�d��ef�C��V�^a�%��%��kV�(@�����?6S�+5{�P.��m���i�Q�Ϧ0s/#���XG�kX�ԊD���d;�S
�c�=���k_����B_�|a���^�HQT�?����$�V q𨍃D�ۊ9 �b�q�)��SZ��>N����TԣTXt�A�,���d����aD�GA�wk������L������:C�N�^�@�S���9�:������nC�s��4�g���1��w�5BR�[�	�S6�ӳB]�	��M���WTJ��^�A��{�b���_`Gƀ`)Ѽ\���O�ȃ'�4<�6P�{q���8$�S$H4�y�
��A�GK�$
� �"M��2��pkdb��6�ڢ��^���33�<ɷ�U�2��>D)��ٷ몷G��D�l��?�߂H���j<���$H�~0�٤P�S�u�ppC�$g��&���Y�޶^By� |L�bE�u���p�<C���r���S��Ұ��A#�[+��ی68E/Q���l{ӕ̹��q�vg�8�Y	��aK�o=�7�3�	�'��k�:��`Q����)h����,Z��/fl `%�����M<��IӶ@o�7ݓJ��֐�w���пba���N�x)5�U���Mr}|KW��A��8<�s�0Z��K֠]����b���1р�0�Ca��H��]�4E ��������P*G�(�d%�qP�YTyTc6�Mۖ�Ƈ� H�%���t�����Ej�	��Vd��P[v]��������e��֤�׵լ^��%��`��[�{B| <���e-E�B'I=6�i]|8�P�����,X�F�F��������v����q�aU�#z�����b�7B���LQ��SdS����8��7wl�+*i���㾀�*N���@.�B_F\K�%�tJ:��%$7���[��Է��eh��D�͇�ү����j���
1�)r�_��6
_�4C���gN��7 �*���D�^�֍�7��2Q�#�I���(Y���G*�5��B�"��O��˪�S_��y{F�N+�����H��o�?�ݲJOz��#9epYr��h��ͺҰY�a<z6��z�Gܡ9��&���0��~߄I�,�~g�R��{��zv�6g�a�����$3k,���n �
���C�+�pA��e�M�����@�ܰkB���+��='�v6�����#Iޞ�Wj'�B�ƙ�=�U&/����$�$Y��z�+:3[�k�,�7��'}Z�s�!#TK��I�ؐ�gy�8��f Yr�-�K�8C^�v� ����OY��X��%U �<�O�9+qڎ�2֘���U։���̤�/�4���s[�1��d�W�T؟�9��$j/P�K�vLd�`gb�q�<�7�ZuB�B�S�s~��A�Ctm:��9����=��s�)��D1p�ݟey��w��?�HU�_�Q���A�8�Xg�n=3agV>�O�E1�ZZ�O�x�J��!�����OA� M�o3�>GU�`��;<F�7�[,����dK��q|�T�(NVY^�f��2 $R�yc��ط�%�9�	O�����@0�=�O�N�A��CsL%�F���Y.x�]�IAL�E�r�
v*�cg���'S�(Z��f��r�Br���՚4�-��#�/��UN��\�Z�5� ;�>�Z�ͫ Rs6~�B�`�����5�w�-��h�f�w�Q7�?t`��\�x��������ڄ�RAw������B9�Wl�h�v���Q���iy��,�YF�ז�X���Qk�<��Ԗ:�F��#+�K���M����'���j�\�p�Aezv��;70bSe��D��M�̢� ?K �Z`ۑ͢et@}$E��g���ɕ[��h�{x��9ʋQ�;�*��e����*�� ��Zj(+�0�xG�(.�Z 
�R\�+\��\�Ub3��~éP�I��h�WU��:,鱯N|�8������e�X��|��j��m_���KRK�T��
��s�%����j�w�mj�1O6��R��:*��Eˤ��õ,��*�{#9��ϣS�/����l�٨�����Df���EĬ���q�[!��{����J���#vj n���WռQ��;���rm�Q�Q�<ҭt�U�� �;��\�P�1>�$��LbU����N�p,Iz+'a}�����J>=�딺�|��k�E]��[�q�23i�����8�G��Pw��.�;�M��bO���yd���J���{�4~D%˾I�����v�D���B�C!y#0�^@SwZ䙨p�K�+� c����l�U���&d�HR��Q�@d�$w�\(I��	� �<�Z��S
\ئ蛹���{�#��h����>u��?�l�	i�oAQݣ���n�P�������5�>� D㧥ޫ���L�TJ�����Ǒ��c���FQ[pҐH���ţ;�0�Լ��K1��Nl?�(��CC���^�Nd�g�y6ˊ_	%��`��b���!nk0-d������L�3:G�����ꊧ����6�
�JX�؊yPI�7eO7z�e
�������{B�� �5#�j/���Xx�c�C��W�\4�~��
ހ��Z���M��D����K�Zj2K����?�t�y��a����Y��S��OwG�p���eW��Z��?�3�����C	a�����O�j	�s�h���SȗXjCVS�����=��m���a�@���A�E�I���7 T�2}�U����	����oB� M��7���������4\��k4�t-?H;[y�[���l��m�iI�y�YQM�<i�W@��
�r�s�?KH"H}�|.8�f܎��:��3_�n|�c!.�}�����"`K�f��k՟��`�/6�ѮIG<D��(e���0��E-�������ݘ��u��w��� ft���r��>�� � �D��|�v`��60t��8�9�JA_����tc�E	! �1�ò~�1�,��5�ل�P ��UM�=6�[CM+�b���Z�kD@��<�q��<w��ba�.�5���R��9@x�-u�XPoӹN��N�2�K&�z������Pp ft#R�i�ޟMxl�d5����O�׆�s�K�}�G\�8neC��Ȳ���Mz��h֞ú��=Ih|�BQZ2��-"�jT�����b�P��L�K�I*��oLmvxG��|R#�q��v
PWQ��<� #tQ���,[�N�,��ޮ��C��u^�Ah�x�_w�f���^EE0�w#,��BIu`U��4�d�Ց����K0�+��%WF�%���M����b�#)���2�v���H��&��z(y�O�%x��ȟ����C%�kw�p*��?�Pt�_��2cQ��&\��J�m�TO^��D��(;xD��Wܕ�n�S�-;�'�Q�U�Q�<��&=J9��'�R�2�@A�1Y�6�S� _e��C�'\a�{�j�*m��=�(��*���q���5,���O�K%d�C��m���r�f;�Yl����O��=|%k���Q�
9;kR[��D��v�iq[�=e����
�3��M�y��<�ɾ�w�������=���0^����;v�1�A��v�2ۅ/{;Y��]ySk|P\9K\��ٯ��(O*nU[{�������%�܂;V���aȘT����&��4��Y���N3a薡�V�P6(Kޤ`"�6�ش����%o
�'�qkrU�wE��ӗ������y�tN@��C�W��(�X4_ὀ$�t��Kt����r�	&�T��d)��~���\�L�Z���|���J4�Lw��J�ᱴ���C��l��\�HD0�P3h�&������n+{^坣�ߑ���bCD��'� ���_{��.� ��>�y�"�cNf��+��Tꞙݲ�x-a�!<??p�a�&��n��gچ�\�̨'6��[o`�t�-��_��3i�m۫���OQF,��]`�U!�1^O�Q� 2moK`�b�?�q�~t�朋:��p�r#c%S�[[ř<Kǐ��������k�)�)���;�T���a�S��K�2�8�x�I�F��0�SA������0$r���/(x��dз�N6%��:�}�D&��w^�.�Z�)���s�q�b�?���L���	�k��	#��f��f�
�G����5���e;vƙ���!�U�ӋE:a�xr���.���D���K�k��9�'딚��B=9O��$WGŔ�l=��m���rL�u#�mbĀs�k��s�q�o��`�A�|h���0'��KN���F�rZ���&ֶAzߞR�)�����q$a�C�;��qe�I;S�u
�*>}��{`P1�X��M����څDW�	�;�`�p��hǻ�o[i���qO�~_�l2��z�SkǆO��ߥ��aܶ�s��q�<L`
�^�i0�H�m�{E^����4��1�|�<SX$�.��C�kA8ՐX�ް�o.m8��e����~1_�+@$S�&f�?�<��[����=��U�1��a�ݣ��yA���nK����r���w�����<�3M���WJ_f���v\!��-�"���kڽ�э�eK��u_��rP]�ۏ;��v�:ԣ��
��Y3��;�ʗD�=��HMv�8��
H�\dX�;�hp4��JE��M+u:.GØܢ��B���)�N���.L�x.��7�7�{,�4��������	� ��%șs���OS�6�B�&#�M��3��8*CS���%\؛}'	;*��Ȳ2��hj!F=�S�-ӡw�D �������+ƣ���WN��P3�~�MK���SܽDo�&�X��#3�`H�'�t*X��u7�KKNV�	ˢ�>�Zʕ6o��|�^�`h��-󸵢`��@����i?Ԑ��� g]eQEG`Rxg��RLZjT_�/�d���d�i,F]�a$�WC.��q�(Z@P��)�۞�ȴI"�oV��	c$d�_��7p�.O�����Hvw��?E�`Z��:?�	7�5ۀRm�~b����}11{�G��P���&�<D���Y�� ��aL�bFnd���f���l�s��b��ܿ&�kp�4��ٱD�;�m���w�P�rf�%��5n8�������5�!u�B)Ė�Gu�{�8�W�J̜O���{;��!���ٱoʄ�:y�@�
t>B�i��'�7�G�@!v��q�Ⱶ�� g/"dI���E:�&���oS���q��q���5�U1y�ȏ��_�="a?߬]⵱})��T���g��@�D:�ӑ	MwV:I����pUmF�!S��풺Ƃ�gY��b����3��b ߓ�=J��?\�����	s��?�~Mx���e1WR���9 ��;�xJ�?�M�@�n�}ƫ*����Y�� �JN���S~��f��� �Sy�=���q��YT�0ͳ������e��� #�m�b�R�_¼yW� n ]R����ާ�X�/}�S.�?��L�0LV�������ڳ@���!��ϛ�na�Y0�n�%3�W�f�|���b��6s�:��X�{��;`��gApX��,-�.�7�FUI���Xŷ�s��u�E�ب�U%��D�,,xOZ��1��'�X�!Ф$r
�@�D�f���o�=���"�ù:;-cB�Ǵ2���W�u�a�	��{6�5�r^0cB[p"��;����N�M_�G(]Ǩ�#u6�H����z������zݍ����i�tC,�ֺ���)2m"u}Y��孶��M�� g��"�^O�V~�eO\g+4��%��3�w���(��T9�^����3$4j�[�|��z��]��@<�^>r�5��a����,���3��M�*Og���<�:�(v�_HH��T�们�zGhj��e*H�S��Fx`-�Er�g �IH�r
�����D���9������{��tq|>�Z��E0�Z<  �b]�g\3E�I�����A��-e&I �,f-X���bĐ�_
~���43�4(\��)ü�zi7�r�+�OosG;2�����vwJ�����y�%
��_���6 �,밑�S�������� {镌�"�G~�<����x8����Od�-̙s�c��Lh��69x����
�s^�ȕNs����̥�Ɯ�? �ޚ�R�	h)�o��,F�:	C\lC���*�qH9��t��_������(�:�z����X�
�r�`���M�$7jkְ�7�x�
�p=U�q��,�&j�^|s��dY���uM �g����5��ޞ�~o���\��pD�ݶ7c{Z[�0φ4n�T��C��Y��
}�����^��ˑ��ҫ,��#�}[-��N����Ʊ�1�]��cy�Miٓ\�8�U.Ǵ2��(6��#�/��X9�����&E8�s6Ǎljrr�A��.>Rwc��o�*)�}���)���+��9吗���L��f'�'+~SJQ���#s5���H�k<F�[Qk�Pe[Ε��� e�ִ���ty���  '�q&�ǿ+��F��2^.��h������b�	?�O����k0׽��AsN���C
@rl�&������<�ۿ9��GĿ���ߤL?9[�Z��6�tP�s�Q��C�=���Э%��Y{d�A/��tJv�~��zjt)idSl�L�k�z��0\q'�l1�igj\��W �wj��1\{��zH���z߉��i�%���	g�	��&�eg�!��6z��n�n9���5ۖ���I���s:���Mp���`N��=��f¯q��>��WU��b*�\�(��]�v'�}��$�g�0J��F{���7��� �F�Fx������LK�8K�Q�;�v�"��]�[�D=V����
^OSe>�#7��5�6��16�aP`A�6�O�pwS]G�9�5��8ֲ��q#.G����7/�>1��l���w����%�9$82
Kq*r�^?�T<0L͛�Sx<��D�S2 /�I_��fkG��`��]L�0����������w�ʅ>�-��)��qvA��J>��]h/�i1�����Z��p�C��&��+s�;F����XN�G�h6���/p���@����:��K�VC�me(��!
>Q�8��ֆ�qߎIψhE�y]�5�&�,b�{��G��g^�Ϧc���܁�U⭂�e<��.���ըC�\�G�2�x��v���7�D[�`N��fI��YHM���@��09p:As��~
���Z ��b�����sN��N�~����c���3u��sw[(��G�cR�rU�]��>i, 6�>0��a��JGd?�+	N}�xN�M��Kj����2�Kָ��c�M��
�+�=�-��B��g+���]����T���A�f�fJ.�Wpx9_���zN���Y���H ~=['����(p��؃*J�w�	����t�7���6<�p5��NJ]��W)�������\�r3U����Ɉ!A��S�cu��4M�ﹹ�.��ŀ�"�wʤK��Fߌ�d!*����lׇ�"����ȭ�����`��HgTZ[�P] <	��������$7��OLʯ�HV:"i0o�$�)��h@&���;�E/��!j��U���w1j�&�5r�"nd�*u�V��w�ܤ�0��W�F���~��Ѳ!����tk�N�WO�y[�`��R4��*���\�����_�WL���Zy��R~.�[c�Z�,C���l�6�Ax6�A7?�
�m��D�
,�4���0l]�8��h�+�ш�h�|�Tm����=3�V|L8Ve�a<&9���R*L������Ԉ�CDW� yI0��c$�e�*��ዬ��.x!8��IG�*>���HW�`�&�u�D����R���s��(�#��>��n/�1��j E�a��8f����ؕK֊*<�D��=��b�ry��P���SU�&���E������Ïp�:_7Nѝ�ޗ���j��l�JI-�{:/G��Zu��