��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q������5Ij@�fK��s�8�Pm;�̘���������RzF��c	�^K�[ߤ���p(�b��:��Ɯf����?1�gؖ�7W�uJEF$'l�q^l\wَf�ͩ[.��6��+�����3��
I���4>�h�|L���Λ0j��a���o'�������MH:b��E=�r
$�?�|>z������rbu�U'b�N�� �CueXȬ#DЙ��Vlm��@-�DɧW^R2�[:��`H(�ߜ��{K׽�n�.��c�,˴g��{y���U���0�*x
,e1C�W�O3
�Z�6N�v��1��z�fչ�[����f[������d�m�=��7�SIXHnV-���~�{��eR*"o�S!N�#���� ��L�ɔ�m�^Ň	s��K����yᝌ�A��������� �Za�63B�����{��7}w����#yN�f�D����{����n���� X��z낲�]{<&�_�Wb��Q�{|}g�X0C�[�B/;�уF�WŜ�����]�0�����@��3��@O0�]n@�Ѱ����
f��Mmh�
��eZ^��K:;�s�}����Lu��
��A�꜓U��Y��8B��f�2!�vA�7��_�]�w�Y�0{�p��)Q�T)���IAP���nD��&�jeX�s����G?F����OO �Hi�ӝ�p��W��;�.����:�:�G ���s�������`Ge#nu��Rk6�t�l#��dR�D!i/��t�$� �ϵ����_|%g�|�J�.C�ieb��H����ڸ/���B*nu�&����S���Y�E�����6d��P�'l�����v�9�2�jrg��\b�Iث�'e	m��zaH��6 C����j�-�y�)��EHn#�a��,!H��np�1DB���������%��W�$�λ�n���N�Ă�񩙪y0�^�w��-�%��X�k��j7-��1��@M#�-�}E_g�����K�m|]��8aq�?t�ba�7T���	];m��������$�2��^��X#�����A����$*l����,����v��F:\9��C[J�"
��L�{�x��7�G�� �����F_��E�K��p\U'�36�q�څJ"d�C.��ߌN���X�6��7���k�|P�߾sP5�n���4��L���H�j�j�I{t�喏��g,�/gh�#"|�D"�u<��1�%l���+M��+���k�����O\VE��8� ��D*�ts.#�ܻ���[�j���� k�_�����jc�$��s�r�Mn��*�ѽCgJ�>yk�|�=��P���}d��Eq3m��j�f����W�E]>lmhޔ�f�W��X0�hF=J��&%��C��"�c��N%|��CB�K/�x��W�q�)F���D�lk����6�˿����ܣ�P��s��82�E�7�GC}�H¤�<u��^��`j:��X��iN&e���;�4k4���H3��{Y��ǻi�I�]vq�L��U>�A�	TE��1b��
����C&��������b�Z� �͢,,�r²�iߦ����0!C��`;�.^��G1(�DZY<�6�������+�S'y}"���3���C-�:����2	B�m"�E�l�_N����N	�񇽝��3;/�P���I��.k��M?��t�m]�94�7�R�1�7����i�sf����^�(횩HV2k��6WT߯�� ��l<�OaI0����y�	�!�P4r����c^mg�� ���� ��h����O
�oe���[߮5 ���:����B���q�#_���E�L�_���YO���"ff���W�R>�R)F�*�Q�pZu�Q� �W;��Vسz`BOr��M���S7��4n���#,FA=J�
�D�}����x:�&Eᦎp��e^ AɆ�M�KC���VQ.`�	�1�Y-�47i�	%o�m�ج�9�K(lr�$�,N�wA�yе4ݛr����^ܜ�=D��� ������(=m��ybqR{�ze��;��*O��4��47t~�����
TO!�XU3�>4�ѕI2R��[{Ջѭ��4�]�CNF	x3�|XСN� ��$Dv�w�B��O��}�Q ��ZX�
FuC�n3�Zɥ�1�2�����I�X�'.x�@�MB���	�8H��g%,i�clª�4cS��	̀��Ӥ�Zo��|@;��3�4��q�SKZ��`��޶H���!���d����xi��6���L�%.DQ|o�Q��������o�;6�3�0�=w|α2m��.����b���v��3��7}�/�����P?����\�S2B+������Qtr�31�����jx�m����-�h푲�<�����^K���VE
U����(#^�{����|)k��Ǐh����l�Ro8��lSJ��y�TP��KMqN�Hhk�1��zk=�>�qC�0�c#"�E�8�s�IC"ܠ@��c���K�ڰ���.P֎%v�t�~�$�������gq��Ѻ���h��(����b��P(j'����,_hJ��j��f�w������sEKl������#T�1�,p\o~�|���^M�o��v�[�����?��� ���,V��]$��~�U�Q *����2���\�I1���ȸ������t�@��(�p�B�m�v#�=&�{��ny�"7�ZN-4��㗸� ���k<#U��7����ߤ8�v�cbu��`H~-w�����t�D��"YH�v��Yo��8��~��&�k�p�Ջ�HF���U�	:��"�%]�
w����n��>�lM����(ڟ(�[X�-��\�MM/ݓ��A��d�\��Y�E<�P��{�3UՏkgv�n�;��1��G�� �t�ԯ$27�\ל��~@��ʅ��X������q�����sir���[LZA�eNBGuVE;��s���]�r�������6�?G7F��q=F� � 3�)�[���9��ۨ���*��#JD��y�g�w�Sp��!�JLt�)��f_�V��/��00C����\Q�J�(����T_���4veh��H�)����W����h��&�g�A,a,W�!����вE
�lX���R�[-#|��Uc�J���E�do:嫒j�}�upL�Xt*"Ӂ�DZ��fg���oP��1��UaO��X��?.Y�a��n�+�m[������7Vm����]���p1���-I�˭�C��o��}�h���ð�0�̣ίa���/qF�HE��\��^�b���O�LTTC�lS�'Q]������;�T��j�������
�W��ۿ��B#��_k�7��ݫ���"O���s�M��8�eS�P��(�y:�����х��>'�*(WWEpR_:��w��\+�FF=�jx+T���42���:�E�����!V'�ktH[e�e����X^��ne�hu�zP�ӭ�Z$C�S�h�c7I�B%�����H�kz��re�S�<V֎�D��޶��.����auRy#fN�;s�ܷ�(^r�x�M��	�Z�+rf���(�PN5{�e� ��˺Q��:��{��!�-�r���zܮ�pj��õ2��9�]�-�%��d�NV��:��G^�]��"z�τ�����I���0��_���Y��OM�GY���j%8 ��º����T�V��g�[چ����H�@u;�y�H�<8{����Z���8�L6��	��eQ퀅"�(FU%d�(֥��C�yko��l��xN+^�b ��6��(W�T|>+T��|#e���z�mT�]�g73}��f�_�ͩ�e��x�8�5Bb�C�{�!�ե c����..5��E�I�R�p5��'@b���\�ǆe@�Y0�I`�6fv�hc�jG��1��t�v�G���]6��S��5(�j,�]�c��~�	N���u�;���9�P*D�¥��E��hGe*��8A�3C����Bf�O��c�Q��3q��Y���:V[,�x��E�3t��&�S}�rѲy
�B���cYz)?��,�{*i6��6�E���1���D	JiA�f�4�ΠSl�r@w���D�k��i�\\�{*%�m�e'�W]�5�責 ��+���(�,���r���d~�?��	&z��*��P�	�8��%t��۠r���މ��k�����F�KD�9"7�.d*hPQ)�v�hvw�a���1��Ztyb���Fz�>��O��҃�Ӓ(e]C6����/�ܝ�v�,��|��ޜ�h��b>GW���O��BBɹ�uY�4���I�J�_�o���K�|;e�/�^��N�(��"ϮR�r�Vuф*ӎs<�7��qv��e�p���2�1����Z[Bp�Ȏ4�X\E+�2�T�1��H㑾��*�5�?�^�{�ĩY�I��!��W�ܪU�Zc;|	���\�nEz��G��u@Ϛ��-ʼf�@{;,�&�U]8���E��,X�M��j?�ކ����+���x@��ř�y���@#���p=M�߼@�R�?�S=��'㰇��ep�������(⨷ѧ��{ƺu�،Q���='������Dw�w@\%:�al�Nk3>T�¥�t��S��� Fc2�ϛ4���Z|��^�=�������ߛ/c���*�VS&N"�D9R��q��V�� �VA:C1��[SrV�0�m���h]��i�za�|Ĭ!��}�"Cp���}~k�|��~��r�3E&9`�c|ISa��g��Z��'�2}f�h�g��Ŝ��'�Lqi,�}�A;Oyu��!2Ea��j�bwD��.��n��I{r�Jǃ14u�x��ۂʍ��CdQ���&�p��*��Bhad�$x��S*��Tp��x_�0��S:@��\�*��N���Iu��]z$)v��jB�7v��7�.y��k8"Y����R]���}Q�@'\�?]��A�楌ERzĀf��]��,�v��{�W]}PU�Uq�}N��Ǔ��pM?��fA����Jݢ�O��J���/G�"_�4���y�q9�P����,O�bx��iOc��s�O����E{�"!1�[��3�>U�7�3�$�
)�'��p�H��9-���+ѱU�4/��^ׁ1����G��i�i��6@$'Yq�ɯ�<��7��f�����~n�qe7�ս��U&���*8�2I�
����i8��|)2���|��Im���͑�igv5�)��WC�C>A�a!�g���f?�MU���y���ę�����	'��Zw̥��Yb�w�d��^�����VY��:�����G&��I��%�ϯ^��Ak��ߧ���PRO����jdu���O�F�Rb�I��ԛ�����Z9�|�ؑ�ް7T���Rd2�1��h����)����;{����v�«�z�=0�7,���|����\Y�����+������!q͒��Rgoܝ���hV�6r�D<�!��e���B�l�fQ-�P��>59.Iq�q��FlV|}��Nr���h��x�T�S��+XG���g��v	
��I�>���Vis�����sbN�
�H�	�R���z1�sf�rg�	x��[6�ٔ�ё4V[�B)�ƺ5������bh���m��^3V�1o��j��ZUf��e��U���-fՂ�
ht����@h(���/�TgU*X��Aېû���^A���e��6�'��E�����m����0��`ڒ�.���o�=q�v�=L,�x�/�3�A�G�:*3����F���3rb)�ɶ�81�P#�T�g��1�u����Bg�t��I���Q$ӕ)iQ����J�.�l�+"����c�:�AL�,_c6���L�bLP��_�s݃fJBTkI���s0�H]��*'�I2A�{rM)]��Q�j�BMp�0L��~�~�������z�[�H��̃�3�o
h> �ڈr/f���/S���.�=���7Z� �Б"imlV#��$���
�[�ڞ�R��]�:��Q�6s�ڹfCu8Xx�W�|�A�YM���@��A��BW?qDy<�^���0'��(��w�ў���	�v�v���W���6g@�g�3q�h�O��6�Ô���M?,ȯ���s`��%H�>�{��$���x�D���q�������	}��A�Ԃp�wUX/Җ2�چ$<�>�L6H�ܤ��%{��)Za�H��VVi{�yd��Ľo��c@㻹XI�ʁ�q��d#A�-�ɔYO3j:���ݜs���ì7Lv
��b��.�M�E���VĤ�J�M�`�o5�M9�Nm�n)u���-�m��Mώ�E�o�1�4w��UTn�������$�������ۍ��D�޿�(eN���|��J�27�X8���rC�h�5�E��Q��3=<=��	��6Bs�ޯ�#������}��[T����Z+:h�G5��e�X�"��@�-|��Cjy6���Q�Q�9cxX����70�J^����3U/t(�CW�"Q<�Z��a���t��A���*�9p4	�=�=�\��y��n!���h�w}j�Z�Wd��R|���-U9oW��Ԇ�v ��M�"�.��K�X�V"99�����42�>:d����_L��p���C>���+"w
�k�7�LK�jYpڙ�!�L�O�3��LǤ���:�43/U�c�[O��^{��
��$�5�z�9���gN�	&�������D�p�eG|SVZ#Aÿ6���H�^ܨ�O�\=��:F���ݸ���,�G�=��>1�~�G`�1]=���kx\�L�zA��C�|�v����j8�1I��e��C.F����w�Q'�9�O�O�R�G"0 H�۞�s��2A-����9K(#��� q���ট��X��w�^o��_����f���m�����Hou��&���Q�nt��b�(��B��#�43	�kL`y��U�����G�"���Eԣ��)��+���#R<~;euz{Li)~Ȉ̸>{Ty,W&�t�i�Y��o�Ҳ�">��
s�/�柃�yAww���$E!�?�ܪxvly�,��Ÿ�:�3&��F��̔���H��w��ҵ�q�(]�DF�;#��%s���Fh#]ز3������E���T��tj@ߨ,���aQ��IX@Y�_e!3UOɱY����C:~+�);ti���j,�rg���ĒV�Y�/aKk{�\X9\��w�$:c���J7{k��$��Gz ub �wA�=1��_D�N�)B�*�R�/3c��������$���vo�^�(G��������7���pqqJE뵺�
74}88��h)�R&B�g�7��.6Ǐ�l:�lN��U�)�E�GKP�t��z���XNz��(�V$�ԛ�z��O�Q@�~��'�����͗��F3�r��D�0g]�5��R�b8Uӹ$���N�Gk:R�Kut��R�!������}��&������\�O�I��_���r <PN�N#��%z����eE���b�i�S�.��x
��"�6�a��t�W�
}{^�9Y��<��5|l*�Y�_�Fn�a���G�"��{(ŏ%L�)4L���]�IdO�2����㪹�p��(�W  C�2Q[Ĉ��/��zH���n.�u��