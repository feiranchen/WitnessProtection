��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX� ��V��P�e�ϧ#��z�����J!�G1t__���/8�
�{9:vS�A�@�j�6�:�`��"��[J��G��6�8�D��~�/�Bl�gl�M�X�Y��G]�����mxK�z_9��[Ʌk!�DP��zqآ��Cj�}�ɺ��x3�t�3B>D�,4�S�&G���������y�ȽM��Q/�''e?'ڡX�þ��2��� +S�cN����Ġ�4 ��1�)ѕ���!8�Z�?��$�I�1
�+F�}H���E̚�o*��H�P�SC|�1��Go�������+I�|l�q2\!S�*�V��!�q''���-0����oj�Uo�l��V��|�;dQ���߿�̃k���Y5!���\r#�0�ך�ߴPT;6B[r�,��`�#�ȷ|�`k�tP���5|[+]�E��b+"ܿ���u�[�hl���\p,��}�����g��,~���JO,��	�N�Cn�H���2)7��x��H.�<������4�!k�M���tk���j� c$��-Tu�e�&ܾN�Ȉ��i�֦巉�N�6|\_��F�Շ��ù&��	��X���T��t.hjёs@��P�Qc�Jm�����Ǎ:���(':̟#V�,��F�*j7�Zfh6���wp�qb�y�cFԿ���?���|Ɂ��Ϻ9�.��R�آ@�>	��f)��yMP��6�g5�EFl�(_��;��8�(,GA-�&F���jF�=�` �H�b��f �u���[��*�R�h�k�.tʕ�fO��Ϩʨ�w�Y*�w�f�3�V)!Jå{/�vE�Y���P�	����^��c ą�ZUդ��*bh/�a��2*­�(������$��>��0/¶B�1����/�����c0���U�`�攄us�!��ˣ�E`�/��_��.�K��;��V��3��n-���YiY���@g���t$2*�6*v9�)��g����x���r =[�G"�;R���e�;l9@�J!r����5Q�) ��V))G֐�V$j��R�x;ꅸ!z�H6U!��_	�����'��\e�Ĕ;,�� �̐�'C����ɭ$��F�8���`����ymD���> 	���������f�8�%@/+�H]	���u�n�,�}}=�<ʃ�;��b��S�k�(k�g�\�<7��$L��1����6C�����4qLq��S���O����6��y`!^*�����t�om�Z��|��U6~ˋ���f[o)���Y��6'N����ʸ��3@It�1�=������xџ�0w�9�~OCN��p���̕���7q��1C�F��.��W�S��������A�a-2�;(���*�V_ж�c�N�9۩�A���땰Aʇ�#�d��/N���k�~��i�6�Ih��p�Ă��������#/���B����X�~`셐����z�����R�5<r7��&ì������,u�[�Z���afiHQ�l<-d����G��\r�y��h&�A=wcw2�%�+h����_�c� �(Ԭ��Y1�	8�xɶ�xAW�_��<�tC�4����e��/�ѧ�[�N����^ak�K\���'7��rw�T��IaV��vZ:y�O�� ���;x;e���C��3�e[
��6����|>��DAfEcx�\�sH4~�"��b���#K�ω/������������a�[vd����:����^��&�b�c�I�����^W�6̖����H���l�y�����ބ\6L]�A]�#��k�a���处�q���$��r��b,Fs5pBk�1�[[��?~��L~���	sE��y/O���i2��l>����݈�J1��}�~+��#=I�5�bϲ(�KJ���/���v�/�������d�m#���-��|g��/�#l���Ba*���^ٚ��!y���i&+�|I6�;6.-pn�Lb��&��kS�5�Z�eA�c��T���X��X6-�v�"�m)�::��~�0dیk��b ��h�IH���QH�s�L�ԃ�����2#�c��bl���R?�M���o�8b⳱>���AC��v}���V��B(7O.H�¾�2r	�o]R��f3f�㪪��K����JR�t������G���V�fꛗh�0˝K�]=���U�M�q��^P�(��n$/]�Ls=o&z��r+[�����'ӡ<��5���+5!ֳ{�}=�N�W*�Ñ�~������?�z��#jQ��Ԓ3)�r!;����!3��w�!c��3���6� @�ܑ������5k/˦Z�5���3��Hy��XAAySN���嚁�Ӎ�!2��������'�ѝ1�k���wü}���lG������e�䁻�Dd.�oK��=KR	�I�*�;�'��������vum�d��Q2�KцM_��w����V�f�`��o���&b�=_~@��s�9R�#�K�����
�U��^�a�� i6*��~��c�!{:�M5:��ް�Aŝ�?8�Tg����D:c'��@�(���z�$KX0vŃG�kdU���a)^�y�\:�C�����t�8B|/�{�|���y�>K�B���'�?4�O�^�=k\�qY�^)_'�N)<\r<��Y�~�������Ӆ��+CZ�+bi	Y ���?Z��� ,�rZ4&�?i�o��@����(��[%4�.�$��b�^	':r'U��&}��(?r�+�=���ܦ\,TUS6�,��l�ņS���4��u&쉧)���z�9�����)��[��f ۚ{��V��.8��ɋj6E:�G�_�:�5B�k������4�J���?.[s2�	�L��o<���4<aAɨ�%?�Z��=����"��+�mW/��C&�˂g��g�nKB��Lvq��xT��K��9�S@q�:�ؠΡ:x"���m��xZ��� S�Cb��*ѥ> 7�I2��zND�v��sp=��5��^���"Ih1�Y���С-SѓXD�!�Զ�� ZX��K�����F`��Y���%�y[�1������+s�0ѱ+���t����4hS�Aiލ%�Am �՞�Y���㨙��)��{�!�z�E~"�}�O�#�TrV+��W�g����m�~�6�;h��T��`6Um��JO���n��Q~�Si� 䓬����}\D_�RJ�k鶊�_��L�r�J^c����N��E��Zv�aԱ-�$݅���]���u��� �0փ��:�>���2c�36���J�Ȟ����.�6�2�!*��K�@��b3��V�{�/b!�}��'/"��nř�/�	�HU���j�7�,��w?¾�Ÿ�c��&���X�S>!���Eа�I�tK�x���xLL_2ك���֘���A�������6�.��T�I|�����̬�̙�p�	�%R���q��K����F*��z���\��Y�B����S
�WϹ���v�BISVA� fp��΍�9Ħ��=���E��~��O'�H:M'���`�������p�n`�hF�/�?�W:�f�Kb�(&v�QҀ�'iŎ��i��G����{�*�&��T�y���7L�a�H�>:?(A|/��Zs��JW�IJ�0�"��;w]��g���U6�E���~�����Q	�<�� �::���L0�@�t�z��Ғ}�7���a
9���9w�(����ّ�1�.�Xu���K�u�9���b�	a��i��������E�B��%��[:�|`�#���ǒ'�
��j�,��ŴX��X�	A����Ԃ��k3��� I��Z�H]!	*j���3ӿS�&�6�؇��EI����V uC�#�}�9��[;ȷ��=?�i�2N[��g��W6f���w�D��Bi�BwOt�np�8[�ׁt����L�R+���}���g�o\p9�D'P�|hyb�Z|�Q;�}��EEp��r��3(-|�5��b@�I�j�5'��>ΰۇb,R��Жwޚ��.�X��MäpeN�
MSkmc�2=�c�OP�yQ&~t� �L1����Uwn�o�2`1�[F��6Sھ����t�����.��_��nlE��%\���9�¸^�����}@�ec��cJ����QӍ�ԕ&��д�f��i��|��?�e�87P�/iV���yP\����$2aʑ1�Z��6Uy����u6UʦΥ�,�W���-�L��3�^D&CbbN���M���rE����!I�O��>��B�#4UG$o�֖ ܇�R�NN�li�Ti��ߴ�T��L;OO�R
����ɣpH��Ng'�Ι1�F2!:wUPY�Vg�$�[v+���Xyb�2�a��4��q{�Q��5��`2��fo�;Wq����G�`F�lp6#��@�܏�0X<�2�X���R�k�L^����A��58�?�^м��ZJ G��>�����ű��Uzq�ɤ�*r�2K{5�
���Mv��r�9,@��㋳�wø~$&[��I"�Co��xl6�(�'�yek���1ch៻����	 P�<���\���&gAj�:°�K,��5��GWh@�hCk�3" �H0�9pn�X%�9����!�	pS���$�.���8		�U����z�Y��M�&t4�s�N�3Z�,�M	�>���k�����G��[	$�$�221;���i<�|~R�`H����6����C��k(Oer^,��4`"%�c6��u@�c��[*�H|�͸Ɩ��v�h��c)�{���i;���`���<���-@����e�U���x{R��/kbS<�:�s��>�t$z?��0��(q�����"`��"���'���QZk-0���15��2�Y$�]�''�PN����8�����g�W� Ɣ����o�l���8�Ar0_@Ҷ�{#��H�:"`����7��7��V�7u���Z>)����HQ��{���lupL�m��y��H���bE�� �8��.�=�K��L��P��=���ۆn M�������Ӳ:e�}:ɒ���.Z4��_��v!�A�:����k����S��) ���:����n��y�d�e+T������I���)�̵~�k�����J~�\[Ӽ��0��/4����{ +:�Z��>��u(��	>�I��1���%��ۅ�'Ȯ� g�ϥ%y` �J\���"-��;��J��	�Ixy_Q�@�ꅙ���1
-&�������V�ݦ���G���]��aLU��s-y��il*s�'~�m��T�Zb��d�K^U�M��#���l��6�ip��XkO�wh�_�7��~1��/S��P�������5��E��GH}5�s��56Łg�L�k�j�Ï�|&�nYlj.-�C�&�j�&�q���1ɷ!�5�����dchi��l�1�$�g_�����!�O����f
Z>E�-�̯,�[�^��}Jr�ۖ���˄8ނ���p��
{[�9�4U4�v3�E;�H�,@D<����-����A������!Ã/�<�Ä���>�T�ro��)�/< �؟�M8�4�:�3��8|���` S�(��1A��\��$3�Lc�E[E�8��l���jydC���o���R�$�Z�J���FY�&���r.��E#���\9\��۵t���(r�,�E��aAۊ
)�F4t�Z�{�J��Gov�Z�q�}���{���Ք����	���`�+\�|��kʒ��Y�Z�t�Y��j�)�{�=��oϦ�Y�KǪ-N�ųf���L�d*8H�V�����{�DXO#�"l �BOܿ�Z���
�1�i3�7Fe��<�IɊ=iB�K���Xj�Z��Bd;+�xSV���[,]�E�9'o�(����B�vO�����T�#(���qLN�;���Η����C�P8	�q�;�z(�tDzN�>�%�1Zq��~�|#ű6���.��|�o�vT͡��V�	tl���2��؄��:�o�D����$�6M�/CؾL���ɱ Y����Q�q��R���@���5j
��Ph !�:X��~�?(v}�wN�q�6��]N�Ʋ
KI�zU��9�/��[��p�f�N�+�}�&z�Sc�~S^$�d���9y�7��Բ^<��r!�2	�X�aQ�F�S����1��+��g��o��������N,?�.�#����L}"�k�r����v������ܓ(ѓj�p����|�ރ6���6ݺ+µ��/��?�^���4�8%��=(�P��B'՘gK�����)�]����^HXaR���3�k�'�mn��.J�yalV�?M�n�Ḛ��d���:�����.2�u/���i��^j���C�:�o�-�גƿ���Q�0˿���X��M%U>G�?��\�#T<��O�u�������
oV�f�w!(-����d������G��� "���&۟a��y���D-�xsf�X�[�&aH�$�FZ����ֆ�g��u�\�9Ô�Ut�����:�K��:Yc�`'TO����t5��Z�x��6�2!�!%sV���Pg����+�|�P��l��q�O�`�fz~L�P!�y�g��z$�6~�^Z>����x�qЛ"��>He;*F� ��0��f ����Tn#M��vY�4Z���
�DX/#� �3�d��샡�������<3#���d番���ulwap��dG��^�a��ؾ���MS�1��s���������.�j��s�A�ϗ����3�!�v��@w��^���="��&fu%����N��"N�.<W��ʓK<ؕ���`�v�c�]n��{ѽ�*��fs��<k�f�?�gKNOh_߹p����L�C+1�1��Џc���$��J~3�ڶ�eF�|��W@LEܲ�o>��=G�q9g܇K����ɐ<K/�ct����IO- =k��\v�an!�ə�B:Q����>i֘ ����N_��^բ)m���Er������*p�<��3�J�[�T��=x��^�!�~�l���=?f�F�B�{y��;�3��[32{Ԅ�߽'2+�j���Cw�ڰ��zo�,�C��>Mj#z3�E#$Qh6c��HH������i#���HIA������"��x*_�5:����!I&g�u-&���,�Y\�S��&�_Д^��\����Tb-� �T���O��Q�<��e�D}>W�h׬X�%��̷��'����� d2����z���(�zP�}"?WY��7ì�kB�܄������b���_�	���O8��C����(�5?Y{��L��Ɩ���H�VJ�/�Q�-�N���*�Ej�J�m\�#�q�p��y�U���������B��A+�Tt8����FcΖS�8g��
�����1�ơ�|e�m�pk��44���0��t�%�Z�b�*�o�Z���8��k-g��Z�3gT�EDv��1�}d��Q �Ӌ2G>�*�{`�V�&�	�A3���eǥhP"׏�֡��+��Z\AX ��c�������͇��ﱹ��s\�7���![�8bF^�<&I�'�$pul��
9#%K���o��|w��I�C$8�" 
X�Pb�t{��w���_N>�>�!6�6"�&�z_X�0fM����]����\����A�+f�������<�6oTV��+�Ŀ��b�@�&K(�	a/z�خ�RC�~��1�����<=�g2Gvh3����n�/���?e4��iN��$��/S)Z�#�Vc_v���\CV�� �S��P�5`����n���p�<PV�}��n�P�p��J�v^���$�3�`5�c��&$�P�ni�B����?����сy^Ne{Ÿ^#[J�������J�i�(��Ip*p�s=�4e��r�!�oz��-)K"U*�ï��!�W��i�h���\�b����Kܮb#�u�YY$)9,�q���f?NHň�Z��{�q�̩/�F�#��y�VaK�7�	#�Ţ�����sR�l��_�ɮe8>�/&��׸7�1`�¤څS��JAi곩�W��ɸS���E�4E,l�?[��H�*-��Kvq��9b��� �$-�V&g
�\4T7P	���ֳy�͉�O(C�n��m��+�L7ǈ�N�����X���o;S�|����a����]ڬ��\T��]=�/Zʴ���l�����>@4y�5�)k�}��K��S�E����
^�v~���A6���]�Ӈ�>�x���V�~�֎��5g�{2�TW����Q���^�O�/�D��+��M�/)-�
\L%�H+rPf�'�؀�E��Y����=���.MOarr_��c
�je�M!t��o�*I�Zk����l�/������o*}������/�{�F}���R��W�,m�V��tē%�Q��!�Z$�8�*V3v�H�Ix����8����66��L_�c���XgH��=�����!ӻ�`4��%��45hk�����c���#yE��KH<�/fC�e��t�t4)O�P&;Q[���f-�j���i#߁���!|p��0e�-c�b�`m�uh���yTzW	�;ٚ���+���������8٭�zP����a��A�{�:�O_���	���:�NT1�����ڲ���Yλ��?��
SR�|���O���N,c�o�>9�
YC<M���w����Zw�;�7ر��lK(~x.����y��4���z��Sz_���Y��Z7ʅ�5�j�������`ָ�,���JL\mC�c�f�\�� L��8�il�,����V>�����G3Qw�V�I�	��.�$���j�䧗 )����Seg���L��$�4e�T�dm�y�8l�E/�8�6���]�}]
��S�Z��ҡ&+P�u���͠N�~Q����9�8�eĸ'2�&
��1xY�(5!ϳ	��sw���G ;iC�4p�җ�pv
��#d��]Mݩ~��(m���Ok�T��
�9[֎|���t�\f$!�;M%褞_o,�W�/!�Y�{H=�UJ��"Z��<:��;ܴڲ��v��%k��T���̖=3ώ�L}���C%��t��N�:���|��8p��fJC.�/M4L��ž���V�U,c�Y%��v��c��_vuBψߍ:�`̡��<\���Pa<Ey��I����(n��#���5���A������)(�@�㯶K��F�&) �rk�	�鎝l7�����!
_��	�93��,/�0�\�݉>��(�u�__[^ՠ��qJ9�o��������N@�`	ϹX7Q'ʸˇZ��}���<�ڪ=��x��A���^˳�xR�U�P�Ծhr��ٵqX܏l�\�"������$E���h���/�Z�[f��43�"Ώ�4��1�p������Q�O�ڡ�y�>��j7s>���z�������,`
�__��wY�ݰ]���!��5���Pv��wh
L�8��m��7龲�t|<� |F����O���՗��%ԗ���fN���`1����G�EW������
�.��?��#?��LKAYe݈j��άqs<�1j�Zj� �֙p�ꯟw��`��� Q�Xeg��M&�X�9�d�f~]�\��|��33`<;��k���˽�tp�k� �w��6��}�,����O&n0��Q����,S�C�Y����~H������W��n��9���� W	%Ѫ���+�����E�v�9��Ł_b)�i��iX�;��03	ৱ~�yF�����~�Wd��c��lW�Id���p(�x�W�qC���~W�N�ZTSR�b�;�v@�U� �mF_�P#��i2v>4�&m6u-�vx��w��_�Mm (� b����qG��j��K�\<6���:�4�7s��'���L&y�c3�Ӈ�R��b�+T1�m?����5'�q�{����1y�)H��С�����{D�
IY,�l7RΑ�0a[L�\
O��Y&�{�ƌ�[����S���0�~�T^|��jN�@��nF�59d�z&3��Z�,&�ђĘ�h��!vV�׺?��36v)���Pٚ�-9T��D"L���G����@[��S�i�Դ9|�t[�����d7��]t���!4}m<o�l�Q�u,d�%gW�]B!�(��-'gO���B�x�i}h���E���r��,A\1����T�Б�x|�+b��	7s�خ���O����|���V�YK� ��[v���ćd�瘘Ern6u��R�_�.��%%�^�~Z,�l��Ybo���;�Sj�"4'G���T��m#��מ`1�LdVO�*$*@�˖�Dm�"��hP++ �H��C�Z�c��&�+�V�3#ZuUym���qKK���}���k�Q�eg�z���n�aG4P	��nd�w=ZH`h�)q�y�x�9c��,��O���N��8����?C�������?�;��#���p�8ؾR�˾�ޛŪ[dt�y����[�71��=^�����p��i�JC.����-`(5��8`̱0��[�HX��ߜ��_�W�JWn�xڣzҥ��]=���a�c���AU1��U����W,Ř�#���L`��rK�4�]u"�N�w&7�;�0�z��)FχS2Q�=�$��A�X���|Ć�7��A���q�(
[�L�������g�M�� �8�bZ�'��#9ߝ� )Z�%��
�p���2QE�������A.��P���S���̀}���������ɍ}����*����~�^c����Wh"C;��~�����[y=�z���B��s��?�0q:ʅ�J��'��hF�F�(P��HZ�Y(՗"��k�0`<��z.\�B�pKp
 3(s�WM�~�}�c8忔�8��ǎ�����A��''�pgy��<��p����$���f�#=�p�JO3b�¨�0�j��D�3��<���t�r�?`��|<�ڃQ�E�����3^��y���s��N2Ҫ3�/ �j×N��v����4
���̐�s��v|�Ě�k�Zk���� ��a�ph�+I�6�O��Wv�'0��^��}��sL�, �}�#v�"�ޛ^����^_�/��rI/�Q�qq|��x�����jR|ϳ���ϴ���g��XX��ӑ!���?�(�Q���\(Y�2q>�\�:�-s�����Aw�d�^J�K�����@��|T���d�$�jd���U�l�kG��J|S�R���G�D%���8���*�֨����I�7M�{��{q~�������Hj�����7z����^'?N�Q�g�]Y�s�?�	U��W��t���w�����"3��9�UmB@���ᤘ��*RM�t����Zp�z�v�5�v0>�������FZ;"*I�ä�8�o	��\|F�Qn��jF{eHL�\�M$@�a '��͚`�OOGpd,�c�1v������6�2Տ���JRfU�CI�Rѧl#7�[�#ڦ��V�%jLVܚ��*�Cu��^%�@@1uP��$�b3ѷ��|0�
�o���K�vV�����szT,���D<8���ݖ��"(��=h��j-ce�n%�J0'���d�OƦ鉇�q&�+��'�U��ts7� ���n'=F�R�r�&�c�ʙ��j�{7٘(��}�k�W���4�́섲��_)Y��+�"� F�����2�bۊ& k��L��V��"�l�����F�3����C�6���O&Kg@�M��A�痳����) �F,�
�HR���kb�獠k2����}�-aΩ���Sr�[�W�:�N�r�.�5C;��VX�W��,��.r#ɠ���	��@��j~%��i��j�*u� 0�\I`�a:Vn�A���-8���=`��S�1|�����y�h9h/��S�֥z�l�N(��$]U��L@��E<�l)D�	��vS�'�LT+4;Z�iV���Hx�Qc��թ���im���� nB8�����\?��O��g�{*��c��?w`��(���ZQ�]K��qx�l4Hh�%q�:�L�Q�����cI���X��V�ۋ����p?�c2c��g�}�j#�&�3���~��3���A�h�ZN:�,������R�p�r��4_R�O��l��3_��#(9��|�?���G>��Z��7b�ףugpn��4Pt�jA�Z�y7���SB�<G^*�J��hW�������mlU
O�A���ᮎ��	8��%qj�����M����Y�H0����	1�Mg������H���!���6>Y6I�n, ]:B4�6B܈
f�(�:��>�Μ?�����略�2u���[���(�1)`bb?���Jᐔ�R+����NO�������.�KL����J6@��H�]���u���ȱxX����Ǯ��$��p�����J�y9�= ���(�/۞�9��6]]��'�����Ē,���Ξ��"��8�K�����)'�V�w����Z�2�mZ�p)��v_0�.�qf�Ôl]q(M�_*7?�_C�
��Qd�{>��
���B��!P�D�<��1�W���F�iC�����F�����@��<s:����)���J��y��K=�&|,��C��:���`��mFH_g؜�Q��+�/��\�4*ꘃ�x/�h�|��:�i�M��s;^�� �5���o�|͐06@GU���%֤S�͝.kt��������R��>>�����<���
R{�5�n�.O)�מđ!g��QR�_J�a��¥�O�;8==��`�w�`��0��靊B9C-���{��+�mI�i�ͼi^�?K�A'��"�\�Ƥ��]������0�6��
4�}~/=�h� o֘j���0�$�+��+q����ķ�����u�L�yx��վ�d
\k�h"��?n^�0`����`��SΞr�8�l����J��@N��sQ�(��?�F��S�n*���oܫw$�h>7EY���ko����*�ڷpoWX�0<F\e���G���sN�~���R�duD$�����T��@C��8��O?�q����I��B��lʍ[}x|��L"�u�W�P޴���-���V�I��|R�}:��7y��[ u��j����M 57!���f^�X�'��sx>p�"�-|/��}v����#�C{��?j�F���H=�xv��#)}�0bi�`��G�'�iS��鐮�c����>��-%����ɐ����OCx�e���m!7�o�o\D�-v���.�L޸H�(	"@��6��q�=x܌ل7��E�f���M^�,"�a`Q������-v�os�n4z(4b�$�s��<�@�v?W�i�(���Enδ�"����<.3����:~��G�؅Li�u�aUpK��e�K铒�2�`u�/�E1>�Fx�ㄌ�0μ[���-��y�$�@���)��?�A���R��Q( G��hLj	!�N�\�o+�
C���oK�o�)����q�ֻ��I;r��Aܙ aO�?�A��d���fRъ�땎��֮����
ª=5�����ͱ�0�ΣJiA���F3��\^L�M��J! vx�I�mn�^�giU�
%n۲��#�cwY���({f�A�8˜pwU��ёn\C��i~����}ԟ��0T{�Y9²�������&�JC������?�1����X�'t�?�{4�(�o�j@��t�0��w��C`����������5�h��F{��91��t�n�΅}��DXB`5�����|:B�4������b2� ު|�5�%Љ��b���ӹj��	v�����6-�;;Fg�\���v�!��%cX�3@��ː�	h��a���|4c���fT���@�s����7O�U�j32�P��Un~`�D͞97��Z+���E� ��Gd����JB�[�%��QÓ��Xa��o���U}b�U�c #.�Y�c5~���������<nX�u���KA�px`���x�1�pF�c�?�Vz�tǻUU����˄!O.x�����M�q� ŗt�U���+=�P]���H���K�:�ۨ2|	�?���u_�<��)W���4�?��1�,�#�P�ς:ϸi�v{ظv�9a�V-`�ax
��&O����d�?�C4���l�%`"�*�Y�5�n'��x���5�Y?�U�J��x��{@�c�7��سIAl�eMMx	C�ke����rD������.����n��eJ���_������I|gcA浬���E�`�o� �N쑭� cwL8�Vѧ��p?˯���7��OMFΈ\>#�I��ٹ��p���"���9�E� ������w.�_<�0Y�?R��2ⲐzV���CN�E�( �2@�M�BJ�ۓbl�=��@�No�׹�����Wx��Gfq��f"~r���M��Ѕ����r�(���a��J�Ȯas|����L%͌��2�g`X:U���\��'Bdd�����g��"]�Aw�!� �����AkQ��8�q4��t��i���?:l���r�r�P�-&$?�~��e'͚�Pҫ�@�Eu#�u���N�����s;��C�܃��д�N��-�|�����<�b|췋B���ݤ�MsQ�ѦO��WS�����bL�t��׿O6�~]���c�mX��j�p�|xwB-XH>q툷�T8|�9-��=�_�i�@��"r��fWl��k=����Hw�i��?ܺ'�1G�KKo"�A�Z<�J�T�\�޳�-�lHν�G�*��;7Ň`[[+��4RfX�ҕu}Xѯ�W���o�a� D��'�HFz\��v�-KV�_��"���0컿�h����';+��s�o�nf���\�f|�Ө`�N��G�'�[f�گ�f�P ���O�����n�<����e�C'�a3%��-z��^zњ ��~�)��#���*����ʚ��n"w����-�Z����¤u�D�cuiV���9����b���������aM�DP��z�h�j���W��H��H����0ǥc��v;2v��# ���[2�;Q���/��yÁ3�N��
ĵ5���;5_���� �3��!ԍ�]�LM���/ql���&��4lVW�Ğ?&�-�m\�(u�9�����HK���zi(�2.������owA�3�d�Y��ZB��3��6��b�����]�,����!�QT����%���;���U�?iN���0f�-�@�'����Lm*�p`�S�i�.q��=�b$�����0�^<AI5�-�Z\��1/UR��a�6m�h��.��5S܋y�\{K%��FR8���#�uS�Ei�u�߲�6{�%5@��N���E�݂�՟�������Lb��h.��\�m����*;P�b J}��Ok!���܉B�͡�:(+�.�Ϧ�Ş��E�c��&���t?�-��"�`ay�'_L���u������
�����׊#�?��ҿ�"��*eW��E�n��jz��E�iin0����}.әaO�ٴ(�Pn�����
��L���7�����P�ѫ^�v[M��qV���3�yU��(�@˙�1�Av�w�.���r߮ �����-�6��3=g�[(�!�FJ�ǏҮ���ߞ��F共wP= �0����>ה�eȶ�U��>Y�߭uF�B�w���  ���x6�~V'����}���|S]��f�b}tݜ�|,�l9B�?rF�|�8���/�s�����ʹuH6��ǘ�ƞ�����K��0��tx��o \gq�H���kv,+�E+�2��p���:P���.ADŨ���:���/�뤢{��Q{<�H���@C�ZUH��jmҲN��<l�{̮h��k_��L�wz�_��C��Ђ�RAX�R�C:� c�#�g��T[5��Q����2T�	M��jR� $c���Ԅ�{���1���h�K��r
���Y4�M'],%�F���IV�,����D�h�]�[������1�B����8�޷%��"w͂4��ѩ}�U��_x��L�3c��z���aT���ib>z��NXDI�_��E��V��ן|�¦x�Vim���U[�W�g̟,�TP�M $��'Y�NPe(�&m��Dowl_���6�f��C�����|a�:̗�RV0�	��:����3$�9>_�4�t�,�/v�W���s�����p���!���s�:�]���yh�W��/J"=>w)p0�\-='��_	,ొ,��oq-ǐV�;=bV5������f��N��������=�`~6���%�xˢ����o,	���SB�<��ѣ�,J��^�hd�z�s{�$7�P6��-Fl��C]mj���F�a)Wp{��ے������Q?�m�71i�V��[���V��{W��U��*e���=0�u�p�j�ڑ����ж��;����,�U�:)���kFv�;^�����	 �g�h������ \,m�AV-��Å�c�$k�ߚ�M��,z��7](�W9���J	sfE��2�� 
B���_/=9p���P�B���*�>1�''l�l+
�y��
"F�'��m���~�褟��� 5���E(-jO�<_���n��.�?Dq��N5W�^᫖�����i�&�"kﰴ~�FJb*Vg� l��[���څ����dN*j�Y�؈lZy�Ca���l��BwW:�d��*�
�+�@�����C�Dx)�s�ە�]:MvhP,k�������W��V9�~�~��8���WJ��7�i�)v\�nc��f�-��me�ڲݯ���@���)�@�F`�T�a�K{u^Q��f�ؐՒ�I�m��������[�t������Z;t#��@�w�Z�n����?p�=��S^="��V%M�-���Wj�KK��������\7bU�%�x̃��20rQ��.���a������O�v��l�C��_�	�X�0im��4lA�9�Rds��S"͙k����Xn�n���1/ɠ���o�Is��1{̲�X������,��S?�/:�*��P߇/��U �B�w%Nt�_@6Gh�y��R`���d�D�d��#F%��vҒ�J��mafD������`ϸ�!�����Uk�O��V��(�2�pZ�XӘ��L�4]�x�]k0#�!%��19��C��f�Ci��Dkm���U�@���������m�a��|�rz=���gtP;mW�&2���0��G+_ ��Oͳ����_�ni��dL��~�?*L�� �f8�r���D8��ױ�l�Wۜ!�i��x|��!a��h��j��p�؅�A�qmG	 �����c�r�M��?�=5	ygAJK� =�8+CTlyS�l�X�a�i�RV����J(��-�	l���B
-j�$�jJc��vb���'��R�����%��X��g�t��*x ��}F�����,`�VG��mj�um���y�)�h�'�,�VȤ�'}�_��@`w2�M^
����۪m��f~��+eqP�{����L`��f������	�� J�5K��|$,���CyB��uØT�F���f�����q#���t*l�V�6�P���G2��u�E"<�M�������1F՘CO+�$��[��������|�Ƹ��n�\�Y+�y�����D�_���s�L�vp��?\�D&Ù��(=5��
�:FjO x���Li�8s s��'�9��� #Y� �N�ڻ#�W!5��Q�>C ����1MA��@�W�`���f���Y��b��q�HF:��u���>���Ki6� ��W�=��r��J�����f�Ʃ.��?k���w���u4A��L��fB�_�A$獠 �t8t�ʔh�Z�3������&;�|���	�~����kC�0�"����Ɂݵꅙ��L2"��%������^k?�#���bi�Y�x��aN+N*���׹
�Q�B�fXR?A��Щ;d�d��,����2�~fɷ�A� �+�048EZ�r7��k��t��;�3J�� �ʔ8^���ɹ{quq��d�J-$Z>��#C�@�j��X��Q���wG��pr�����_��A���8P��� ��t�� h�o��c�F7sֺ�sDۉ[B�p֙�:��`���-�0v͞qH!�!K2�FD^n]7::-a���#�4<�H;����-�FP��;�˭�^�,���BO0iKl�CaR�����Y W�;���ڤ7=�d���4Ii�8(}�t�K��h��0s!Ή��W~3O}w�D�-[#�6w�9�ub>|�G�H?�����/���LX+<���q9r�}\����#��&���]	 s�Q�"�yQ'�XxuM�7�j+W�=���kq� x�/�.1��A���0  ��DS�倚`"��oJWf[��� �ꍢ>��&ר+�~�������ӻ\�N�t&(���iD
�o�����HɈ����e&kP��v�u�me����=rXz ,�z��a��2��7����4Zn����T�=���E�g$�p���{��ڳw���+�5
��)�3���W�S��>�X݇��}��r����'���b���f�;��d�ݍu�ù�JM�9~����0�i�j>~8����@��D��Ϡ���fl��m�@K�w�Z�R��c7>d�E�`\��u�yI�n�LW�qX|H��D��Z�F,�H"m�/TZ����Jv��J�f���/�C��f?��t�(i�|8���?���<R��ff��ؘ)C>l��6��d���]�#8��v��=!�.ΎJa���QOV*�E�]�[he�L�[|�}PHe��~׷O�H�� a�e��!��%�A�w�d��p���^8m�g)x2�����j�3y4��H�⨤���,����Є��"Er�.`w�۝9��l�N!�-G�����|}8<���a���������IW���`����S�`��W->�&��#i`Ck����n�,��R��:� �'K6�AK-ܰ|��Nk�Ca�=x�������\Z��Y~�GT���ix���߰f���2�:pJT ��gg�I�o�U7�H G��˘�M)jȞ3)!8Y�� ��T
zˎ�l�:�i@�1f7o��kJ�^s��z���f8ӊ�o�*/I��^Nf	�<��l��Q��K�a�����o$��<U�����^h��V�+1$D�o��[Y2��P����y`���ׁ�}��P�a:���[/�Y�o�Ҏ-��dN�A�<�/k�4��Rr޸s���:*�v��d�����Ǚ͛��`YM�Yq���ܱ��r��a%�F}���J�cʂ�U��;���t��,������;��m�ׅ�<&�XO��3�����^���h�,Dt�i\�{ϜVV#D}�(�0ą��qNN��K*�x(�ٿip��,z���q�cɡ��E�Fڙߔ�߼g�Ѩ�i�v�Os�y_(��C]3A���S ��Y�����4��e7��s�}��YԿ��+�ũa˜v�������W�p~�E�3(D��~�����_I!����k�w��N
�=��$2��1�5������PD�A��,�nz��?4���6
>4�ƷG���� n�������'����ى9�<�J,;R�&���V����#_�!�$y �,�1��$_�����hlZ<�����P�D��s=H���J�l�fEY�;��]���^8����Km�%��V��|�VD�EV�Y
��7�4�'{�W2u	Dhqmu�GH����`nea^�b���n
ɿ��S��4��杻���,��f��/���]/@�8N�L�FI�D�
q-�����k�~�?���Z���fB�a���h�Ay���f12A��%��L�����=.I�uID�)����x�uW ����}G��|�Q�&M$`i�#_��J�B�V�?(�H���p�*��#�sG���pA�=�z�	0�-�T6�H�q�w�[��C9و��ը���r�4T���`+��e�~+#>rfJ|����.�[F�e�N�v�-�(�Gw\���0�Vd��'?UI�ԏ�M��M(����N�����Y�����@����D�ȇ�� Z�g��l���02�bﾤ�^�t��e*rzт�UgR���졅D6����	D����N'<U��,�!q�?���ᛠ��%�4<E�
42��_c�AT���8H�����֛1$dP�O����y�+?s�F�������T����(�捭ζ&B�?-��g����G`Y�)�|{jG�v�����ڶ�B(-�r��@M/#V���M?�����&.��R+�*e�z�p�K�vZ�@Z��ے�j�L����U�3��LFR*�͔8��0;�^�{�\E��F�_��[���������jᄽh����iS��K��ޒ����V�� Xo��'�p)�9���_���'�sz�QO�b�N�= �S��6�V�'�"����E^��)B�(�Z|���$'�#J؇_@<d{��b�V7������� �����Bu�e��L@�|��nJWl�B����#�\'q��T�S�����<��pk�|�F��K
b#xqg��G� �("Y`��]��g�/���=ӹF�ι,s��۷Õ3��H.:G���zV�ɾf;���� ���F�REi���gf���4uRR��v9Y6�����V�ܚ֞���>J��ǉ��I��ƜP�(�J���w�:�T�ڇ���h�G�o"�r� z������@� 4/@:B�j[c��BŶ���\��C)qH��@&+�N~-&$Y����k�,:��N��Q\��f ��H�G�fV���U��נ8&��E�� 1x��R՘ŗ3��b���Y��������@�w�N��Uؙ+��(��D���./S�����(~���WOѪ����e��md׷Z�5X�p=6��\�#m�b> �̩��֪܏�17�����Tʗ�i;���o����������M�}k�l���B] 2`A��ԙ���;NH�\���.�T��;���`�@�P�,��<�VWPq&�̀J~���)�������e�Vq�,�AW83��,F�ib�)�'���#������Uh��
�(A��㥑�\����$��(�׉���A��5n��3�+{xV���mZej��I�h��mD��HE ��DCӵ߰������������|=���#Gv"Qc-���D^�7���w�kY������>7�v���ȭOW�O���'��g�:����H·��-���[���xc{���S��9]iP�B+�O�{{Mcj�$�s���A²���
�}+�[!�[O��AG�E��]!��@��6�FI:u��W�]�W������5"���������s�܍ש�i�x�h�s�	bK�8�x_�ɀ����^(�� sO���k�%�`cGg���3�L��1d'����;8YD����.�J�SD��K{��3H�J�ke�B	��L��H��� �]|]}��n9��n�UH�O<�i��w�\j$���a��˓�u���U:4l���x�!B��D��=�_HĚP��0�v��G�:2ԊCH��6Z��<4�q��h�萣<"F�/��pX3	��k�ݼ^�h�5nj�:f�"O�����mZ��>�>�����]��������F��O�?[�?6�����0�\�S���撐�)�}�e�wKa���>r�8X��Gf]?d�H7��72�?�5�`�K���,���C3���W�w>�?�u��� V�#�u{b��
l:�R3�n]����&��r�E2Z{j�E�5��N]�US�I��:qd�xq�����θׯ^.X�h\,���'n+�y�fN�AO�Qr���w�a�V([��ׇ�S��mYzd��ڵ!��%�Zt�>� �.�]/�֘�맓�nl��]�|h�l�6hN��9��F�����/�%�]K��삀P��86��F��tQ�;ԣY^��)"]����O4tbQ ��7,���x�Gt�Vm�Y��%t%��(q<�w���E䄠.c"�Tj�E�s�yeژn(����`�����7i��_�o���	|hDl�'���.�`2A&"B�oC�U����C
�k�9h��`X_S�������h�J�/�]l�Y3��{���8�0�m�=�Zoغ�����.�Bw�[�9/В'�\iO-O����y��K�*��/�V�|��s� ��e[����ؘ��՛5Kcr��-�Ȯ�i2b��g��4�v�����zv)t�В����CX�0���S��M4�P ooY����6�T�Vd�x��A`�_��/n�:��ѭ�3��!`>����1W��MS�������t�6��s1Ƭ�^�� $ֱuլ��3��T�8,�! -B�b�ZD�?׾�w�RuO��h�5�/*
������#�:�n,u(�?k��aڍ`�ګ���ۑ��I�{U+�샏�a�n]W��V�������{���F�֬x}ޝ��|�L��Bv�.j	������T��ܥh^~S*�� ��k8E����꜂��8�'��O�L�Q���v�Y2����%�Y�'5�"qF�ȝd�P���}�¿��hY�owx�{t��K; VG�T�~H�V��\I�q@�e����x#B�@nN�}��c�>"X�[��3s;Mb�����q^�p'}i�{�i�~I�v0��~ib����T�}M�RM2s�ҩ?!/h�(�W����_��[J�X˴�0��g_�$9*ySY?����j��N7��߇=A�꼈-c)�5����>n)��9nG{�)PS|���R��̂�`��p���c�n�Jv|���қ�}�Lm�Qg�����lKkYł���?sFG�i�,1�i?����g�����4���u��<�K ���u��AOx��j�*[k�`�Zu���s.	n�)�6�О�)�~��?���j/� �EY�Ym�[�&�:=���sR���q���}���b�]EI������f�^Cw��>�V�������''�HK=7
s׺��5���w�3c��<[u>X���TyM�W�%?�U\jH��H��g� �Z@&o������Glg0N������>S�s5�ռM[X�%HtC�C�hgj� ���;$�8EL��y����O�2�5M����=�����M'QJ8Օ�55X�x6�p��_��ɓ
'[�I2>Y���~N�UG��3�CT�B�sid�}�' �|Q.6Q���6�;r3<��I��=G?�������3Z�<Ip��wp���'�=w@Υv/�j�����Ń���.[��g3���W�)��U|�i�E'� jZŁ�^����Y���]-��p_���'�x39?
�����x
�ɖ���w]��PE]a{u���T��h�w|�X��mZK�.�ok�vZcf3ނ`�9��V��u��z�ʾ����W�2�0�+�z���\2dUex���
��U���67Rr���0#�zM;�1q��	�|�;p��	r���i�~9�s�N�w!l����(Ce��Ձ�qsO�G�q�4*��|��>����w�]Sˍ�g��D��]�]�I��3��g�?^f��׎[O�C���ugJ̖y��=�瓖��Aq�cWד'�S
�}%r���l�L�bhg���Ci�p�U�.S�)ݤ��ng-�C-A`I�6^v0Kd��v��A_��=�k'A��ym���&�L�=�Ff!^o�V�=�a-���I�Ř(XhP��j�80�@�G\�T���#��	��I1�¯D��0���UQ�8�v���-��N�3c��%�3]L��}�~w�m�m���Zd4���B�`?���_Āx�a��?>�21/���mL=Ǚ��m�N]���2����1���d]��ƒ�fVr�	Z.sX*��jG��i"ߔ����W= &��!�N:���N`�a9�
��ԯ"�A.#jp\&\�v����RΨ��z�<��7 <�7�78.�J==j�ڹ���Ess��k�M�|�'��^��8��q+@&��f j�A��,�YG�����J}9��Kg��im���m� �{C�6A�4��{y~��Udt�SK�s���գ
������8�}9��O�]���K��lݸ(Sn	�B�W���"q�C
����6:M:^O���yTs�Y��M���(_����)4�F��aRI	{[�h�P�?�ϯ��D�"jQz���޺�ԂIZ׈��U
�;N��nY��F��3�J_/ T6�P���M=~�c+��A+:��X)(͈@BgJ㛩m<3�?�OhR1��6C��T��}����ئ9��&�^�*��������G^�T�����u.�Ǐcݎ	O����)	p�Q��/-2k��HQE�|(a1Ğ�:!���0V��yغ��9��~Y��ޟ#͊u��'�-&7�`&l�|�I���Vo���V:rє�w$��q`��u���3R�۞�^��_Qκl��7U	:}�'_������a�Յ���N���'�L�d�'���f_�/n
>�j�G��E��!�=b®�T��$f&�]������WE-��AQ��{T*#�l�o����l���➴R��+B�ǜ��z`T�࡛�d�3"�t6�����\ȿv��,"�B����Z*/�F�n�"��uZG��(�ss�IP�X�!��_��F6�oz�9�4��i��:��҈���R!�\�R��>~B���qH8ޑ�F��`y�g�9=,�W@ hS4��e�j\���,kk5�x(�q���,�����=���s�d~��H��SI)a��턈�L�lA#{S���=u����w����	�f'=L%�'Ԩ^�
h
.��i����H2Ɗ>��8�=�����@]�ki#D�v��ses& �i�h�^
�鯟iDLܽ%Yo�"d	_�T~V��-Չ�8�eB��(*�`��:W�Jv�t6�J^e_&��?@	-�9a�WT�=��z+��%h'm��= �C:��\����˙��H{[3�8������JjC�����T.���wD�ՌJg/�%���N��v90G�����g� Z���A*�|�YO�w�Luž���������p:�Ʌ)�`��e^3�g����F�4v\s��G�ױP�ЉQi\�|.D��F߸;�������N�I�(Gf'^6����w���ι1�T��lA�d�v�����1|L���x�$�W���>@C���t$���BI�8Jn�'��@SLJf3 �͐�����5�>н,���+���j6�ȅ��K�|o�ol�����T5H����fS��M��D+0T���r�]�ب�!Bqi�pN�:J��9���\<u7�C��?_Nom��yɡ(�#�x��cmⱎĔ0�l�S�Z+����ղn�-i�Z�uqv�
�����>zd{)v	m�����ԙI�\�Z��lz�P�-�4~���}�c�gC��R�N�8H��H�g/�
�g��rq5dAu��T~IƐ��������q&;�q �~���/�go�Q����좜&�gc�Y�R
���()j�3UYg�:�m%����J>�)���{:�:��']c'Y!��*��x���	��2 EFdsߓ�D�&���y�$�Ψ�`$x���~'�^��N�D#a:����V�s4�z+��PW��L��.�J�BЅv�Nd�Ɲ��[�I�:��lEu�d`���6��������J$b�dC�����%\b��H*�ck>𪶻l#A}�a�;�E�4$��(e���u�2l�V���:�N-��7?��~��M�6 G��0����@��C�
|�d�ؚe�u%�\B�=	8L����F]��y���`��UTA��]m;b�6(���?!餁I��������D�FZ�@[�NB~�
a���ټ��i��H��}�谂2N�cqb�f >FJN�_2����=I˦Z_���i�0�^��\�]Hz4i�[�;�������T����U�Э|ڵ�e-7KO�I���ߑ��+�zkT���l��C߆�1�����^s���<�Z�����B������)bU��fd�{;�D��>��_fw���%�(hg:P���E�#�f�f�$�m�6y�K�<�yɄ�ߔ,���T_df��a ���(����_��Ī���N0{Z���O3���lC�o����x7t���{�����&��Ɍ�Ur�1"Z�Ջ9��8펬����Y�@�s&~� Ì�Nͫ���n�����_����R�)���	;',����⌥��H N��j{��i��B�O�u7]iYO��X%��W�=g@����T��ۀ�����Y�YCT�gΔn���Ο�׎�ɤ���1˯�����S��lک�\s�w(����[n����©�sqڲ�H�[���p0ybB(xg��#�1��CD��ye��o�ß�Z����+<��Y��*��֡��f��w��6N�f�T�Ҁ�{+��ٻ�CV_�ߠ�Ek6��O6�.���d��� \��yT��?��(��$,�.����K8�x	s�[jB���6������69�Y)��v� �"����=؈-��+�7]��Xm�)8�s3���#s6�H�D4�y����Ħ���{,�1�r�p�/ls��wQ�H��>��0a�6�`��.gcA���$8�(�{��V2N��v�g�j䓴���4����2zC�fƺ�\�l{�$��[��u|�箷���đ�Ykͭ7�;}>{I�������đ,�6$
����q�
�j� ���ߐ�]�dJ����)=��d&���v��U��Oܕ�@�z��į�D�~pH�T]͋�G0��М�7S4�yn)v��pc�Z���Ms�HYC�fё9��QD�vO������ǋ+g( b+�2й�\^��iv c�߄z�S5����fy��^Q�!f>+�{�n3z���M��3'����^2�K3W˖�v����,?xqAg�o��W�H����ou�5�I���޷}G��}bޕ�V��UB�#��c|;N�y����qO���る�w&�Bob�y�l�ח4���ϊ2Vz��Jd��)�0͢C*�[H�ߩ���ʒP�K�
ȉކ�W@Yf"�+/���d���fV�$���mc�?� (�[Ũ��z%��(bN��@G�L$U�XU� ��ͷG(�����W�,��E�*qdl����g2]q!@QЗ��՗5���um�1O���䎋љB��N,��H�+�<��*)oG6 -��cn�f�E1�.x���%Lߩ��ŭ���t��m����{�F�.�PX;��U��/&a����R㓟����YVa0Xd�༎��a���jܓ;�	W[M��m��,���	�=��+:B����c��0���z%�SN) h��ti����*����Վ�"�4�2y�}���x�[ck,,�9>�/�Z���@_Chn�[U�hN�Z}��O�F�5���f�<��7E@l�w���cx����gS��G�,��i����Ő�X铮�쎚�>U's�,�L	v��i�x�ӗg�6W7ڮ�IL�^S[^.
:��C��ѻ�%<n�ؔ�:K��"�;��hg6��Y�SD$��bm$F���<���ba���&,?0�c�:&a %Hm����G��~�ʋAl=)�r)����� �$;R,�(���D�Tp�:����&�=M�n9���9�ܭy@�!�����gJ�WG����"G����t	�Rl���ᚢq��ݿ>�N}�ī�(����F�_>Q�:,��Yw�=�֜2$���B��IdB2v���B���'h�b�ΥY���������_�J��l�an=��C���0��T ��_O�y̐��R���S��U���	q�J��8��?�3��%@�#�D ��[���am���͂{�B�z��As���|�j�b�� 	}����aՀ��_&�M�q�0�/y?:��
	^����5�u͕gw�k�,��$�����{�M�F�Z��!7p�:��]+���n`��|���}Tj�#zd�/��Cy��~��,U (�QM���T���v�N'��]��ܓtG1UXŶGt��%���7�a�P��e..���z+yٌ���#��V˟�0�����}�sκ>mJHy�6�కLd��H
��V����4b�Ϛ��I��8��?,XC�j���訩�v�A�����i�ߒ�.��ES85�m\}[YY�
	�d�r�pF/Pz{��U�j���T�Kl����`K>��!�+�g�ٹY�L��_w,��_J�I�ڌG�>�o����WQP؜��9!�wʜ�^Y��@��V=��bg�=NR�h?��	���i�6+XÕ��
����O���L�N��a�5jv0�	&G�"����Q�@7�M���F�n��ȡ^{0�i�i?����fS��Klɡ$��#���k�G���RZy��`�ƃN���A������{���8#a���7��1�$*��FC�)�I;K�϶���VN#d�1�Z���?�3VYR瓌���.�����ķ�
~�^4L�<;kzW��Y�Q��`Q�g����_�zli��ݓ%�X?���ʕi�΋7m��#�;��VE!C����h�J�Q�CG29S'�Aȕ>ԩU_v��+�y\<D�C5v��bb��!g+�4�|���O��ѫ���@쑅 5�Ģ���+�zY�D�ř��5��_�j��+7q/�|,�;"��Oz՘cr���=6� YTK�o:�|9D	L+��w��8�l��gV|c:|���6y��1�o�-*��XL���ywX��A�4���dT�����c��6��[�Bޠ��
0�J1����&��_��7���$n*b��Bѭ�2W<3[�L�*�I,L����4����7?��;I/��ǈ�wƸ���O�=�H}$ɠ��dzr��pԀi�}b<��I؆:�g$f��/{�7/�I���>^?�����xG1ɦ�>8�c��E�A}&�A �E���MhHw�/�r\���S0Y�L7���~!�d��i9����KnO�SE�y�� ,֟�����>�v�#`�/���u����$�\tZ�E�8y0�,�X��D&�Jq~2Yv�
���T@�=d���'��Fqq��������vP���&�!����7�ʗ�ܤUIk�I-�,�FE�#n�f�|�n��p� U:D�^���ןET�X�_���5��T�2+%��9��P�zy�������7�|���y_�g~U>eK����,*�f�]�:�.���O�����3��=Sx�u>����p:�l���5����,�E Y�3Lԧ1�W�A«�c��?��a�挻��ƹgCG�j��]�� �EG��Ͳiɒ F^�_�s��� >��R�oqT�/��O��Sс9z�9[�fDUb�����t��t�Dj/K��8T���W�RR$;��j��k�tWo�Ō���=%�눯J��;;G_Z�PLd��_D�� #3��-1�_O�/Y��&>�zK����G�GH��e���4#�=ŕUKQ:�n�(�͇y~��"�G��Z_ x�RYa5����X(�'N�ԓ���@�l�ը�����W�gzc$�"P ���5�x�3��Y�)Pj`ǆ�v��`�~��E�7�B�	��*"�KL�i����kv���w����}�dN�/�t�F��xE3����G!IU����+�u�nI�B��42ܪL�{��'ME��z�,ړep0�����<I1Z���yl
��,��mPꘑ�Ne�O	@�)��Bk'g�r�$�d/8���փ��[W"�.����'G���2��:�u���hY6�k`������jgM8	oI;}����U˕n�7�P��w��48�4
�9J��.\:�#�1u�7&�#���|Xt��mZ/:*�@��uZ��65�U-L$圈qV�NMXt��5��wX�:�U7�yR9R`"�Y�a
v'�A��M��ﲨN�����N���9�4𰰞XT�t2���4=�z�W̒�42�)�p@�Pw'��b��A�����7��\o�^�C���QK�����[�������U�k)��?��s6މ�s.w�݉�#�����z�:��,�k4_��ϥ���)��nTo�H�i���K��`'� ��[+�Vi�^x�[�Sڣ�J;v�3�,��\�$�x
�;hR]Q��4!��o�[#!~�f�:M�Ϗ�)�J�+s���MUD�>u��E�����2�3&#���s���X,�Y
i��~�в��kJ��ږ�&�e������vGn���My�RT�~�&�\b@�6Z�k�\fsbݦ�����{�u����q��2������y@����☮0l3f�{�� �:�����,���]r��T�+�6�d��v��w���!^��N����WO74t؀�M��?&�/��h�hӄ��6�HW���<���W��]u4��C:�B�H� ���)���֐@Y)D}D�1!�wKuD���8��aM�`�
���D�٦ųs�Q�'�LHx4|�����ˤv�_�2Yൔ��a���|����(��U�v�f;%I��֐�c�ά��ύ@�-�f+!<:fɩ#u�Q�0*���% ���j�w��vLH�4�PdB'g��8`'�QJݰ�o�[#%��
��6��6���p��t�R�)��x����N�:� 7��D��-`�N���-�Zeg�n�ڹD9��(�{/C�րsd�U��,��P�_���� ���x"�K�Z�:Yh�R�4���u�f�٩�Ef���M5�/��04bC	�ʿ������R�Y�C�y��"�-�\��]7�4�2���t�w����Z��I` f^�6ˋ V�I���'��	�Ps���\��w_t��U���qǯ��>~*�t�0�@5������,�:�2�V�g���)Á�7N�=�� J�r烢���ǩ�
�p���>��ڧ_���p�1�m�~/̣(��L����Ն� ��
��㟘}��\�XLj�p͌��5}�:g[�h���.�o�*L�=O��x|����w����s� �s�^ 0/'��щ��\x�����r�_G/,'�4<��Ǳ�E
Z2�?���9�T���غ�Pm}&�{Ђ�a뫰UzD[kX�3+�(>�-�nN}q���l�Z��~��J*uЩ�9�s�V�X��#��\n�^��"FDv�K��+��&֌�}���Wc�L��d�4
F��h�PnVu�F@xf|Z�Go��;�w:�� �+K���<��<G ���!�Z�����{i�F�n{�bd�*�[�wV��%���dHb�V	�%��7���wܰ���۳����pAߎ;;v��C>��rH����<��g��F[�|�>�f$!���Č��"{)���[�9G��鰋����	/�=4y�����N���lOF�'�
�CݵO�=��InGn251�g6K( 5���w�ǌS�ao\#������p~8m���UL��\0��s�!�����U��Y	^i���-��S�Uƽ%K��K�X9��3k� �3O᱊�A�-��v�f�������_!D���� �M�]�~�[p�i/1M���R��_��1r�ia��J�<��i��~�Ĉ&�dw;kɿ������+�L������"�Ƅ�/��Gd	��~��]|V�t��_J:�"�<~e�uK����p��ph����T�b���9�IŁ@[U��J��A�Ձ�Fe'>h��&"�n5%���p�`a��	�?��إ:`bK�?5�ԋ��pi�DZwʎ�Mb�	`5��'�2#�I`s��d �Ư����/��hK�Z_�8X��4��r���a���t�Ul�5���_�xNg �C��ЯF��1��[�Ԃ\&�}����3�S3��^�w��!�@ԋ��������'��l
3O�o��(�� �} ����8�-�t�]Q�����l� �8*��0����ZRp�����=�ا�ȃ��BR��u$ly��FƊ�H��i�8��5�6�p��̃�s�I�jV �W�����+���"N݁�ƟlL@_�U���H��VV&�{leT:�(���c�FFԺ:O�Y�W�O������k��B����4�d���8��c�L��bmNjbnդY�-�+�o�c:
��t<]�瘍]
�P7���r}�HV��A�r��6퉀���&g)y�RZ�ST��|�Xq�F.�nP�PV����-(jom��|S4D�.���g_j��2����{�ov�Ҝ7�#]
'+��pT���"o j���Xej��+�z t�%�ݭJ�q\F_O��7�aC��t+�V�@�!;!Q�e��.���H�Տ�r�&�H�v�����