��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�Xn��8��ՍM`P/��8TRV�Ox�	���es�&������Q�i}��+��:*�}��( Ą!p��1����,2Д��M�O�8&/�r����}�ŵ.�����_60�=}���A�_��"��Ƽ��T�,�*�!�S�>}6���P̠��_E�֛�#3���M86�W]02�5�4n߲5*�y�%�M8܏�-^�;De�J�����"L�C�/�e�&%'/MT�>�]����E(ko^{
@*��^�`ǉ���VC��A�i��L�#�H�F5ho������iG�[�]m��()�� Vy��f?l:������
(hqb�r4O1Ї��*w�=,�V�P��uo�z7}s��p��| Ӂ�Y49�Pgu��öy&�@=�d�}���M�_����k��˄E�U�o�ιSg0�^��c@�M��R��������3�C��t�F�"�rI��Dx�)b,B�2R���T8�I�n0W�ĕ��1�+$mPdLNu��{��^'�Rw�~�O��$K��\*����t%��"ߧބ�� ��&l���ق��H�$�}��m��ꗇ8@�	� �����׎D�5֤�����M�%"�7�
�5��r�ʧR�k]g� ���:FYȌ�@#mʽ�,N����LbTj�n�=�X��i �;*��>�d�A�"�hF�r����6or�^3�m�3lG$��b��Qp<������e���,�����P��2�{u6�(ֈ�Ψf�	f���nw��D���,�G�*�y�+�hM�,g��Б��n1/�z��8q��7���2B�u=o��tfv~B�$ɰd�(_:W,���A�V~-��X�����W)����WU�:�a�����l���{�-X�=��?���KKD��f&��~�'87� �s5.�����%ue�'H�RI���sPIW�?A�d<�ZX�!x ���scd��>w����Ȩ���s��;��"�`�3<���Y"~X�}���Ͻ˷k�ޥ��L�H��W��8*6�F�CԥR��L`���޵�И��0kFiƼ+b���qiE�Z�>�~~	�;ȸSb������P��Yl�-(a���AsQ��h��(��	Gnd��΢�8�((��s^a��Jt�|ad�"Գ�݄,ˣi{���j<E�ˉ�SS 7�M'Z~	�Hn�;3`6�����������R-�o�+4C${-���)�|u�o�ʞL}_��LY��������@EG����lc��r~K�Ր>X;٥����Q��s��ȇ�]���9�4p�d���^�xv��|7п���h���x*��ըә�ţi�$�;��#+6�� ��-�c�_>Ӥ���C0D�Ŏ�����x�f�O��ltq�7�A�!���'��xb{br���A`�ú���xPeF�1`-����!���M\�,`�!���V߿�ǸZm��zfs��l��ޘ�V��B�G�Ty�@�f�[9�|9D�=�%y
�KZ`�]�Q7@(��g��n텻4\P9�H�b{�80��,ʐ!�"��_]l��E��{��tD�͊�S[�z���aLQ����idU'��s�Q#�*A�^'ϴ9��Ȍ*��:Y�,F"�s
��S����\䡳|hZ�܁]H��*k)P�0Zp
t�G' D�^U�Z�i��+�at��	k����	���b��:�>��v�0�?N��)kY]�|����艻�	mv
]���ߏ�ߘx!�"�bUc�x�8C��eL��k����rG�hі�	~�i��]^~zLo^E(�`jkY��?`����p |�jV���
(#� T="{A�t�:^�o冲Z�I[�Kq�z+�v,�h���~�c��,M�7��MZf[�:DB����oaV��;B1�,�.j?~H��X��S|)T�����)/n�Wn@��̭?�$QZ�x><nB�6!0g��qK���#s��W�ƻ~�Y�ǣt�f� �'�j{�]�!�mms�Gɞ�!�͆ �c��h[a���u]ѠF�m��8�LKY%u~��
ѭ�A���B7 �ib�L�^��O)t�I&
F�	�OY��g��\Y
WT�Bhެ�j��z����C1Q��N�~[�l{��p��%!7r3�2��"�nM	O��s� �I��&B�Dw��>��	����\�bU4b/�Z��ӌ>W��{�$��b��W�|'1}Y3��a�Y�0D<*i�+�Q���U4��k���S��N�]�)i�3p}��~G�k�+ށĨ�(mR�S��g��0�A#z��t��ӏ5�y:���7�I4u���r��&���{@��P��O��!O^���W�H	�N��l��j.����縲9�{A�����M{9}���n�p�Q��Q�aZ�B�G�m�Adc��r�-�P���W��CC2�Co��()P!64yOpƙ���h���q���б�>�E�
�����6*����zk +�"܁B�l!y2*q��a0ut;��O)r_hj��ki@�<�~��K�~-���@A�i�<��O!�����[s/v��_��:'%��w��)_H���tc����_@��*I2����`O��C���x���U��ߣv��N�8�!�@h����V���̶�3�54LG���
����	h{�KM�Q`}�V�ſ98�M2�ө� ;���,W⅗���*E���ϫw.3(���7a^�5Y��w�����7	���N�
)�RSPx��`k
�0���w��>RUZ�[u��\=~g�Of�d� +�Ғ�uD�ٞ��|e��0�8�z�gŦx=R5�I�����r*�Sx��f�ʚ��,[8�"����n�%CX�[(��v'r%���p�lu�~R6i��%~��K)u0�;�y����b�㄂}��T@m��#�U�C���R�}�2쯉��"�`xHv�o�����J��������?���µ�d�m���9�S������
���8��a��@�k0�c��ڟ5�9�a`'>z	���Z��|��Y4�`�P���F�M�y��ӥQ�++ uXmUs5��azV�̸t,o>N��۹(�(�e�8^������Z��E��cm�G!p�M�=T\T�ƫ����!<��7��)�P��P.�,��f��Dٱ=��Wa2.���@-葧�0!B��<Q�,e�:�z�d�b�W3�]\��ǉ�j� ݤ=e]�)
pH�9B���}��	+��4�] њ]�F�KV%�|�L���/�O>7���W��
���&���2z�4ך�zn��@�����ԣDL�2�o$��iKƛ�{�����S
o���CE�B�!��?�9p�a4�|����@��)E�-��^3���<|(�>�w'	��M8�r�4,����r�JE��,9%�� ����
Q����ր�b���g�xC?v�C-Ѹ�A�J%�;��f��./TbǲiLw�@�T]+��l���%���^�Fm���N<� d1Ԯ ����?8�8+"y#�&ieKΑ�zMʟ)�j��ʦ)��x�B�=<��y8�x\�����7=X�0��_�r��M�>�r�K����&�?$-�����%e��$^�O�Z��cSz�}^��9	o g0��Zid�x���ũY�iG�"�T�����a���7�~��=�כG4���֐pO�l;��f,>���k�������y������v3,2	Ԫ�0ު�".q���߃��4�2�0觰��|'����9d!�ѦYȻ����mfȝ_�Y;��/|��VT��g6n�|o��A�e���Ke����J�}�O��4* �Y��������VTt?Gl�f��&�j�,�6TUw5O��=HrW�8����ol�V�d������F�{ykܕֹ-�'+����q�����:���b��c�b
S�,�S]�h����?��	4��m�h�,9^�c!�YJ�M��\7:uU_�#��zVY{�Xj���R��G+y�pk�ƀ��Cդ�	�x0<�kn���+�b4##��n�zE`0�Ӫ����t�Bނ�F��2��Ҙ.w���L��%��-��F����IЙ( �~h''jZ]���C���l��D�6[#�w��*8���B�8S�3�	徾Ў[~�m���P|��쎹>Z���C�9�"B�Z���Ѧ�=�B_~��&�zjog[In���#�8S�V*q�yύO�^��P؅�����=��nc�L�;�h��6Õ ����Q�^Ր�:�ִ����t�|t�M������}�>���L�%���d��a�� �����ͮ�f�����n׈M�9s��&x�@/�JW~x�"M��k-���t0��2�."�����," 2E����k��Lp�	4/gL�x"�F�K�%k��kk>ɗ�����U���sik#����}�l#\�4P9��ғ:($��o�+oa/m�$RgM�	\wi��w�׊�G��+c\ 5�4Of���+AW�W���Ɵl
�;P�����RQ���w�#�?io��;Q'M��d��]j��o�'�>B �1܉Y=��Z��:aۉ�Q!�,���hR�e��K�m~�t��D�s�� ��q�7@p�Z��3 c2Z��Z�f��A�33���c��)�"=�tp��hf�5��c%�[��yo���s�뭼���m���M	�ga��
??���6OY��_E���ܠ�$�c���9|�Rd=/~���"]���h9�$@�5��9�&$'�4�{Hkْ+�震2���2�1א֣qd�!�|�Ol���ެ2�u(���nd�9�e�m㜺�b|�,�DA�g|�+A�7�����Ur��>��X&#*�2q��9�,��`�I�w�TՓ�� b��2�Y\���������;��W�Y���x������D�_�?q�f����Y�!���/��m�e��Q�,B>=E�C�WdU/~�:�pа��.�l��������LZ��r�Nȩq�>h� o/��춤a2�D�jOqJ�/_E�������z�`h@�6K�G7W��n�(��P򇴦^���l?��p |�N%��Z�� k̡&�
��8`�x���lH�����V�o!�`2�ɘw�?�]vz�綫�BOQT�`��w$���b��>
�qo�+�����Ǖ��Y���b���HߢϏZ��"p9kIقr�$��c)0O��f#y�T/��<�(c8}/����:V}����
?13���ݺm"6H��!?X��dgad����2f��X,{Z�t�=�A�\#_�BP�X!������΂|g��*�_1�N�$F�3�`4ݶ�+®(.�籪 ���A >		u�'���;��=���w[*�Q��c�u���W]��e
0p7��^Ϥ2��4�n�1Ӫ�_��vj��m�m���������uZ�����f64&�� ������ir$S�̊��,j��)z���8i���z�!��W��9��O}�H�i)��j� �N25�� ��9���A�uS��+=�����~n�	ta��&��� ��H���@牿G��z�#JO��j�C�"���9�h�Fe�v�`��0!�����'���6��u�8z{�C"]z�$ �����l��GPݭ[�C<K�A��jp��}�W���6:L	�Ny���v��څ�De.��*�WB��ए��5����,�<��@�G�n�1f��@������n�ܦLhe�Q��E�U�����K����f���bꇴ(ҡ<��),�/l�(0.WH�D�ƶg-)�ūI� *>�����AQ�~�R���?&{"N���
u�����w N��=Cަ	(
��#4�D�h+���@J��Iwd�'�b�teD�Bˑ��n�g>P�}�υu�9�-l�^�I�
P���X;�\��ǖ@�T�?��iK�q��byk��l�؄\�Ϙ~?��y�.�=`�����j��L{2C����T���?ȴ�tXk�O�����=Y���c��|~kM+x��A�L�j�pxU]������M;���O�6���8\�v���\��ҠkdZ� {�EiEw��ȧ�ە�'��o�(&�����ߠ3T�%��{��$'k/��]��%�Dn����:�	v���$W��i)�>�P���0���ᗼl>^��I\^�7�������˷�º[�~��^�/h%���`+t{ _�2UC��g-�V���K����6��?4AVyB!۹[cj}� 
x.�9QZG9����q��B^��A�&"FQRE78�מ�
m�\K���ɴ��vr�Ğ1���g���U�g#`���̊?Ҧw�I(�jfX���UPq=���:�{wmQ�N���^沱�o��W=���J����n���d?�zG �
a������a�J���7:��	��i!:�R���G�و��z�V�s�b�m�E�t4���S����]��F�4mr�4�$���X���Ɓ�l�f�4;y�n��Z�yA���5B�3ч�b�c㩱�%��ILSxo�"�f��ʯ�W;�������d=�����o^��Ц������X(�5�<W�q��_��	�f˘��z�jh(�o{��/�;F���,)���)��ȡ(�����{Fҿ߽S#���*��ז�������
�G�����`��;|N���,#<��r��"cz�|��@��^"��Ƭ��SnBV��T��73>ws���ط���T>�������[ēUK�ˑ�#��5�F��*�+�u1T2�<Bc9�d*@ǄA�p�����B`Fgǘ�Ɣ��\&$�� G*���uRpI+V��Db1�Ј��He[�|�mz�]����sq�`)]���0+>��� Qv�@���e#��}���mhN�V󎚦�B�m2��!�2-Gİ0CDRS����j+�:�I`a��:	�����oh��m�����-4Z#�P:2r�x�=��&.�$�\��0���I�L��������Rjq��ǔ`����]��R����W��K�HL�����;���C����b�Mǅ��T�P
��d�UԀ�h��j����"$1�V�G[��a}��<&���d�� ��w�ۈ��d7���Y�s2�sS�Um=��� !$��U�c�W۹?T��U��c���n
x��h9k6)|�.�&�I
aB�!�e��듈m!�
B�Ii>{�"��@E�Nl�M�xEN�܈�R��wg;�RD�9�x>o\��3�
��@S�bّ���t� $����piyLq���P���<��r�=��'���Sy�h���/K�2���cNKR͢t�B�V�@+��E��w!�X����}
%�5����F�KP����雂�hո��)7VTڃ)Z�8���Z+@��/�?S�����m����.�a�M��rHsd��I}T�������${Oie��92B��V�~!���B).ĳ�b転��Ȕ�W��m"�tC�F��E���M縣Q0T_�b]��b�%�)��cL�����P�1��55|�c�Q��Ϋ�V6R�Tf<������{�'��æ��7t�ɱ��F|/z�FV�.�����Vi0v0��r|�pD��kL�����@G^�f3"�����j���T!�s�i8�FXA�67>#|�\.����h�y=w��ڈ�j<�#Շ���d�od+��r�rm~?-�1������R�_Q���k�4�䰫�!�YJq�k���u���&"�O!U����=�h�]5BM�J��h6�F��*_��7}����0�Tt�oلT�Zf�}z �t���=�2��|�٘��/N���	�b���N�P�,	r��p~��`1�B9�Py�};;@Q!�T�_���+��r��V0E ��-C���2��&�P|^�\�N��4_vM���z$�st7Y���xrL�4��,l�]Ey"�N�M�O�^{��ŗ���.�T�*�ǵu1�%s�ĸk+��$��Lg<���(��.a���TZ
�����f��W�gӾ���̾��]��k=-I�g	��ڱ5�IQ��]ش$�rum�O@�l���;�S+R2�_�@�@��R�����%���#۞����]8X(�nq/k�q2�	v�(��F]N�!W�sx�͵ot��.OHd�o0���4L�ղIV��#$;4�
7�|�i<d(&�"rt/�`�d�y㳴'y,w��h$ g��f�~�L���V���nz/����ܟ��u��.~���1`O�h=�-��^Ft(uM4���Oȶ,F �3�a>����♿E\�dr���ؠH�b�ط�^&,Ǳ��k��pt�y@4p�6[�r5VJ�:I�x�h���͙�a�ڠzmF�F��f��g������P^%&���1��$Pw�n�goܵ7B�r��y��|�\�$������U2E\���K��(@�u{b�7w6K�ٯ?��-~�̂iΕ}�׹&ҿi�VeaP�2�H��8�r�e���v!���Z+�O�W<�_�uӱȾ"�����V$��F'��jG\ȉX�P�X��va��a/K��(�^�oI�-��QP��D�2LH�H�"��PQ��lgE�6�;<���K�M}ۮ�5�����"1��qBٳ�v��8�2�g,j��8�W6���6�Dġ�����sq�g�,wz�-����O�bߓA�ɰ�����Z[9��_�N 1g�ږi�oܒe���+�Z�8s�Nf��B��F%�!������<��P�h5Wй���=�a
Mj��.<�r��"!ke���t�������ب�l�R�ܞ�E�\�`����_A�����OEZ��ح��t���^D�f1�W��U�Up����ē�Ъ�������:���̓����ˆ���b-W������M�ۈ/�9��֟�`F��k��S��d�A��&����7���xb��uF�����U���W���)��!�2�kht��@\�D��x�J�(Sn(���ͥb����eg�J��j��̀奲�YJ�
� ���0�VEk�R�����h�j�ib�x8��#��AOŠ�Xq�M v�O�T�Ke���`�78���
��"�h��$����z� ��A�H������G@�:��k�E��B^�q@�{o˭�U�Pٱ;�We�z5.B�cI��}�9�9'A���$������<�� ��)�ʨ8�	�v���E�����w܌�f���L��$��	y���W��IYdh1_�����ʺP-PM�v@�^:Y�����;�Xi���-�A���4���8M�_@8��?-���ŷ����Ҥr���2z?|��EG����A?��ωB��"�ju{s8�8�4\�|���SG ��N�	�1|׺�u�)��l��8742���I�i�9�hYTwS���W��o!���i�ͧ�'�9�y}�޵Yz�n�)�)�&�#��H�F	>p;�6u��o�d�B߻�0Z؞i�3rr���5���Y�h
�c\
��o)�^{���ج�w��W"K,b��ϒ�M��/&(ؿ|�M�Q_Ae�v��\��%��D�7�K����E�e	V�7bAq���zuEmԕ���+�.b<LA��'�k	C���� q�Ӂ�����u�G�KCz۫��|(h���� ����d"�� �
Y�����%��@+�g�Lȋ�.P�/jĀ1iӸ_��2,��ת��͑X�Γ�Ӝ*��[��0+;N�4��}������h�	��J2��ߪ�40jH_��][{��� ��b3��?P���
r+�����Us/5��7W\���4e�;�rwd�tݹk��5CFR/�F���h��Ā$��V;Cz�y�ז�1[��	�'k1��,���`w�N+��]�^6�.�pW����P��K�ɬ��Xd�=ʪ?������`�V�늛}귢��=_2�i3>*��u<9����MΓ�u�M�� �(�Yf���8�sN��HC�uF���|���V�ݼ�~S�{+���/
�E�C��ĝxd�-�Q�L��Q��} c(��%P`�y?�V��\lD=nK�?��P��65����[�R�e��f��x���U^�}G࡭�>U�H�d=5���#J��Y�}KLX�3��f���yv����+?��b���6k��ٲ�C�Ţ鱴;tU���&�-�����5��o?j�Ü����4��i���?�X��<e\�=����b+Pxn#�����M��@���N�"fP�"� �9��ԅ���x�ѕ��KY�,C��M���}�Y���oj����g���IMj؞;P,5>\�Rs���^����t�,|?<D�?����e9r���^��a��C�?�-n�#޴c&�HjW��S���q?K@4k�8k�Fؓ�s���5"�1���E2f=���X�S�'�@dy�<-��P��L��L#UD�%ô�ݓ����'�(���0�&�𽽜[�p����o����Y0O�����F���2�>/��eq�]��m+2�L��v �kQz�C��.�tP���*��s�1����`���l��&�#D��]^�r��W�c��8�H7�[9���ɽ�lb˲W��$i	'�J��7�N�;v�n��	�w�z�
�W?c�%�:�.���l>�iE�L����A��$��z�L�5%��L���X�����6>l���$�sL��8lG��E�o��E����U�z��k>lό�|�3��r��12ѯ8a��+$%����6�~{Q��8r#3�#��I�A��X�ap��M:7<9}�nR�\�����a�A�t&6f4�vT������E�E��!Im���ݳk`�|�F���c��l��"�$���'
��Q�cy�Ԉl�'�I�D9vf���ꊟs��.�S�U;��h�`ĳ۾BG�e����X�`�����~�7)��&^��H-��EZ|}c���K*Q��[na��Uo���#��7��⣼��w�p�AU�Ӎ�@c�M �f�JݓX1�^�]v�S��¤e	���-1	�D��˽�P�h����QW?m]L���KPu�v=��Z7N���IRt9B?WV�耺��1�6��D��Td�N�t���.&�0#{!����#������H�����S�L�Y��c���>B+JU!�048�QV�Ud:x��?ғ�2k�H��tģ���`��:3��C�q������3(�1���r6���g�Z���u���A�����+CFJn�y�@e�	�=
�O�Ϙ++�\壁[���{��daisxZ�L��%2l�.�sł��@��RA�{9?29�`�F�=��&Fd����+�.���q=y"�k����%����l6�J��/Ӟ
�����FI!���p�Z4nQ6�} �]txai`�+^��.���Xb���&�%Ck(x���j��&X~ii�"* {���]�[����<|�i��?8? ��П0\؉f��+�g8�g����(,D�b�PX���(�n�YCYp	.]�����ҁ��$���L���p#���R�ۏZ�댟Ѭv����m�,��4����$��PD�I��Tí�W_mu�a�._�Ynb�#P�� �� 	�~#J������Q�+�;��K@֢��.��#�,I	=A��/�@0��R�A"oұ��),��Ml��V��ę���<SFyZP2AP[��#������|�/�¶6�|A*�� k�t�8�`�F7��	���V5���Y"��Sթ�o�^Ǎ�P�t���~��"V	��4�0��HȮi.����N�����-�,�c���C�)���(���;=�V��o[��q��l9J����ftN�!��:�15-���s����N�K~L���D�(��L�z�况��{m�H�W(bPy�IW2�w�7��F��1��f5��*���4N�|���4�j4�t�,/\:�é���Ъ�T7���:�h5ĥM;���8
i_�J;+����"�n�2vvT�~�ID���AE�����z�<nP��vaztܸ�3�bc��À}I��I���d�}{��æ���$�����璯����Qt|U�VYJ>��L�¾�'ԍR�p
pt��V���а����$��:��w�����R���z�"����~����k��/���mFP���ϭ�A��cKjBՋ�]���$r��
@���}�\���2eݕ N�N��t"d���:*^D�ҸR>�h7��2�k�>�Xx͡Ja�S�,�����(��N:<��c�ZP'���������8�_��:�%8�e�t��`��č�1����9���tW �B�A�ҋ޴1{��׵%ߴdU�1�OAn^�^כ���+��4=bD\�;����oٛ���&+t�k��Ӵm�˴#�|��:~�<�Z���Z+G����J-���ۃ���VM���i)�E�JϷ�I�~`���.�qcŎUD��A� �aE;w��d �U5�Vr�V�Ou�k���.��+Y䎽9h�89%��HC�_K/%`���t���L�5n"�0�8�0����P:��b=���I���� �NYd0��f�G+���VDU�x��3��'#�ss�4�Щ�7Fֽv1.����.����>b��5�'M���;�����IF{�CE;��\9����ͤa���/��w��ж�~�?��g�
�YI#�lf��g����-ms�a>�dh�����aCA�󠈐#�e�
@U�T��R�藻Ӓ�{��?�<'�����Bi�_4�P#���N=�y�6��x���W�mZ��$��=���bC�+�|��'wlD�hU����(jPu���䧥�Jڇ���\��Gaw��"Kp�]����(���\����f���'���F]��b3�}�0�E�F�C�Կ2����/ꈬέ�$b@��C���mp� r�)�e]a5�8��|������vB��L�]H���	��^����䙤(��<���-��� 2�`��Kp$���#�_3N l�.7{Hh ����}T6��n��ަ[dQ�O����|H�䷹z"8��Lt|��#C��L��g&����b67-�]�8��[/|�ba�+���֍�3�~#4nXd�^Y��o���i"�ۑ�dS��4b'�C��1�b��Q�
��5�@\?����?#�?+�$a��_e���;�ɳ��g
�F~�n�s��������>R�XMj����$��-\�l돭�.�0�n��J��*�����}_ va����e��w��Q��)�O�N4�D��RbgO��&]>}���)xJ�Βs�xY�t�%��M������8�������������T�uCw4��u:R��n6��X#R�a�r�f�D�r��=��W)_�_[8
�x�٥���cS �E���I�	/q�I��+�KA��X���eY@�ƍ,{�:��z�ϩB�Z�lO�ed1��/Nt�� ���\�{@1ԛ����`�z�l�X�$���v�L����)��
#liH��W
X����H��]��.1m��*$��MH���i�>$`H0�Wԕ�F��\�m���.�u��KJ-P��F�>.KP�~a2�$���D�bR{ �$����<��k�qs����W��)o��4)g�烝��[ίL�-,�O|�\����;��3��5L�ë��%���ս��ӝ�I�p�у�	�g;�F�$�?�Q��w��(��1M���ͦa	�޿\'���ERo�Ὕa�#fyz��nn,�}�V:��IECf��/���?&~}��?�(vLDJ���Ws [���&5.��Q�Z�k�"r�<bO�ϼ�>I��:��� ��4A��01f�d0OL^4�)2<��w��E���_��
�46��u�".+$����l*�"��@���H����k�)�|5���\���ԕ�U͸���LiS�����oQ0M]>A0�O/S�B)'.�@��S��{�K .d ����:��e��@dԵ=kJH.��/�y���vK�2	��.��:�y٤F�3ѠL�*�yg6$����J{�"�Y��,[��1P"r����Z�����<s+<� "����y��Z�A�0���1%* �HY�)��߇�Z{��3;���l�(��3�SD���>����{�+_��t&{�0�t�k���ILr��|����YjPawvS��}]���!�e�i���Q#��a���v��g�j������?Ƙ�"�"`z1�Ź���iyZ-����sm����PӒܢ�ڡ��){y[Ul�Lwח^%o<ޠ�jGz��pSJC���]s�K�L����j��WwO�W�H9��D�k,���9�Y�\v����p=S�<x�1�?�:"�՛��.8�gd��ޡ��q�[�d����)96�
��@)����tl��Ս�h�2�F�>� N���Q!�)�u�G�!1:2q��*��#��(��q�kA;��&��S  �^c���A�Q���iB/Z���4D zŅ(��ƀW-�Zx�!����upA�`7��m��rra��d��}�0�����p�~�_S=���1Y��J�#6�]��9Ufݷp�Z:�\��$�o� w�Ty���`�{C|�j�P�n@_��6�^�g�>T.TZ\{���n}F�@�ߔl��7�FI�+�e�O�B�q;w�-�b��8럠�B�a�\�B��:Xg���a'v���N4sY��1c,�v���8q��84���Q�nq�&XU�X�i�7��#NoZ��QV�=�X��p���R��o�F�S*�o켗���d5�@�΀���ENԼ�&І�%#�O�9��@sA�����H��R����~8����6{�K`����+XFMx�X� �c�'�?��I<�?��sJ��Q
��io|��R��c���V���%ˡ����S;d �v˘[�#��[�$�8�J��)i}@���@����>6�wE�4q��c���81��c�Ĭ��䩍����0[�T���i�,��,����c"Of���&5�C(P	��x3�f�5_�:�a�3Ì��SF`�G��31�Iq�����9R!ΠO�K�$2<59(�|�^Ce�۩��dC�,N:X�D���7�<��.)��q醸�aJ�1��~��C>��ħQ�I��)1<�M���[�8�	6���Z��UGxN�%�d9 �(�e!�dR�K���¼�;3��?�Kj��9�EpCcb-MGc93ui�Y0��a������I��y���I����w�V=�*hƈ�M��{([|��d�yepm���CD�sf�3n4�-�{$��"��#�V��s���/�lw d�,�:�u)Ʊ A1:�[�_�T���V�����7�_��7˿G͒�q1���9��O���>UI���� ��m�\[")�"'�����[a�D����[��G7�����'���J�b���I(�ۃ>:��H); �)�����i�%h0��C�9��R���S�ta��h2�v�_a���E����ILj� �&:�-�?���>,�?��E��G��|�h&س`���f�0��m�����%��m�w�}m{nH�02h��)����<P�;ҟ�A�v��ɬJ�۵���<:ƎGz��r���ˢ����U����S������lG���gS\���>]Ա�P��E��1I�w��k��A�=�V�?���ῃN��˼������4��+W#��(��������&Lq��*�������y(��>�� >�5�NnPV�t)��Y[+P��j5pg��o�������x�zyǻ�gKڼ����g��T}��.�!����b����D�!W;TnLO�~+�+�Kb�IMb}����� �-OAZН��Ԇq!���s�CZ�zJ|���y�+�g�[ќ���.�e`!�X{�Qxk��Enqc:--�͸��fR�#q+���<I�"�u�߈�����=�aH?S֨*Q�Yp��s���� ��� @I-���[P�*)���OՒo<�r&�XKG�{�S�3�r,p��G{g�N"�2�j��X���4ܒ������'�v/��2��P�3n/I]~�Z�J:k\M*�\�C�臐(t���h:�N� e5��	`r%��/"r����Y�����q��u�Ni�α�Hj��6�	�������}v��} �`�*$���� t�,9�u*��MMj��E�1�z��� ��-=�k^����;>V�B�B^pS�X�K�A�Nr��֋&������]C-�u%0�>��<�H�r� '[�=Q�M��U〥@���� Ǉ�d�;�kc��}�J�t��C;5=���s3�y�#MY�Y�����]�64o�#(�C��.@<��ln���~F�:�!.B�9�~��vc�M�η���u��573{W�-��ǐ����;����q����7yנY:Jk1��k�E����?������S<#�/��O�RB���"�eь����0����p4$ny"��8/Ss5��+U�;��Ȕ,L�X��>��g��S�#�f����Ɔg���?,{�.���Q��=�)�p6� ]�@@��WG��nĲ���:r�W�l`�﬿Y��y���|l�b�yޓ`c8����d􍱅��"���4�
B��i�oᒉ������5��^&]+�Y �M���|p���t˞�j��:<��� ��\�Q����+�ˈ�s������i�$�Ѯ���R���.���-}鱹ۉ{�+�ZK��C+�~��
��僶ߘ���Wc�ՄdE��޵�����B��o"�o�'L_�Jh�@6�/�ə�;�+$�z]�Bb�}������-�����ӭ�t-�e���Ro �P����]�0�K�!��M9
�HYˉ�{[A4��ػ[7� 6/zV�a��`_�����d'9����p��,� Nt �t�:+.n,)��� $�{�)���y�zyZB|=o���ԁ��U��9�x���N&��Ņ8vn��"l��^"��s�$5 9�lZ����G&�F����{�q�̪�4#�������E��DP�y9�jIA�Z-\-�ȃ�ʵ>Hʸ�(�Q�ʘ�dG`h���)�Z�Ff2����o��}@~����R3�U� t�M�;�0�$����:�?	�Wȩ�K�T �}�����P������\�o�_�n�%� �ȁ��)a�r�˜�k%���^����)�k�4�'˝hj��$��&3ҧ�����!O�ѭ���@K�|jo�/��콀�P��L��[��2T�9���pwr(��t�[�6IB�Ǒr��|Z�kk4�8i�z+��������}@���tp� �Ӟma����4 � �;]��ݗ�����$�:���z�Y����#�ǳG3��GgH4i���"Ӿۏ��m�f\�49�����������;���U��3��z�
��� C=� '���A�I�u7*�r�p���dȪ��:�`5�5���""��Lދ_�_ܚ���.fe<�tf��ȹvIagK�I�ǵ�� ���X���:�m��/�b�����b`0J��C�5�&u4qe�X��Ys�:���wz)�Y}��P�{8Ղ�q[��Vc9,����ǰ:��Bv��,��K�e�v�����cPn��'�����)���,�ˍ��'���:�h,�sC���f�E�N.H���򣣎Ƀ�MG,`���7�����bTZwJ�H����&�كߖҡ�x���vD)x-�EyѲ0;g\�u'(��Q���d��
t�(
��l5BI�%�C^�/r��/�nȝg���[ԕ��=Z���Jy�B�eB��߬�q����[C )�j��@�{M�A����)R�����Q���}��o��g]9��;�f �-b���P{���h�OՓFSYJ�j5Q�7ژ��KS{ct�Ɂ��.8t�@ݪW�~�r��ߍ2�v��\�Lu�H��u�������O�9�j$hg���w�ӭ��~�'&>U�pǦaӏ�
3�'|�ь@A�P�@��˅�Db�����>d"���Tw�u��T��"�����/��B�CIT�ꋽp����U��)U���A���QP���*�b1`e�j@�ʴ���@7f����r�t�o�;��n��&�<>�mp3�n����$��^��9��)��B������A[x����D��p@Q���dI�CX �(�:��B�h*}mA���7�um5�J�<V��2ٍ��S��m���?��u�f�N��!����ԩq��=��IVB�8R���򒾮�|�M��&n��J?�ɵt1��ތ�FA?h�@����YU�6�:��e*7�1���a����J�}<�y�4*�z�d�ՑA�z�%���:K���n��>CFA�z܏/C_�8�n�JɁ���E0�)?u�;��E�Ѽ~�Ϙ`�q0���b�/x���g}���`��� J��^}�T���an���t�v�5K�-E�}�7g����>k���&���2������"嫟�RDFϝ�LF,ͱ�9`/,Һ4ҍ�߾�$��L>�����p���O���v5��s(�$2
u�w�/	,5���c[}LC`}We[�OtF8�(bS9��*db�M���ore����������:�Bfs��JW�^�l�B�E��'�[����D΄@��rt���dcF �lCe�̿^��>����d�����U�H�5�2��O��AP��c��8�������s��\9���@U�=��4���\]�����ml��[���ϽH���[��Cn
F3{!���o��';2���ݺ/�2��b ��hT��+-2W�.&e�G[r���F��eǤĭ��A��k��рN�4 ��l��k��vHL�](����"ެ8��!�Cc1Ï�<B��	�bncG��˜a@*�~�.�)��9�q��+#�j��T��$�m�-��
�qWեK[�C�re�.7��{+�'���0�I8�����7��˔��8~b2�|g.����{��*F>�C�!"A�6H�.��d��!�goe ��k��vl�������EO�^�̹�?���?b��oFq�tRx�m�kZ��Erq&�K�lk���3C��8<��Q�t�0b���7�D�����3R�,G�oV�B[�0����vF�_^D��f�V]+�xk8Y��F����R�[ mz$�#��g���tJ�����ut2�w��O-�k��ߞ���D=�3�f��Ռ�}HZ<FFV ah�D�E50�������Bzla�4�	�[�Ñgd~���|�q�_۠�(5��VbeT�0�oM6_�?�wH x�9D�E����iɓpOӌ���!����՞{~d���hL
�էp@-�Qs��,����;�؁��Q�U�ih�!n�eN��Qm�o9?C=�M����@��a}���A���1���YZ7�70?�&l�o�_�,[���ɓhw4暰v���u������ Z�i�7��vU�/���"�e���]��Ө�&C������ߑ�7T�����n>�N��Wo8 �3�Ҷ,�s�V�<ϖ�^0AO#��D���QS}e ��Ʉ2�?�<�<!
5�j;č���@��ʼL9��\�lw�^�`x��}#�����˱âEB-�BJx���K���è��4k>��8n��`V� ��>hrS����C'`����2^��(�h�O�HUZ�^����l�0.OH�����D��[L�a�)�&r���3��2��+��`d���Yy�X�`^қϗZYֈ��P�=!���Li7�%n��l�=7��>u���_mO[�r�t�eP�}�<۷�|DC��W�,�� tQ*�0����x�!�i @�c.)�S�:i_��=ͬ�[��x�HD�gNG;�ѐќ�0+�E9�虎S�%0ֹil�_1����#t8\!����-�����1��9����Ǖ�T����(c�kIy�nK*���λ�[�]K>��z1�|[�I����ɨ�����7� \ ���{��Ί���pTY{S�+�6����YJ�!�]N��)^}�w6�X:�� *J*�,@=���Z���}o�調��H�A�j3e��M��'��kjGT������L)2v`س|rw��;��(ѷ+�7f��([�$���Zl�6��L�*Y7@�^����hȵ�p�_��nI'ipfOZ�|]���Y���wq�4�(�=��˗��+M�d�jG�TǙ�WZg��.���r9����HU��x�,6E
�5o�ڊ��ա�p:�e�;��A}ɬ�x��f�e�JF��D P��oLxW+2�qŖ���l%�vEq���1��K.�8��2�N�~-@�\[��/z����(XtN&*r}k(B��l
w��>�KcCᨵ��sY��)�~ʹ��� �י��D��ۅ �)gס�������u�-aV���4t� ����?t���~+w�2��c���`�K����1'����54�U�:ƪ�7���:���M58��a�]�3���|�+[��:��^J��4ʧ�kY�4�*����V��ə�D���7���mvL�[@��Q�r�G�_����U\���<q�ٛ5˵WD� բ�����t��ݍx�a7�t){�_������#���L��IZ��H�f{X �:��n����Ϯ��Z'rL	, -ZqV���ՉQ��6�Ҥ�G��,R[�H|1��99<�3�r�`�M�_d���:�֬&G���#0ܸ�]�^�1� ���y]ˋ�S[�G��#�s��XϙD�uk�$>
s� �*,g�Q��%҆��p��Ă�뻬\��Fm��l��jC3�����kQf�c<uW;,���q���='I�f�T�-���y��8�����Ae�ķ��ԕ_ڑ�ﵑ�wc��x1r@a�������c4�c�J8�u����,5��u<hr}q�wU��8�� ѸxrfOz�0g*�8DGU�M�n�X�\�@�Y\ƙ+)�iPK�;�q�cd�t�?-�5�6.�v�T�ȉ�&��&���LƩ�r��[-(
4��@d6�yĈx+���g��4�ҡ����W�C���6濅h%������`P
Ƥȇd[o�,]-��z���cQD��NCߝ�����z|�ƤpHw�q��^O���"�@������	K��z�u�&Y���{���?�w�����hɧE���JB�����-2q=t�9aê8��?�.�����\�;�}V�|���l_�[�f �����XAӇ)&T��}��)�[Y�=ěl�� iY�~��Ղ܂?�Vʉ~����OJ��.eP�q~C�&�ݛ�<7l�%X���n�0{T9�!:i���J��_�	?���i+��Ub`f%7N[U��"�*�(�E���)����8�1�MX�٧k���lvOg���x�Ã,��/�FG�6�^Z}�x���nJ�osW���M�|�����d����su�
���&���0&�j������ʯ�YT��i�4Z�s�z���o�!=.���^b�D�:S�~}�����ݗ@K��vx����意x˦���o;�^G�u�x!����ug�KC���Mj5�(w9ڢI$j�d1�Q>�:�<B�Z��u�d�ŝ��/c
�Ǽ	.S���2�|���I��D�(]V�2����9zL�� ��������]HӶ�KP�'2f�K�����`���i����+��bq�00q�C�|���օ��_�k�8�l�uƏݔD�
d��W�!v�0A��m�ۀWd�;%2�ϐ��`6k��P�������`�c��=
K�qh�J) �Ŭ!Y�TEz�ݷ��(�5��Z9��,H��+G���~ڭ�_�i��Ǩ�f�Y(�ҵ�1B��O�X�Ē�5�N~�4 x��j���!�7<k&�B?��G!�]��8�6EA�gd�mD�Ԙ	�<!4ɊЧ5L�#�kYug��rj�(yaS�n%����8��������d�j��N\��J��t�g��I�����'�#3Q�G�6��4�#�<A(��;���ߐm���Ά#���Ϡ�7���.en+�	?��x�y�o���*��2�����&Rm�>d��m��-�u\Pʂ� �EZ`Dү�t4�q�uj�T9��P[���M�9zM���ϭ���/q��S�׵D��xI�,�?&��}�mQ�hX�'���� w9�~�%g��P0����>S�F��߹�]��V�!��FT݅[:�~	حP�lk�|�mf�h��W��0�/�=�t��Kgf��BЯ�����G0��:�!�1�/t�7�:�M�Lz�	]�eS�����󿳭d�Hx®2��_�#f��T��s��Iӄ���e�"xK{�!���u:�p�7WH�k�F�  g�;ڤ/��T��b�u�~�l*��qC�OSA{s��g�l�;�w�;9�;Fx@� uG�phR�����R�uMe�l���˴�W�>�5�������7D3�J�u9wq	��RTT9B�Tr���+P�@DZ���O� ���S�́��:�v7����|?�M_4)���KD���y+��_��La�S����g�E�F����q9(��Ҷ/My-@\�=v��5���GB�r��	>M.�O<|G����������^J�T<u��F��e�_+��qg/���i�m���(��k���٪68��Q�QL�9�+����q�:[�&d�����%��yZڤJAA��d�Y'����ħ�9l�k1��H��WM�������m;� �`9��D��J��o�|��+!��Mb�^��Ɨg�˕�R���Xpq�������#�O�X�V�i�:o�d���z>Q���F��b�3�Q��X�#!E��jRٿ�VS�+ֲ�L7�C���OĢ����D�V���)�l�m*��� �������j�ٞOI��)�r|�_�%��Ĭ��ruR=��[�>���S�$�"-o���D�8,�Q{	�qL�������	m7��Oq�(c%iH+�@�~�ާ?�=��+R����3;�I[�9�f̂�(ވm����
@���O��BRƗ���4�A��[��EI�m��{31S�l_�'�u?m���Kc�2��"��v{���`��Mˠ1
�	��ak!Gsɧ	 z�2Xś�~Z�ڦ�e].[B���pAڠ�e�ђ�ߞH�l��L��so
ڂ�íH���У��*p�;=��'��$p�d��3�q`��1�(�x�cFO�T��&plmD�) @�ê�X�/v�F���(Y����ڥV��������6kIi���n���Sx.�GF��li�ˇX�n���Z��˕Сc`&���RO�Ik
�@�*�x!��Wn�#	b:Y���@e��ֻLm}Q���-g���w-/�HI�?����}в���I��#�i��`Nc�a�C�Pz]�wi��hsњ����8�n�ގU���-��o(�q����4��`ir�w���)�� ��v*�.Z�/��҆�Ϛ�jM|�i�gx�����Q3�_|	Q��lNb�R��61�	�O;U���17�t�ռ=?�A�t����3zs��%������
6����#���PY��q@$˷��[bf�R��j��b�^GS�نzi��-XO�nT�]�I���E�6�Æ�O8T5�����|�U�,-O3FJT��H+ߦz[$��튬BB��T���>/�r��˶�<β��z����)C�?�����1SJ����W�?��_^�T�M�F���⋔���,�߭�{K�VS��/D�,@��e�.}]p>/�Q*]�Б!mv:������D��9�6|$� A�>6ߔ�Yj�$�>,�:�9����35���Q5��"��ù���Ѿ��pl���]�n�4�ƥ��/G��~WF���C���u;Fy�"wB	��c�.x�2S~Xp�|�3WT����.쾥n��X��[=Aqjd����V+��"���n�S!�ܕ�w2	��J��7IK�Շ�3�(&�}/�^'&�"-���Ʃv˫�
F�7�}%6�\�=�#��D�j_ �黩LT=
�a��tueS3W�)|Q���S�^B����jXA�v���Qa���'w6':��6��;��HO~�N���d�7Pڄ���)]ڐ�З��&�>�&��|�/E�b0��D��<�D�E�;8�.�@�IĘK�,�<Ϝ{{7Q< ���@�ܳ���^̢�w,��\�O�/��b�4#I����P�P���.��&�ѳ��SM��e�!E��	�Y:O�[!ҝa��?`�!q7�
:^5������"����(�1K'�9����*�s@�����[�<��^�h�Ď�&,��e9��t�fbWs�O=����G����P3�+��ľ�Eh�ƍ���oO�4��}��Დ�~�?d6�3�l7��'KJs���.0�*ŷ��ʦ�~��"(�\@���W&{�l$�Ȟ���2���$���e��91Ox��QG���Y�w����&H��2���I��,���yg���a��AD����R���D�u¨4���d��1�� 1D[j���Ap���_���6��\�6�K�<�۸����W��c�d���$J L��n��ˈ���^�k�J��6+�;�ҭ|2�m�p{,�C��4Uq�G����ȿ�%3vj9���Zۏ��3)�����c�Ye`���xs��'x��;4��c�&'M���{��w�.n:�{�F���m�7�4���^e�N����&F�qۇ���e�.���Z��k��A��?5�C(�8��D7ǿ��2�j�{Q����_�����27�E(���u�5y#$nTX�zvZs<����ouL����������"�i�`f@���5Q�B� �Tx��jٮ�u2���uFV���z:oM��5��=�!M!X�2O"�'��}��1�A��h���B��C��u̿�L��p��(���paȯ{W��/Ŕ��]�X4+��A2F�p?UJ������я����p%;̀���*��{�x�_��}dh �JLFB�>S�Q�+8O5�}��n��
d���s�N�*ZPl3Z�2�2��'��,Ӓ�_C
�9G �]���wyy��]`�M�*�-����/K�2�.堆� �� <d�[���B���%�q�F�����F��>�F	�%�t��J�&Z$0������}HVM������V�rMZ׻�tR���A�Yz��-�Ay�����ξj�u^�Ό5����f��"!?q�-�^���8�	x�t���u���pũh9O�B�_�0$��᣻�I�Y���HP�_N��?�仳p綳��4�gE�D�`��y7��6�N��j�e�����~���.�����c��h2��V��8��.Q=���Z	�oW4�߿��{�F�F��oR"7=���
�NϮO���A4ҽ<"0�L���
�ٷS������7}:K7`>�F���)@p��h;�^���NA������#�3�r�l��-�n�#�J'w:�K9�M���^B_|�rfe�®8o=M�u?_d�(�"vo �Fl&�t� n���N~�����([lLd�ӁM9���*x����rE�˕����B���γ���`@ �ɥL�ٰP:��R�;>��B��,ypH7��T�-^Ou)
U���n=H��{^��Kꊣ:��-Y�94�~	b*�d��6��_��n��������MY��X"��P�?�t�{��}!���Z�R��lc}���j��̃�I9(��O�W\
p=_���<B�+���N�@(3�E����iܽ��*1 �TY|��1��\������,!]���N�j(#���ԋim7J"��@`��'3}���=�X�785A��/� ���F�K��_�2z$�T͇�7�ǰw��]�U�?_p�=� L�5���5}!V�L\)hG�I3ѧ�N�8���Ǩ{W��g;b`4`��Z�Kw�{��e�x^��VT3x��bue#���{�]�H����3�΍���͆[{�%~nm�DzS��!̍�-dC)j��aq���M]��������)�-P�T�4�hh��.H,�_�M��oׇ*�d����0I�i∩�6���-6�I:�+�����z��n����m�E��-@7,ct����=�r������ބ�EW�|��LS](HS'"ɓJ'̀C��ݯ�DY���aE1" ��L�IL5��;��2�d
��TXſ1�s�¢v�����ӫbc�����	�eTA�����^��c�����w�S�����F��;b��=�fޠE���ۑ��j�d�oХ��4͠
�{W+��N�����I���?	}�"Sfe�-����ưz({K�^73���ȡF��"g^,XX��Fz.IӠz�K�����g�|M#��%͌gGH�Z䩈H�˝,�e�ӏn����6�:=�Y���~����H�H�'|�v�� (���3�Nϓ'/�''����E��c�
�P��71��Z�s�Dr	�^�ln�Fj*��	�B0��ա0��H�2�C2���ܩ�2�Fμ��<U�ݨ���tQ�T����}�m�1���F\���
F����1��q�(�ۊ����!��ɾ/i*�	�~�Y��\`�)�����[I�Hy�1)�a�;cS�i�bq<yr�!�Om�u$�.��+���a���i�wRJ0�6�+aN��V������Y���޺�����X)�}I9Y��N	�<�"�Oj��`Q��7/ͣ��L�9 �[�3/�l�"����r 0t��p�c��ƖMŗ˭��� �R��4�2H��K���'U{eNH!��X�aиZ_@S`�Ӈ#;`�2��bI�m;�~��TL 
�ɰ�"�`4�΋�T�Z �@�G������uym�tBF��T������;R0|�|�/=`�I���i>��;u�hF#�{���v��	eݕ0E��fE�?�<��k�vªkեA��v�Ϡx�#�H�l�[4@�?g��l���M�˫��(	�H�4�`E��F~H���~���~2���9q�A��d������cܬ&#��:�W����A�FR�I�d4�
�(pGtƑg
K��d�z���]j`���<�!�	��9�Sm���Kš{�����)*`��F*�\jY��0Q	�P�؃�6�ڝ`a�����
x�ɠ
��9���7U���z�W���_X�<>I�)�/S�T���@򴔩@Os?M�c�&Hi�TpK�4�V#���W��HWɝ{�x���{� �����~k�zC�S���^m�/�GR��'G��8�D���̽�I��t����-r���QyK�E�{�|(�7nSz|~*��O7d;!�RG�����L�� �	X�f���[jC�l�����v�?#��+�`���%^���L����\�ͅ��"��U e�HZN�T�]�KmG�h��)�U(��x���x'�8!�H9��%�!�r4h,��";
ǐf���Wv?���qAtq�FX�w�U�}`�X��/v	X
�Ö-�ea�I~�r���R�(�`>,mOy�1�%sw4�)�ZÓ��)Sɤ�mW�܊�7���z�L���p�U�8 b��9���=��8����X���핡�L���-�G`�S�g��V�.��UY��e�!f�#�P	:�n"gӠH��>S�9LI��B�P'o�h�;���'%�n�-�j#�����,R7K��-34O��v4S�BH5��j�_�HƑ2�8b�C~��@Z%J�D�P�bp��3��[����u�E2"� Kd(��Ks�կb�|E>��}�Mۀ���+ﴯ�^op�#�kZi�G�{���a*"I{ 5�}�m��b��i�`��4V��Mޗ~C�[,(�W�>I�#AisZB�(㕘'S��rb\F�|����b?$ׁ�(L�EYtL�,$�6[XQ��K��o�1�!���Hz�C�L���J7�|W>#\�M0=��k�훀�FT�����E�bԄ�()1%�����ʰaAw8��d����(	�.�3	����N&����Jh��w(�,���k����������U|���q�
cMD�V�4�iǺi�l��WF�5 ����2F��{��C7�d��V�i�U���%���Z�PT��C��J�3^~lXnX�"���L�P�jD ��{���Df@9V��ﺻ����P)��iVˣ���������ֶ���jWy����_�7�&Ĥ"@iZi�]%�Յ����y�A>|�-�6fN��'�kk2�S���<a�a�݄�& ���� U�U�Q2�K�
���o�T�q4*7�4�EѢm}�ޣ���UG��R�6H��-;��\ͷ�4m��K�qyʌ�8�%i�M� �pU��&��*�2�)��էW<��g���O�"����R�9�s�
���QXP�CH��;v3.�/_����']/U9��:QG��[?���L����ؚ	�w��_�;� �HU�UXV��r=+��6�1î:Bd�����&�d�yO:NsZ��z��%�f3w�I�k��T�v>1w#��0����� ��7ɪ6H��ȡ���(jy^�����yr�����������r(P�WWϤz�/��Tg�ۍ�J���;�����P���G��m�X�5���D�dv.�F��E�2F!��fN'�L5\�wǴ����uW�_�'ݣ�r,���m<����fL��i7ָ���W�(,�t��0Hyv��AyM t���]ˉ�U�EO�k��M���ur� ���q�g���[�oM�K�d���t~냟����O]T�{ǧ1�Ȋ�O!�t��-�ؗV�q�NT�+b�6�Y�d(�`�������X��v7�������s_l�H�H�k~��#�=�[�*\?m3��3�6�G&[q��'�+
���t�c��_e4�S��F�tUA�o�\ڶe�, %e����:R:�+�1�챐�˯�
Z�/*p+P-&��#l7���J�vq��X@����9]>@��B�W�V�@<��N%��U}���T��ڒ�M��L�$��X�*E^Gx�Um5�w�k�?��}��ͱ�z�gY�y��ڽ<����&�����L�����E�!�%�����XW���-�p��iu��2ǆ}�����,t���>4�(7�o���-��oK���Ƭ]X����?Z.!`k�Ɯ��dR�\���'�[N��+���M[1��<�z3���B�]���Y����j�%Wi��4O0���g/������� ��-p�B�O�T@�{�ϓ��
����W�.���]��(����dU�����2��,����Eu�N��4���8Ekgׅ���鑤7��GZ3Dڈتd��$�4�jU+��]�K�M�5\�q��1��Y������ګ5��cO�B+��C��(���?.4�	,�T������O�:9���A���9X(e�J�(tZuFGM�Wu�/*6̈�lo`O�z�qa�l9��L}b��h��b����!J���F�_�@��*��N��+���.S���,~@�@�k�k@o�t�V|�&�/��Z�7��^?Z��G=(@t��B�H��u�(��:�F�:y�^��Χ#�U]�Kga!��m̕����/��!C��!��� � �?6	 �/��O�>��-P�j�����~2p���&+�Wu���#�z�ݮ�@��I�� !X�y������|��8�0XH�9qѪ:#��CGS�~�0q�!�RҠ��S�y�"b��
�O~��?�M���܀��ܲ�`�׈�Yd5D_j�E.��2�LHo"���ڴ�nU�t���EĤn��B�֦�|pi�v�eT�ۀ���=>ݗ�+�����dX�Vx���zs��,�N�v#V�)���x3ǎ�]�-;ӯ	0�Bᝂ�A͓)��i}MJ��Ն��^zVĤ�:ZL�_7G��]b��VvΓ?!�\��V""�g���aW͗�-���1�$�g�?���#إ�- �1ɢ}�ݥ/#fi�m�R'員�i��RF�G��|m;�K{�˾~�6�-Hzy[R�^��Q�j Q���HJ�g硭a-�\h����|����X>׵$���a��9�'UV�#ֵ�(��z�Kۚ�&�E�Yk2B~'K�/����Q��< ,a�. ���Gt�cc2��T3!��j�G�Z���}�r��(K��k����V�<�)*��(�Q=��@�W͉�P�W����bq�����`��a�
Wn���rkp�����3���A�p���Q�K(��c)�ӆq�*%����}��I�*�z���s�r1����#"T0�O���c�K�hL"��'n��'��Y�g�ɰ7[��#"Q�;9���q�-��/p��V�B"�����MS|���Ol�F8�Y͵�G�J���-
1�$�M�r�N����r�O�u��I�^��N�h!hH������.@Qq ��ԝt�o��!�t5Y|@i0I���c�R���7.1M�����n�e�>��r������5�o�>7f�l;!~1��1㲨@<D�Ԏ����Y���y��&ͣ_$4�G�4簤X�
0p�-�A(s@¨i�[��8{���@�
>�9��	#6�!ht�}M�z����(ûq�1�z_o2#�����l��=����y����L�~�6E���˺E���LĦ\	�W�/�z>�����F�Qk�8�;|�.�H*K?}�q�{�ذB�&�& ��������O`�=tˮ��V88p�?e ���n#J��O�+��,̶�H�1]�,rUF胾�;��%�ן�
@�A������ gQ:���'����U�^�vK��$�_���"�B�s c	�dY�Џ�g�nr��I���ʫ���iΕ���)�#�9SSF��\����ܗG��^j|Da�3�޴�g�G�_s77�bR)핡�`&����[�R=�(����X���V�ϑ�H�4b��Mbu��Q���r�"� [G�n��QvSU^>ڑ��'�qu���xB#�u��Y|�~����o��C���vpJ0f݁��~������𳑕 ȥ�t��:���/��0{g�I=���"�#�mp�V���Q�8�k���2�U�T�Ū�!C:�0*�I��x�6|��,���]?S$��o�+}�n��^����?�z*��RK�"7 \�[z���D7Z
��D���	��G6}�q@.��,�d����P_�f+�$K{��aT�9��%��6b����R�� ]��_$5�	��\OV���Z=L�;��N���!l2xDOR3�
}���/�;p��#�v��P�n�4�l��fc�wh�u��1�9IL�`GܬVz��Yg3Z�J ��~ޟ9�^<H���r�f}��pD	��j�!��z��8H�[��C�=��X�8�w�9���~@��@��u���v�373�C��n�$����OP��Lzw/�W��-��'����Z2��#�58�[l�@A�v�ڹ��a�_�g~v��t��g�_��a�%��1ä�@2�°*�6�񠽥V�B�ǯh���1����,�:$(��l���ѿ��@��1N"�#���b�/�܍�,c�lW�,U�-��>@�`��jʯW7��7�P��s�{�Ӱ��s�^�3���g
	4��Jغ��?�]���ن�<�Y1�V4��x|ⴌx������WB�ƀ`Y4��l}�����#��6���#: �e��A�g:R=wH�7)!�[b��3���5x����M�%�V}8�~���C�\W������C
ʀ@H��:�f.����

���J�y-AU�H�U �s�A�����>Ms��V�ΩD�Mbޢ���K��E���t�K��7a��i�3�'���`����r��1C/����%<��Y|����пE�R逭C:� C��|�q��TZ�ϥ2B=�Jm�~�vW��a;���u���<d�I�wV�ZWJO����"�b�'f9��`�$��d��O�����|�~�����_����QL�7�Mr;�@ 5�o�{�i噦k�J�����4=��`�Ye^V����TH ��.���Y<b�@�"�z��^��"O���=��w/ ��:wzV��4S$f�PZ2��[��9X��י�_P�E��#\|��b����L�~w�ݨ!Q�-��R$�HzBV@�u��Ѥd��E��ج�r!+�n�-�n
�g�X�
=���d4 �+�?ޚ��P}�#D!��b����5T
���o�txxZ�����HUQ��F ��������"@@Z1���@l������2����(o�]f�:�n�\��J����u�;��-�n��ȦtJ.sh� �{sd	���_�V�.Ws�����y'
م(g-H�5�,�qՆ/�+ڗ �ϻO��)n`Mzj���G�P���M�����t3>T�m��a¦�e=���V��5���q�`��`�B�:s吴9� ���_ry#ƍ��&:0���P�;j���>O����+T���h���!^`8�]PT��k}#�ff5�1��`$z9�WY��}���g^o���@f�Uc���w>��I*)!XR|�ᕘ�AtLeE���q�������A�<3B���G?�L���x���𙹱����|��4#�[�@F���f���u�>j�뷌��<�C��0�C}����j'�ݟ6lN�b�"���K� ����d�tܯ(0����R�\�H!�5{��@o;{�d��x*��G; R�F�-��S��aDc?�Vz�鬣�5��ܓc�=,p�?�K6�@,m���:�4m�+Gv���+Ε����$y�9{~?}���a��N`�~�"��o���Ϸ�5�1�
�*�g�p����W��%ۊ���S�q],j>�b��Bl�,���^�J?�f%�5Εi�U�mdUI3q{���W��h=�<���_��L�f-������\��`>G��K������+�)�5v/E��>quPy(Z�b�Nam;Z^��umf/�t��[���R�-�����)+A4�'j�� L�G�bt����HϺ�Ɍ�߄%��KW��5֜uV|���4�aT����PC�J���ep&\�:��Bm(H�P�	cߍx�;�h�/�u��ĵ�_4J�Ё2ej�"�j8�7{*��]�H�5���}���0b�Ԓ�"�`�����h+�X����$�?����MT�:Ri�V��^o!��8�jX���x>U��a��!�&t�nߪyL����{��p��n�*U�@CD���SX��w��V�Y[�#Tt�i��r��F�]+�c��~E�͒ǘ�ܑe��x�������Vgwۻm@��y73��˱;l$s����0j��T�)���7�a����Eyڒə�.��M�6�&R��'��U�p�zZ�=�d��߫�7�G;�!(Quw=CO�:�� ?���o3��{�w�r�X�����W�~?1�+۟�=�被���d�˙�8�ݜ­����fu��1���w�O���L�vx;�K� ο��%�I��M��x�z����m�v؝���x6w8
@+��Kȇz�JȞ&W�aA�k`���HA�O�� <v�C�#��V�[����ާ���`<#𴞁���⒕�Tԣ�,��bkߖ�'?~�s �ƌ��7��O�L���nuqkZ����m�̳�j�"�ō����0: �GX��qӔ�q9f$�NMi��A6G0�g����`�� �骕��u��Ң�py?�lԓ��V6L!Ѩd�W�����~��5�V]\B 	����~�c	HK�D\S��{��	>�+w�KI���/y���k�ʹ��M�O�]%�J`����LeUozJ��ZƘ��2��ōS�D��n�֝x�튢�}��m��zT�~w|;���a� �<����^�/�=�&��b��0=�ϭz�hd����c�,��7+O��?Sr��R���!kP����y�	P9	>�ך����?"OWtW��yb^�dH:q��Hu����de���[:�`�i%�ʌd9�Z��˂�[�7�z�G�*�7��Ci�%cV3���?�Y1z�Y����
,$ml�VA܋)z,�H�cM�w1�����[��h�B���X�r`Y�͑�'s����$�fGD�-��OE�w���礌��XjH�C��e��>�V�f25��_�ś�� 0���{���;Kܜ'��O��D0#�c����#E"�^{	���hoͷ�zA@�ȗ@��g�r!�5�9d�s��

�8�O�T, �bS�>��X�f)�������^��dp�pa�:h:��BP���2'���_|�U��$G��@��ޭu6�&���c��Y:I��v��tw���΁��������е�^߯��fJ�pBG+�m��x+���xr�N���-fl�=b����5���O�1>�b�g���<��t��ϭx/|*��븪�,}�y��z:��N�X���������K9k��My(
���dߟ^s���Q:�h�Է��ơ@�5��hM"��N�(�w�|\.�Щ�T��1O�*�;�ƭ� ��z��fN���Fx��ZZe��Q�d����]�����i8'�Z��T�P�+�Il��1D�!Lԭ`��FnL�@8A�`� ŝ��'�0~�*8���}�1�����=���v]{��!�sژ
�$�e�1"����!Pv����pr�Tx�X`���q�����5���!��]�A��$���1����8�qj�-PŸ����ol�.�m���1�@VE�$B>8#���F�c���.מX�s4�W/���{l����]7ͺ�Q�w�9c�YPG�6^�LH3,s���x��+�19v��<�����V)���@+6���j8!���ڛ���%:�
ߠ�+��xe;�W��J�U.ه|:b�;tFfG#�����	d���9z�7��X����3T򻥕�� �Yz�X<�a�ŐD�
|F�p����� j�8�Y���^뫎��A��7Z<x�W��;�bp�,I�2�6�%%��D�2yď.H;�W�4 �n���0UK�i�D^�1H�>7��`/8S͒�tO?K�.�}	���_��x�:�ug��R,�x�=e@ݙ����I�r��X��0H�p��{��|�v�8w�S&�g�/�ǚ����>?"�6��f�T�"�Ȥ/��΢f�������S���\�?��O�7���d�R:8[X6]~�I^��@�y�X��3�
z*�Ti3�WF/�x��<�*��h-������u*۸i��P����i~��n�����f�׸�8�Fx}7.�L���g����-���>K��y�_w�,��x3��"]��AFL+EI��t�0V5��@(%
VdJD��Zt���I��q,#�95��&���	Y	��w�����܎�v�]0�/�I���:z)�U��[^�'��c����pB�5�%�w���ެ5PYudS@�q�B�Q�c�qc��ɦR+ОVtJ$�ߌ	2�$:y�1.�Oضi��AEzF�R���9?�Yo�w����>���v��V6�2e�_J"����dA�^�� ���J�O���\0��Z�G�C�p�n������	�<b�?!�}$|98��N@�F�߭�K�@Ju�69�jQs_��[�XF^����Y�>���`�X����m�u�o�v4������V�)��䲺W�G�������Y�j?ME��B�H� p9���'S�S����7]�v�/��\���"8��n+⹐ui��o�&�Ҧ�����[��v�Ŏ4n�맰�Q���QG�`�Wv��w:����T��U ��ϥ�7�+�}�i��;�1�H^V�;*�0 A�;D#���t��YV!�Y�9� �ҥ([�	���Y��� !,�;�T:P��Eϖmf��T0���r�zK˞��qC���[�l��օ��Orq�F��R�+����w�]�lB/f�sI�W�q��r ,eU�����iG�m%Z��:i��}�8�\�خ�<�UȲJ0�;Nd���\��������|"�(�E'7B�U�p�M��J����N*�*{)�(�1�������7�9��z�� �ij�4d��Eޫ`@Hs��<)���h��1��0AESZBٱ��d* 7�M%.�WBe?�A���(�o��>h4c������S;=��]�l5���k��&X�_������"��j֑Sd��*��F���|��{���h������벊O�X��?t�T����א�AK
�J�.�mgP�Ѕ�1��4�1QS�8��!i�M�G7O�Ї����76�;w�8�Sç�e�b|	����J/�V�[�
O�)bϫxP�)�����,���ʄ��ρ�YQ���z��<lwP�`dq��l2 ���5�&+Ȓ��p��*�������W?]Q�4I��T��8�J�@��f���O�J���~��W1Ry��ko�e�
5��d&�76I���I$���;�� խE+o<�L�� �u������^'7�R}�<Q�]�<���§AÒ�2�ǰ��4^�  ���1�"q<�_"�c�}h
���H�:�������+��ϴ�A��2V�|����E����d{T%37�@�/T��&_�'�~��B��{<�t�������I�`�W���6�k��#�]����u�)+`z�Eo���%|B+�;�$3�`Vr�
����Ң���D]5��*��:�7[%�r)e������V�/݁[�C{��-�=�}{TP����01	~u{�W���2�"�1���_����ɷ7�E���d^��q�)М+���\"����#����X��9k�2쁜̇.Q&���Ox�d� !A�v~��ÉO�`���	lp���ܡ1�(e��H���)���S�nW�0����$n⍠��*�7o/��n�Ee�/�7�y��Pr�N�"���2��;{��7���s����13{��x��J}r'�
���w.�7���;��۬���c|x�xF%D�k�mf�֯�����HH��ahѕ���"ζ������&�H*{��fǰ�`i�y�W)�Kd��$�A�����9�m�u�_I#��`5
�")��B��T�x����%��nx��#�t��
�L'&..MkM`3;�p<V��<��k���+�X��lb7�đ}J�s�{�9:�Jվ��+�j�:���������Z��i��F��s�>��6��hx�?B�r�	��e���$Dy��w�1����no��#�&V!�岐�vE��/6��QlW&й�|��)��U�1Íc��A�$�pW����L��ߙ���{�_d�Z�ِ��|H��b�K3k")�[��61#�f0%�[qr�k�5n������1��G��櫇�9�Ǣ�]AҌݓ(��.��o͉+�Mm�.�p� *ݟD�Y���"yߏhé��Ʌ��-yB����T��j��w�w _M����k�u=b�$��n y�N
�Խ���C�8�ԐY�aX��Z��c��������<hjڬ�&�ގ�)�ￂlT5�X��ԟ���{o|zX:m��m0[U�h���:i�����̈f����z䣭�\�&���E�v�ۖ�j���|�1�5RC�1�>W4�k���7���H���}w�^�̔0ޤ��	c���@Ё��Kz6�7�� �~9V` ����8�d�*���xp��jA��l{�۳�[����>"��q@��q�Z���L��\NfU����ZY-���;pO����F��r����KnpO��8Q��y��7��Ϻ��˚�����_=}"8f�smHuGf��B☶�d�*}��l�����ѱ��Z�[>s+�GN����������\��Z��,Ǧ�W�)W��<�r�d�J_^�2F�z��R�$��$�y�g�]}�����h�T�վ�Q%jsV��x���k��+�}�vX��4�"Zi�m~Ui�^�4�������-[����sg�aP됮Ac٦����LH���Tf��3Dn�86���u��v��E���!����*�9��R:�dQ^Wv*5%�1��E���R��cp�/��7�i����6�V�Z��:L8�G:��Y]��(R Sg�];���M��#��ɈM��g�k ����۟~L�*QD�K�Q䁰��4�i�j1K��gg�*�4a���:9��H���YM�C �����݃�ob̆Ӛ"�+!�t��L�!���i���¼�Zq(ϿE2U&}�%]�3����g�QMƾ�%":ʯ���a�5��뙤o1�����71J��Q�':!h��}�v�߄��Y	�0;��L~���Y(��e�0�ߔ��K�윎C�zKk��$�B�S�R�}��</�O{�'������8�~b"�����bH�2|��?�;�i�K�40Ul�:���DP'�0�B���`�VS-���>�1#��?K��˹����gNp���SAj��I�c@GS��!`'qR�m�e���w�&�׽�c8�Y�T$T�+����~���=���}�aVr�D��ʚ���-��,����aV��F��؂`��&�eo�M�'&o��3Y�n1���Ӹx�[7���Y�,������,v��Ԯ��>`�?�Cq���Y4Z��	���q����f֊̑k(㵿�:��<	h������h��
��7!0�q(3?XGa	����nOi6��/$�y��L�w-��9���� 4��w�L �o�빡��r�y���h��kiw�G0�����m���!/S�Ҫ*�a���c�]���|=y�c��_B_�S��'we�"�R��&/����ޕ�N.�LroM]�-g��-��v�K�IdkPDS���%�}�7\�a�.T�&�]�ĩ'IOIw�ш�4�4m�z��l�T��0zp��>���=[D�`�'3=#����2%���-�2��Tq.c#!���@[Xg^JX=�� PNtD�r�?�X� ���Y���F����׳X.A�%�ȇ�{�c'$`�;����c2�=�~�Ň��%�_l!��a����4�T�������E�$��D���w��Y�W���'��w��&h>x�Jht��� ��ɵ��ܠ����#��>�[��B�|B�*�fi�LH��͵2�k���h�˨ �o�˦.�_���6ɍ%�\N=��^EĉZ��r�S���;�@��WY]_s����Ra��Mi�[�l���|_s�R[����S��!��4|`�N:��k��THS��@�'�)�ڏ�n�W/9C�l2��@
�dw\W�w q]���e�4��'u�H��6�N�L��իh�	|�nc�=!���	��A����ک�}C8'�-4���g��s���� �7I\�<{wu����֍��?�oV������ޛ]�H�ѻI���I5���v5ʝD����gޥ���~�S	�΅f���$1���ހ�X������d ��$t���R]�����W�1-��\��uA`�Eٯ KIoʓ9q4Xv�]Xt�0d)���#]�)�;	��y�SV{�Pz)��h� �����~�[����"j�uv�"�B�?�P�J>����`�㡧PcE>���o{[�3o�U<�ʥ����\'�s��jhW�5�M�iN��9@{jo�c<��O3�rd�B�:�I�����+[M�=�_�mKo���/�Ψ�K�o�i�t��dR~h�a�4)P���W�^c��YN������I[����z/(��@���B�Wq
�y�sbS?]Yp���q~{y���{յ}��ZE�Mz����`6���iFCz��T!ݫA���Qg=��v]~��-�"B��[�|����g0�s�~��p������|
v��G�DSu�$n6���r'�E�m!d��[Mݺ�+F��J�.!��Z�M#�(�:�n:�8_� ς����	=?WHS�@��Ԭˀ=��-$��a��4�d]���d�>���g�D�:*G�Uߞ`�:�7rz��s@���C N����~I%�c�$W��£�n�ӏ�y�F�V��㹷�����pDq�b��Ʋ�Et2�n-~i�kw��|�����+�G�''iJ�wg4.a�w4P�;��K����0�V���	p������� Կ�Y�D�Q��S��������(�����tji�Y]��f���O#WgB������y�n��ư(w��T��e���4��J��Ǜ�ia���tZ7���6�ח���;s�UQ��)��cm/�J^O��7���E.�pL���Id�	S�*�HU�Y��	_��n<7���xī�.�h=J�g8Ţb��)�@J�Vp9���y���s�&n�����a�'u[[�)}��O�o̭����#;���@'���(NU��	rB�!�=��-D$�(y��Olm]�t������D��öKU�nsB��5�,��N���Y�PxN}�>O��Z9N�e��i�c�]iY�>�zc*H�7�w/W����;�6��.L�4������7Y+·|y"�SE����U��O�Ci�ÕcZP���,#���
��UDh�#5_8P?ӭ }� �q��5!Ŋ��I�ޫ"b[9���<d���h�]�2�X��,�tp���L������z$Z�G�Ǭ�z�f��W�����<�\�mN���ؘ �ǎ^3�Uڎl{P\�J$��? �٠]�C�D�=I���Q5o���R�����L@�_y5`�N!gi�9�
T]j ~�����r~V���Cն��̚&P���Y$Z�Yd%��a�HKbvrΐ��XL�G��E[��U1,�;%�'����zrU�D�z_���٬��e��|� 	)�&M�c���m�اN�Ų�`���t�k�ero|���޴��:��η#Eخ	�\ާH3�{@���a�]��vWwt���KL/��߅1zuR��1��J�@�F8̬�p���DT���	%7\���mU �K����C~�n��FL#�u��=���u��n���K/�25� 0$T W|��G�L��AOA�������H�޽N��p�L�v�^��VnKm���b
�zż�Wm��y���LV�rw�N?�̱v�i���i`�N�"y����:p�8�� �pK�84c��8�Q���I���J�$����	�!Vp3�>��9�qO*�c�]�^����3C?�(M�4]�Sd#���2�{��,�B!�N�n�#jvT�Z%�9C��QI�N{�� ����{�@`���oR���,0��|�r�V���
��r���I��p���;��k�J����$Ð��%����L�Cw쀪r*W� �c�^1��ԎP��+�A�玥�3�P�s�o܅�W�jJ}�ek3�8���E��x��	v;��Y#����i�7O�?�X (�t���p��;a;_�z�h���F#mJ��1�&V�~K3#�t���|eqO�� +d�Y��<"�a}��<�0�"��{&l���,(lcWC�-����٘����ꀏ���i�ט��I�9��Njg@���z������,�t���E���PQ�;��P7�C@̠�>��ni���n����@�N"�c3HN�8@�ܩ�2�=���=#(�ðF�D�jY������F��=�@ig#v�_�*��r���;�v�G��:CL���b�Tj<Kf�D�Oz���R��<���ɷL�W��m>�f��S�h>�{��GU�^0���s�D���a����T.�1}�8^H���@�(�o�'6���B�U�q���)�!c�s��2�����vRވ�$+b�� �!y���d{�T(AQ�n���y�	rܟs�7O&�J+�kj��m�
5ю�>�C�b���]g�Y��s3�.v Z��JSkh��M��$8��l<O�_�x��ip~���I��~스�x���H,��j\��V��{x��>Z��&}Ǻ@q�I��fC�h��<e`jD���p�q���M��Ui���_�&�=4�u9N9���j�B�-Ǎ�ޥF��,��6R�>��X����JVp-��+��aZ��s�l��������:?�\*7TqBFk�$>E�o���8~%�0r�'�d=�S� ɽ�r̳D��xovN�$z����\s�S�����5���ȩi^w!�s��� e���rc��!��~J,�kZ5��	q�
�w�lLˇ�'��T}�W�iB��ұO,��W*)�a�_.O���΋u_y~cQEs!K�֠�*���U�h$_@y�܇�����VŢ�6� �*X�.�"�T�5
)�q�C��ƽf�+"ι�wG�����E�j����Q��i* �K��v�x��<�7�{_oR�N����צ�қ��mM^G��aDf�Q�����z�A�g�R>a	A��RHwt��$�ռQ]]������`���%T�ι�O�[s|N�){L�lE�)|f9Q���=?�	�qT�&����7�=���vϑ9x�(5�>ZL���|�a� i��mk�n�̿Bj�m�eYۛǚ�j�]�8Ҡ0�
�Z�h6����b�����=�"6:��^��M�Eؾ_�������t�Lª����TE*�k��sE��;�eG��b�
=B��1l�Q2�{x�1�BT���gHJ�Ks�u�i����.Jp=��	����f�I��3] ���8�x9�[G{n�W��K|�ylKZM���.u��Ħ��n����c'�٣'�wZ|���5t1j:�I���OU�H��*Hxbw���eF�mdR��y�-G�N�8 �v�]�ᴘ@vީ[�=��^�{�[$u~� <Р �ź�)V����^=�TnuT@]�/Jy}f/p=Rw�%9��S��m��}���6T�\!s�$Ѧ��WB�GޏZM�0�x5V������L/���*�\���sj���b��V�"FOc���-�;פ�]ҾUb*�r#�+l���G��_i�<����M��>0[#��Uv��zd�i4Q�U�ѨD����Y"�~��n��$Uė�-b�,��9'�&�-�'E�&bJ�2&͡��b��10�X�ƌ@�a8
�� �0](��Vk� B�y|N	�{�v�{�d�?C�v�}�)?�t���^��bG8��>�Mէ����?�r��W��H4?�њ�	H�=�
��K�IC����<��ɖ�Y�+<��B�q��D�o�����>��Aw�T��(4Ӄ7/wːw��x-䃑�]��K`O]ҁ�Ĩ���e��9XX�mգ^��pTَh��Co��n�=�uh�>�Qe�5���lz�R��tn߂3�V�#�8
�`
�I����z�{��c�t�8��� �S�6H���b�_��])�cjn���|�4���R�QWDft�R�9��m~�QA�~JQ�CN��8TݺZ犒,��k;�.�ZP��D|Y��@%]�:&����gL�D����,K�����#!F����h�m�c}�h�M�h���}��)�mtj�"6ø�;�h�0Yz���0��!ntbnszҫX���\��У1����G�ѩ?��ƞ��zt�LIt ��a���Q{^1\Ա�8����]ַtEu)ڜ?�䶒�zV�׬�1[�/`a�H�%���OXVJ�2iuJ�C�sw������5�m���I�Mka�X��,��m���h�U3t�����Ḩ��F ��Π�)8���)��8���*Ŧ�"��ϗ]Gg��e���8&�榆X��ER��w�nEC.�H��m�;9vػ��GoS���2(��)���
i��<���-�n*p�lE�A���n;�=��
t<�,�bw���j��k�X��I?��Ӕ����!A�%݅�63T2C���$��	�|tdrT̠�1;��`1�EsI�}�#�,�^E��Ls
e�����	��|��C4����ݰ6Z���VH_�g #�׻8����*|���������NN�^}��;Q$�C��X��"��7���kl&��c�ԷE���Ki��L�v���܄�(/��M�U������G_�����CM���j�%Xۘi5.��%���`P�O���:�^��,_~�2J�iPh���-�;��F9�)U\<6m#��m�ھw�{�ww�	�����Y��$vt|1q�]!��l�[^��n�׎����t���`�H�c�A�S��&���HT��n��`��-�x-N0t��\M��zq5 Don��5��+�I`���<Q_$)���Kl��3p� l{���1b]�{~�L)�ɵ�'x9�m��95`�S8�=v�%��>=>��z�^(f�:u�O�Y�~4�X����A���st�����iA|�<ݸ�+ \q�ϳ� t2#*&����z~��?�?!Z@z��U�A�q����ƶyQ�^�=ZX2��ޡ>����A�f,չX\��搠8��Sa����r��g�3�7X�����ɬ�P�D��Q8� ;�)����*ǲ�fS�C��Ov��K��U\m(�/���H�
G��$���4[iAE�dkx0Z�����J��w�2
�4M\�T� r��J2k�W���hZv+�qY�B�R�B�?���0A�U�ZYڇ�->���b]�7`���W��}�G�	ig����S
�l�?�����͠1^�'�F>1F���{q�%�g�#:�-��o�G{/W		؞��k_�߶Ɣ�L�hZ�CqE�~��-���(��թ�P��G0���F���)~��C�忭���3#��qP���Җ�a~>�ɡG�z�Aٌ�?�I��}�n����%��	�-`��#5�W �.M�喍���2��h��Yzu��/Mb���FC��;F�t����Y�ԥ�9�����&�\�n�M6���僶8W�;+"Q��jd��:�=7C�~��c�/��
�b�jN�z��c�g��c���5Yob�'�@hy"׊�[�Td8@?oh��(�U�o�x�0���a�n]Ԩ� oŵ�Ñ\���������O:ZҹS�&��"z���O�{�)�c���Z�T^3C
M�[�/"tZY���n�!Z�s���3�1"�zj�ڬ^9���0��nǙ<�QȜ��V�c���Z���,	�^u?�MU��,쯯w;�[�j�E1sg�B)���ё{�}GI�n��������9e�D��C��4��y�T��Z�H�[Ѷ��G`��u	��.��r-m��M�ʹ3�㿍�k3����f10Ʀs�a�u	q jZ�%���u���*� �\Ʒ{��I�@�.s�����Ҍ;�'�ǝ�,Zp��t���|���˙δ�f_Gv%�F���V��Ȕf�}�O6e���c��A$��¿��l�}O�sdF�ЅPJzԑ G�`���?;�2���{���"���-���'A�2:��^a��Q+����fT�M��oh���!�I���*Q0gOt1�Ln�ke'�w�=WAcv�nqz2)י���?��F[|�6���y(#� gꋴ�VƆ�V,�Cӛ�	I�c�g���� :C\���*� D��)�|�ɟ��2�t��ľ[�
�7M�~�u��[��//e��ì�k�Y�[���g��S�ֺGB\i%�'}ʙ@�0K��Nߺ�:dn��G�g��6Ըl2"뙗e�]_��{ؓ����b�}�����u��qc*46f�0��#&ZY��`
%kC�cjA_�ju:��zM���eK�urE�E�
8Y�#��U񒥥�
��W��u�/�r4���*�xr�oB@�(;d!7��1��r�u�F �P��X	�e��6G�M��Q����bofs~�a_V�w��-UR�u��~�z߰ǆ{�Ԛ�X8�����c����w�dᷲ�dً;�����^/G�a��D�}�KP��� r�Z�m�P��P�bqz�eb' z_�xC�y���7�}��кk�D��_0��'v|��6h�YK������.��Ex���A�=��{���!��dP����i�Nʃ�?neM�f��p�7&���B�8���8x�#3���/	4���<n�~���rs�����(���1,ng���''8,z��/� sRVo­��ca�@��p܏dǱ|�m,��&1Ԁwۿ�?��"��P�h��8�;"Z/�Ș��TM�������Y�2��ۘ\q�<�>E*g�싸O7���+���($d!6���eH;ݿȐg���R˥\\Dc�1�#�� �*����Έ(�4�X
g���^��v$XP;s�K�Aϛ�^��2�8�f��⊂��L�ij���P��5Lt��e*���:�<z�~t�����b5��ɾ�6�6�E�R�>�����	xu���9��_q&���I�D��`����r�pA3���K��-�]�=��+����0GY���uI:r��BQ�儖���=��A�hcD��u���Be�U�UXdjuhʲ�Y�Ӄ򈺉�a��_k	�,��t�1��c+{�>�����IZÞܷ)U������H�kSDBd�0{����^���S������n�xr�ﰛ^,��>ʅq%�]`jh����0��56�� ��Aooq����wMbd�lDa�%~r�$��'ƚ}�&�XMfQ-�7��i+���8�%��J˼$��y9?��1�+���B{��$_6}�g3�?"�>�;�X�5NGʃr���������!m[�e��zpC���n�m8X
��lH&�]�+���N�����Rw�ok��
?]4����1?��=xԮ:�t>P�/�EDfƍ�E%��@��u�]� �!�{��ߞ��H/��J���+�����m�#��ԡ*�З^K�E�!)w3�G���2�0��
4�3Wf?�`8�g��j�����D�6+lR7����+�*��X���s0unfF�:)D��w��A����i͠�Gy�S����h���Z�s@���\I�\ɒt�5u�(:�KYOl�lu����`���]�s��`q1~צ~���SDE�BI�1�n�ƐE<�L�m���>ym-���+���!������sԃ#�6Ʌ$�8<�_�A���m{T|Dɩ�9��T�v�K�o�W�L�_���Ũ�y�āya-	��<x���ofí&ԫjf�[{ l-cC3@b�591X�oa�Y�eY���Z���Y��DǊ�����	Y{���M�I�rWP<Gj��v�C;���Y�����IU�s�iWT�bbo)�-�мʖ�����-vQ,������J|�Z���@E,맢ŀa��\�ܷ�v�@P֥W+]=�u�ݑ�i��;x��r%�w�J����{N�OW8!5�ݓ�Yقd@)A��k��	�Xi����Ƞq�
�U'�^��9e�6��G��&mFT#���ނ>W)�	�e�5�W������o�W�FO����Q��n�I<)�~q-���H9e��|	���+(�.�$�ٴ�I[��Lm�J��.�Ĝ+��������,����c��?�<'���B�}ԭ�R������{�^��d��Ŕ���h�r�2T�H�����н	�^�bYlm�S#�	�G�Z�
��թ����h��k�|o+�}�Y���)�_I�o��Yv�Dhd���\B!��9��ټl�=p�;���9����Y�dT��p��G��x��{��ayM{�'I��o��gi���;9sP���j�k}�X����p8���}`K
ś~��Yқ�k�T��0�f��RS[����n������Z�Y�K����ԧT��^��s�K����ӯ�_�`(�ht���g��A�������k���LH��*�)��F/DrmN�����|���й��rz��c���W,oaZ�U�`��f�3��)8���R��~f���H|v�q�ŏ��P��,��p��H�e�B��?K�&���G�&�^V�pF�������;�/� �O��K��_��������n�ַ�t���M}�S+ P@�+�b����<*�]�}��_��v�
邏Pt,��v�g/�q� �`�6���ک4���t�|����$+	U8�$X�:�`T�v�+A:0B�d�XB��C���Z�i����Or��%�<9WU� "��Oϋ(�
�*4b��P^��Q#��yU�/��-(��wlS#d��Brۯ�n�j4>O���y��C��Ɖ�@6_���x���ԧ�zq,�i#�����,�K�.�g�P�7d(��N�#H<�dύ��-!�q;��6Q:�a9�ȩw	Fa/�����Awx�d+%ħrꖷŤ�vt���erYE��&A�9��R���
n��{��:����Z,���~�ڄޏZ�a6�������"���T�C�Op��S��X���gyD =^�7��3i���+�B���m�d�[u>�!�^#�����6E. i��C��m���U�Cb���o�fL%�D֗��~�lK<c7�ȭJٲ�,%�͝��F�3�#�n2�E�9����M��h���S�����\y�pA�H�o��b��|F�|.E��U�3�/��C�Tߔ�-B���to� ��c�{�nε���HfzO�(��E7����x���%̉  �ϷwN���v^^EhoRڣ��eP���ܘ-������T!�@�vǓ�Վ �W "'��
��S��e�'s
�K������Kn�L��>�z9�=f��TN�R���3�kp�f�>pB��C�$���t2F�#+������"�CKW���&p��	*�QF�w���*$$Ƕ��[SA����0���NsѸH%}�l}�����ˆ�a��O\�c�	�!�{u�n�$�Q��~%, 8��^x�w���(3�u�e��0'ѝ�R\
����
Ebd�����^CXí�S �=t9�{�@��%^�� ��x�B[1+�ٍ�[��sPYi.T��N������\��MJ@���Kz��/j�I,>�
e����EI6�mZi�0� �����rG��Z�7����Jc4/ �by����
�^:��;�J[��uc��W'c.��gN]ȭ5�����M辁j�rR��|T@R�&]���|J��/��7�/7<v��O\��8�G�6�%ͤ�~e�� a^�]�j۩Kc8���=����Z�P�U�Sz�&�%?v�t���y����Ӵ�)Hyt2j��i�3�;^�W���|F̕ѪN�H>��Ş�1'��� �(�ؼ0�f��P�-Q<���uoȂ� /��"J���  �m�g��or1�2x=tb�y��,���g�7�����|q�=ěb^�?�v86�I�60M���{��}�۔��ޝ�ž�����l�j�S�ݶ�,�K¨�d�O�a��E�趬ۯE��3�Mo��K���D��ߓ��-6g�7ѐ�dl�g�b�N��Q�H�9�����ѕ��hO�����'{�_˿I�zO>�1������_i��#X!���Kw�9�=�����]]O.P��]�col����z<�h��%Zvy�`�>A��8H��Z��ױx]��f��f0oCy��UsA������-��#��\�aq�#26��DB�)p3lDk����R��8ġϝuI�^o���ی#CIxeƾ�6�#��;�e���J�	;`I.���E�ȑ�D�z�$Ν��kX�
KW��K\^Ġ����g��i�[���#�x�vTvfJ�������G�4FT3s.����"u7���T�ǚzU�n8R�yX��2 QK>���u�9��zϸ"q~��e�\,lv͡\�l�\E`鼱��y-�v�{�w�!9ASv���P{ꍌJ��J�-�6Ba���=�h+T��͂U��_{��N'��.�n�/j���^Ax8K����y	�'�}�]�O�Ѷ1Өgv�021d�U�Q�Hk>#9�&!�ȗ���C�.�}�%1V�4l����TD/��{�b U]�C�ةT�h��j�oij�vL�����z���~K�s���Ě�$��.!#�r��zD�m`Ɓ��IT�a��|���Iݥ%f���;�m,H�6��NN���:��ȝb/,��ݔ�����>�i�~�T6<@�x����'CU���/}T����z$H��K�(xK����X���1c�������T�E�-Gg}B��(�"U��
Qi�Dp��z$ �y��rT%]m�l�7]���������6U���'��O�BC�����K����h��uuh/)��Y�67��Z������dX~�KGX��Ε��?Z -�H7^wńԷ�`�&��O��]�<�:%�XWm��Y�S�CtN�l>lym�a��g��,���H>}1/$�P~�E�BVy<���Āgk���STaS��T�3r���c�^���栣U�
Km��l4�RU{���gھ����v8 ���g�'L�]Y�m��\��̗8�}̘\2���k;�k?���#l�f���*Ҍ���(H4+��b���m��E��m>2a���<�z�#9������&ƿ�Bt�?����r�͋��9!$�@6m8��k�݃;3�5Ý��8���k�;�����,x�K'~`�@�qۺ�X; }��HV7��+�qt�:d�U	X �Ǉ��zK�:X�vN:4-�N��pSw�*����Qx�+�h"��`֭�ap����-O*S*Fe�D���@EY�
e�q�CT�'F�U-+\�C,���o�(O`F7�o��¬@��x�x���\�"���3|����31��
$�ހU쳙c���~�������X�;kH3j��h�:�K�01�ҍ*42f|͚]�C��ז4�r>2�B&�`���p{�z�,b��&�J�\r��\��Ǯ64jZ^d7y�9����iK�OE�ׅ����8��ͭv{�\5vҎ8�1����!Y`-�1�rr�+�� ��F�7��%(���׈���/�'�O���s�BC����oS�\�m�N�~;�&��jVg}c#��P�3��$�b���y�}���Aj�fa ��>������o�޺U����3�6p��r�;f���6�����uv��U����Ӂ�i�M'�C�f�ﶰv�J����ǹ`8*���Z�ٵ�R����e8N6��<֤�[�ǻ�{qk��,��re�H�F�/�^��'��R�N~74�x�$�E�+i]e�]�\���|�����)i`Uu���-Jt&P���~c���2�{ә������%�����&�ۧ�
P�;�����_�M(@D
Xj��=��][�������]�F=����M3�S�lۧ/�^�1YH�r����v�}6��7��E��@H����sb��6�Y��M�o�(hRvEۍI2�<O|�5Z��J���ɰo,Y3̪��Gu`?��])�:�z�Ur�{K]�u�#lМ�>ʹ�#��=
�ۃdʪ�9*;L�o���������J;�=!l(�)-�(��\��^k��`il�DJ�w�"���<PҶ�	$/B'�<Z��֮�a�]���Ͻl��lS�LaGE{@V��^�F��(�Y͐�����K�ܵ��ҫ��4'�D�L�f�uw�E�rA���: cM�\`��2�#p� h�Jlx�\�'��fg;H�4�r+7~�J��\��*��.��*c\%˒cLx9M��
#� o|���`����$�=����-�y]ȯ�=��W,��H����T����&\ a�Է�x7D��D'9��Rtȵd ������&�Ⱥ�|xm�E��?��W�W��u*��ý��^P�:�H�{�c4 �^��}q	O]���䙼X_O�5>[��DI\�3��S��g�`����-�Z��� ����9��o&�k9/[��\8�L<��M�]x�%g��oAyROurg�O�i�J�ݑ���.& �
nI��9��$I1|�#�X�E޺��sk*�{���2��$3F���	(Zd�dVJ-?�io>3�mЈ���z�q��H�nM�u���O�!)0�=��A�����4*�۶,FT�|��Y�����P��O�d�Ϥ��f����3�<�������{������w����+V�"�e?��C2�zq�_����[R� B&�Q�S�
	�(�ЗK�~�w6���$��|�2C��@$_�7�IO�ʓ;�p���6�~w�k����:����7��F�Q���W�A����F�8��.4��܋X+Ҳ�
�	��=}����	0	���%��[<�7��k!�M8�L�~S__�(x�z9����~��n�dl_
i(v�NˡY�a8��!RCf�'6͗�ʜp���O��t"�e<�5��ِ�%�6��P��;l�J�f��BE�3S�(�Dm=���o��W^���sg��$N��=�a,U�kdt�ȥ��J>p�&��Ji�Y����C���X�G#�./����	Q��'����r���,�5�g�����뎜$�sO^K�@��Q������	��*I���|��9��uj��{����F�Vρu$�@k�`�Zy�K�α��	:�h�я:��dϣ�$5��9c�m��A9Guʿ��h¶l	��n�,�J�3����P����4�=���K�q�ĄS}�H`�y;���<|��~,��j�y��zZ3}��c�w�$����zF�ӧ�Ho{hoԡB1��Qp���c��4�!���iK��� �Χ=_̊�s�f���:��|��킺�AI�b�^���Vlv6�Q�Ml+w��Q=��۲���u��e!��E!_#�O��V�U\������t[�[�L(M�ϫ��/F���&����e���7F���`�i+Y������U_)��f�%�G;P#ԕ���Ō̖f�L�_�p�iic*o���?b�$F�� �h
���8�k��r8�{�:��RD�P�����L���Y��a�~�}����Z��@tז�R&v��Z��Q���g����(�Mk���_���~DD<�����.�y�|kw�!Ey�U�0�ɾ�?{Ğ��D�-�a���M���^��aI=~\��c?�%�:w�-����ӏr��M�-Z��+c��t8��
o��-�,�����+t��֖�Ά ��f�3H�����*6VT���PՓk�Yru�����S�Ý�����A��G���M	k�b��RLL�=�JF����Tg����[]s��:���� �|i�N��6��P�W�q��2�6�HrOHb��c����~��5(�߼2�^�K��	�@Q�()Ɔ8~�%W�.�*�P�;�|�����4(�n��46�C���3�x�,+�D�~�$��O�[Q2���L�i�tڑ&Ճ꧃�i"�\6�M�<�~mH�W���V�U׀.K*�c0[�D��(鍓��Cn����H�ų>�ƺ%a�N�9x��A��8ށ��fާ��](�8��6��QZs�ys�zw�}"�����Qo@U��{��w�P}IkW��2��\��ʏ'� uݹ�~�E�۷����YAW�c� ,��$+u���ȃ�����ƒ7 �׌��e�c�����j��A.�Ɣ��0"��S��g�,�X�$�b�=�S��/Y"�L(��Ѱ6��E/)4!#tg�.���r�9��h��Һ�~,'I;�cp>��Uw|^�V�e�7뚥-��@�h�����T�H�ŷM�nBd����Ֆ)˜��+lf���I�m�L/�=��BNϦ�-�{�*1�R��؁Fd�8ml<d�[ː�o��zj�_<��¦#�Q9���?��F�kŬ�f;ؠ!| ��> �x�p��m�+��v�0�!�䠬�r��͓�^��| �s�&2Nӊ�h��!�{��l�'ߥ�7�5[�zy$E�������������-^Ȋ����[ M
�9 Tj'�Yl�b_�6ΉT�o8lj�W�6�a.i5����w�3���܄��̃Z��:ec91> b���m���L����"9�XX`~��)#V�?!]��O�|���KqSzK�u3h HI&���e�>�	#�.���XЀ��;��[G�F�P$�����+MM��A�A��GS+�R�g��+ꦂ��M.S���p
v̅�m�8\�B�!3��`�P����#��L��=��&��� ��	���B����׌r�E����R���Q�l�񫊴�_C��.'#��$�����@ߎJ�0)ɺ>�l�u����lir^�T.��J�P�2�r����d��&�TL�ow�\�A�զ8�f٥y=%����%��۾b�V�(�3�ތ�� ����oL2���P��Nf*4+��u�{ɕ����DA��d`LY�>��,��Q�b<sчz�B޹��i�<0�� �Ή5��M��(�c!�Ji��ct��{6� h"�'0ǣ�,F55���`�j�4�ӉJ�j��߼{S�\��I����e����R4+�Ѓ����إ�,�}��n�X.����#n����p��v�]r��3�3ߛ��Ȥ1�6��h�5��V���&E�_�ބ��Ў��&Jܥ܄�����(X���2,���X�r�'[|�-���*+H�j$x�� �����2�[8ؒ���@�$";��Ӫ����S/G:1�E�&&a:���� j�d��o��	�`�u͈k�\�j�uW�Ƕ��IE����V9w_,�#G|ulK@8����m���Y[�	��\�#������>��Mvգ��&�h�#�yn4
��2}\#����<t�����Rw���j�Zr� �rN����
�ROTC��Ø{6���`k~E��%5�L���HNxd�b�1طy[t�ES}թ�U0(��#h�W8���M��b�?X�s�pj����T�O5 NH'�v��u�kBq����Pj,�9��w�3������3y~Ǿ��N)p�c%WE�+"Li�p5/m�3	6�W_����>�E�0�V���z]�͐������ �\�C�@�h\&
�N��9&d�}<�wUr\��7�J����[��2������h�����j��	!޳��::��@�R.� ֈ��>9�@%��}���%�W(���"�)�55��V	�E��IK���^�ۤ��:D<B*3�ޥFv��Y�xp�#�v��wXBC��G��0�y�M�iO�6P|��K�3άX�#V׎ԕ3n!-t�����JD���|��A��i?��c�+w���ж�e{Eecz?A�4��Z)T��{S����T<��,v���D�Ǎ�R�{Hzr�&��/��N�\S�bp��, ���2p������^��t�C[E/��B$��\;��C�Us��{z��g�Zr�����Wz�L�f�e���]�`�T�n�G�x�q���P=, C6̹$���,��v�g��_��Z�|���@d����C%��o�0�g��{J�;�mZ��-�kG2ցՃ��5G�J- �<���� []�!�Fb_r(��fZ���>�{m%���m��g�ʉ�b��Ŏ�p�n]�6ՊP'	�a3�eE�n�%j�6 y�����ًL���Dz�D��A�+��k�k��c␃�-`u��CKv��m�����7#u�H�A�������|�+�a?�v߫���&��5XV��`������N.��*�������]�e��H��Ժ��Fa�3̼c�p��,�T�0����@�����2������2�/���c�*c�X��(�����[x�҈/��{�k�2w
�q!��Ab�m�֓'���ԂyD_������<w�����r'Ug���˱�3ܧA��D<B�b��8.%ySS�36	�ͺ㍀�l�m��}�Q�$j��p��M�ȝ�$���h��6���WT]���^�ƌ����G��4Y�>2��}�fDV��7ie+�0�5����Z�<)�%��50���0/��,+��*���&�T�d5�����5�����:wI�����m=ߩ�9�vfފ��d��$e^��'�@����$�)E��_R���ء}�]�����ڡΎ $7C�hS<����7�P�%�	��qQ��:�&���gf_��|�b6浸�`%��ߢ�%6��s�=	�G��loP�Y΍��3�n���"�^?���.:��2��:icfh\B�c��ΜU���� �Le)��T�`��:	���W�� d�q�W&9��������>��3�/�/�Bՠ��ӣ}j�M����"�)����.�-}��/�~G�"�2��/%b&���(�$�Q~r|���rX
շ�%�z����.Q��/n�Fs&�+�i��6��9���06����mS���Jh����S���P� 9��0N}7m����N�u}�@�?����W/���0}��ŶU��n֡bV��O@��by���W�,/-����q�TtѰ��ۡ�3]���YaMH
	�T~� ��K�.��tE�k(y�C��>�4��]6&��tEb���7��nѓ��b����vn���Q(X����ۇpE��9GL�l���z#���bp*Ɉ<�z��[�@O��<^߷ί�.�5"I��q�_;�W3�[��9�����KIHs7C��%�]�P�R����v�y�����^t�cw�OJ*˿��uom�� gƆu[Y3+Ffd����N�_��hO
3g���#��8A���~�Nt�r�6����r'��u D>��Gc1�S�O���{"��3�I��0��Fe��:{Z��[��caþ��UB���+9�^��}��eM�$��1��ީė�ѳ�.�2|�ݖ����kg�Ʀ	�zy��~Z̼���w���C^�
��<�5�K.����ϵ�����i�>�Y�YD6X�v<r8�=A)'<��8�1��o�ñ;�����vN��_ PLE�����Hq������b_i�����2���>iDAn\!L<�=�������V��w�c�@)7�	z$�6��\-	g-\��]_
3���'v����`~��k�k����(�����o}ޝ=À#��X_p�Q\?H=����ݚ��C����4�)~e�=eFE�퍯�_�@�2�e�X��r�J�T]崾	��Y����e��q1)p�C���>�f��Gr1�k���
�#t�'{[��I�N,M!p��$8DG��Oz3����d#�԰Ml�{��;�g��諩�5�7���r�F3���E��}���m�-HYJ�lO\jBQP�¿�����L|q�����PX�HG����^$1Q��5�ͥ'��\�E�߹�b��*��t�������^�TD"f'[]v.���ė�^����z���ւ9���9��ᖲk��aCD,%Z�wOW�:~b�Qi��P����V��m�k!�uQ|h��mOqNF� ��w��~�3���f4���{�@H K՗I�=&�c�_�It��՞I��A�Z��8�A��*��[�i�}>3�6,��ȿ�ד�jb�j킌4}D�Ě�ii$؝������v�]ڴ=6|[��r�ڥ.$b�T��ș`m�^�����G��nQ��W�}�g��T �p����g�`3m&��k��y�_�̩U����[k^^����A�v�F8��H�V^�u',�[^��m�lN���4�,�/�\2�l4>'ϛe`��̕>�L�9�a�*q�|�X�R�O�
ZY?�|����Y�Ns�{��;BB��
�>���R1�J���i'f�0�b�!�뷢������g��u�dدXv>���p���UR�L�^s=�H8F7���D�v`�
3<@q��?�O hN�6�f�����	��І��5b\h92tכԹ��1NSWM�� �)w���ܫ"d��V��n{D���7�L�δ�=���\��t!w)�64�t�tG�?n���M4p=�wc�w=�'���⦸�Q�si����t-��c�v|Ӄ�/3�	;��3=r���v<7�9WI?�6��x}>+Z��y���։s��m)�<����>�ŷ��\�.�bAwJ`����0m��,�m�h�W*��p�Ý��|m�|F�AY�ޱ�㷭(ߦ郩=����+�b&�k+������~�A��no�`�[վ]W#�����bP���|��$55���R�U/��:�ĞS]�pU��޴3�iеϭQq �ILK�)�c������D��� �O�:'��鐛*~���ųRi�Aj�y�Hg���#�Q%�v�x4ɢ~��smm~n�����%�� a�1�	��q����M	lE��W{��:����b�ʌ!�.E"h��d��@*�K�9�\�y&7^�r��]�ql�:�~@�*��M�с8ގ��Ze5t;I�ϒ&��ǜj}�->�siU`���Aܺ`�|,vF�Ne�6��r%1Y̡��ҫ]^j��%�^�e��`������R�zǭ�r:��6v_V�P/AZX %}>}��4��«�CY�𩣣gcb����=��U��{�q|��|��PkMcr��k6Ӂ��x�h�v��S���c0�;�c���u+����II܀
aV��Ձ�)h��s;_���cUq���˺sS-�k�h�"�vv��U7�R��BG�jwq[x~������8���Zܨ&`p���%�[�`�#V^fy�G�6�)��Av�y�s(}>��_�P,�#懭����>2Mya�Bu/��.X?��ZUW2HÂ�{��1���R��@���z5X�O9+� &>@��^��Hc�_J�0�,�� ��Pm�*��N�Ze�dp����5�[�ӣc�}͸�����QNЊ� I�S��quڦ��AOl1�iܸ ����B�G!f��Z�k�L3�>T��fvR��溘\N�F���}2��ׂ*�D�J��ƚr�EЊQG+�5"8���͊�0j��=����BC�p�\��0��XCpv�'d�{F�������,	�w��i4e���8P�����𾺝m�p̓�o�fL�FN<l��F=�B��j��{{��k'����|+�_U� |B�^�E3������,W�3AZ���i��*���0��5ri�x�On���.��2��pE���a�LC|%���b�GK�X��7Y��&��j�U.^:h� [m��4p�'���SW�6�oK�T�_��(5D%��^��O�;�p�e����2�R�<D��q$� ����LīB�"zO���B��"A$�;�*5���̸KK�S��I��?ꕙ!��	�?�9�{���2��V�(��i�Ƌ)ȥ[*x���.��b��@qS��z�\��J;B?W�#
����\�Nܮ\�u�5�N�Y�,�v�T����I���n�4,y�((z�L��?өZ�,�*�]�˄���V@�nW� �����|�����P�\�1��
���.B�۫��٠��%̇Ϸ�2xEJ����`_��߃Y������f"_+���JT�B���?�u��ve@����Xk���f~qi�I�w���R�)��s6��?Q$j����Iu�?S�G�aP"=_����wpi��0��ʒ��?GoW�Gyg���Lf}�0�6>f�&K�{ �=Q|F��kk�~���!ݖ��c���;�#���Zd�0�@��.��cmo�x�6%c�$"e:���=5��?�|��\�E����ɯ���{��)ٴ�2x#)�)��� sf��;}_>�H�.� "�&-#ɒ-Vu�����e�ʣ��e8�tP=��W��'��m����O6��K��^{B�g�{�{fҤ ���|���T,j)���)��x*��C�)�� B���9��;���|C�,���
�(.�Lscs�?�4���Z;R���iv�ѵXĦ1�4��e���t�b9Tf����p��Q����D�6f��!�
��T(���n�,�Do�I�}����D)Go��C��n ��.6�����i;�������g�5���K�͂i����ZԒ`��;���
�ܗ-��C�lgvm�h@t��qD��nl���+^@k϶��6
&�H[��ӑb�r.�mʋ]���܃�?L�N�z�m�}I{[D7��>5��e`�Q?L�d��7V��j��^��mK�%�l��q��~�$E��d�����ro  HU�����Dh80��� w�dE-\�.��u`Ad�?����R������~ǉ4,ծi��HJ�=5�i�Q��?��ܙT���P{rd|\4|�A�`Y��p�`��|\5w���o��~v�s�.�u�$L���s����-v�����q�\!k˓!=Y���ҝ�Bq �C��fMZ��:�w��l\~<Amtc�ٝ�@5A�;?�6���_z���?�����Ou�����E��攰������?r��17c�Q�d>_^?��=5�����m�ʋ�m�U����6z��j�gm�t��X��̈���hv\g��ċj�-���!����Hcnn�O)��y�o&╰[��lrЬk6R1����9��h�(Nũ��˟a@�RSMj ���K�v0N������������XX�'Δ���Q�\�!/2\U�Q��Xm,Y3���gm$��1z ��ye�m������C�G����h�1�0w��y��Նc�u�s�j�;O�!ɲ)��Ă�\�AC��/�aG=NFnP<:=��p��3XK �=!S��#;�j�������z̍�؋�΀�(4�&O�����U�F����ވ�����E0� ]kN�x
�]`먬u�k�)�La�m�2հ{Fw�/�U�U¿m���X�V%M'���G���J�82��D<ۻ�('Л�����S���4*;>�J=J�r��^�����i���)D�wy�#i�+'J]I��f�0� ����:/�t���n��q�7񫚅�<y�YܹM���n}j����kPވ���n�U��{dC
E��\�/��ae�3�d�랑��q�С�ꀄ�T�Ɔ��#�{����d��zQ��	�SؓrO��!��eEH�W�R�(�H�k�u�ɓ�[�ni���Vu���1k�z��Z�XSav#3E��<�#O��^��Nf��*�`\��~�vw������\qd��E�,����Ađ�����-�Tt4�8R����׸a�_o6"��qdu�9�xT(+�ˀ0Y$徤�)�� o\�{��?�	}:nA�L 1�g��y��_�#/�������L�̒�Y���;a(G�������UVM6,�?����z�G��+0��'Ep��	�b���G�I���V[&lY�˽��xM�#�\���R�ጤ�'���!P�<��>����@S�g}���\g#�?xI��N���(omp��]V�z��|84�`<I	�t�cp�ZH�Ҟ9hi�3!�R]u�[�r�+Q��t뭫����L���ח����$*.$���z����Ù�U!�{�].�|s����3h�"EžJ��UR�[�����5x��Bf7J����2F� �}���{����~C�)�D��B�#^�
g'�Un�8I`��] $�_^V���#_ F/*@X�]�mB"��+�����-JQ��?��۸�н�����ئh:��%LTe�����4+��39��ܴfQ![-r��=��"7)�K��8@}M˽���>�*�����ڼ��=��.f-`.���uFԧ�j��H��)R(���:���5#k�
�
��\m�)(V��/ͥ����!S��V[{\|���ɇ�U�F�q�g?}>0�5L�,�Aҫ�MPM1����Ŋ��Ń�Z$Z�����'�_1�M���?��A/����K]�����D�$�3`�_��_�H2�c�c���GN!��3���i7؏���4k���Mڔ�p�v��N^��'���6���Ŧ����}��O�� w掏��P����N��0M�x���Ǉ؃��(b�s�Iʚّ�r���oZj��	}��A�%���5�+�ߟ#l{��k`!Ա�%�"V{�t�Q�>c�X�4�#hN�L�
���pǳ�q��ۋ����Pr0p�`�Di�k~Ȇ++�R8��0���ܠ���M���2��d�u�Ɠ�k�8��G,����h��^�1��r�76Eu%r1A�h�����O~k�e*��}���ET-�Q��t�2�AZ�������ޟ�]�4D�]V��6d�h_����˗�����`�8�eK�A[�=vG�̶[Њc���˄н.���v���:M�cG�	�X��y���%￢6�-�s������=����տ���߽�9�'�g'�:�Ni��X�`!�@SΒ�9��K�(���@��@kߧD"R�.ui����O�C����5V����9�d������
�����H"P�4��	[S�U����đw���B�/xm�0zg�0���a�a�+��U8��Y�
�d�ޭ;�+[YB��?��U�ՄA@R}M�}����j��1M$􊓐 ���X��t���u������˔���
\��������
J���%֧x+����,0�Ʋ3�Żz��6�h��y1��7@�Q�a���m,u���!�� �h0t�`������#��g�zgfV;��=�KѨY4b�V�F0�k�8��hB'��ޤ�c�ZS�W�i"Q���� ����Y�VH	y���O�@��|�1��O��� �:&n>�����1 ]�(?�=򶐯Ny���+�P'�f��e�@KRq�]���&�<���Δ���=Oi�	4�?!p�ט�[�HJ��z�n�@x`�WJ���0v��8i�9���( `�Rk�vqޚ��>P�{)�����ՔRw��H�^�_��={9����Y���#��J<@#;$Y�8���B�q ��ddf�?p����\8�
Khx���F��?ݞ�_i�Wuc��O�ݴ.'G��Iƣr�2�>.�i}��x�vi�B�Ē�\h@����
�j�|���y��B��b��1�+eę�{�	�ݱ����L�PG]O\�@g���D�{X����m/I�Qr�sA��_��Q%��w~�v��g��Ѵ�.�!��\4�1����6�}�;�(F!v�u[��ņXNR��!�w�rf����d�^l�ݡ��1E[��w|7P��N��]�˧�+��ۤ7sMS�R���W���"�ѻ��<�'(6B'<�A�YaH�I_�g��Ɏ��P�[UaR��l�D�#�Ґ�2k�ZW�͉����.C��`���M�uR��Z���bЀ]��~�9;f���Q��pe���#��W�����߁I�)?�>�	!�_��F��@�S�C�'�Lc�h�	1&w��
�Prv5��C�׷�>�B�V�}�����p��uT>��0�8��/��{O�d#�!
��9l��9��G
�� �x�;�Z�i:a3MuX}k#��J� ΐ+ˎ;'�IX�S��H��I'm�;0��l,V��q[�!o����,0����@8NWb$�X`�h  �E��ߣ���
j�Ms-k��7���w�2RՉ��I�Z|���y�(���W^����v��	s�"����!��ȶ�(+����x���8[�a�U�{ҙf����jߜ�&�zy���C�d[��눽�����r�Ne�sɄ��4��dor�h/�N��Dbs�&^��je�̥-�}$��~ƽ�~m�����)�[�Md��t���1���.c�[/�ybIċzV��5�s�,�����d����sqRe�kr@i�G���*�qx hј -H�� ʈ�j��̔��Ҽp�9B��*Σ"+W,�D�� �q]�����ʹ%��G�s5,��$�9U����D�ٮ�y+ri�?jv����9"O}�.ddb-�>E%����a5�:��T�y*�4l��M�)j>���xJ����l��i�|Rln_�6Y51.�[v����#��>S���GGW�pū���-Ơ9Ƽ�c��,�����R�mG��Y3$���u��d�I\��3�'��,6a(�7/HP��F� h�R����u9��i�[�J�Lq'��06��8���V�`	�o�8�}M8zR�#y���i
��3h�=l7a�o�j�T�u�@M�Ōc���#Z�t�2�2j-��Z�X�l�_Cjb��G7П17^�&�rIXY�1*�����Ã���r\�.��]5�_�Qg�	].�#wpV��OmV��o3i1B�{���S�I갂�C4#�a��,S*Ȼ�wJ*��nj���'���*�Ts�*��U���1�y����!欼fT{�
c��% �ؼK�7̛\d?l��%��ْ])����y"��'�J;#>���C��o����Ts$o.!�Z�8tn�wB��U��;	������1�Q"��2Ĥ����p�!�����E��YE�CRBvn��ٗ)1U�)�ISQ�U�i�@��sK�����5���T�.LJdzMV#YX�?1�^}Ƽ�r��/x�F�1�L��P�HO��7p(�2����A�J��D<�&�l�Y�2J�Pb�Wc�=�8_VZ]�1����_`���E`:(`qt��v	�ln���O;��v��E��A�7�U�1		�M)Q�1�R�'n�d���߻A��U����q��2�֣�E/yYa�����瓊v�SB~�ǝ^NG����_�f)k�AG_ˉ��ǉ��ն��4O�.���~�j:������4�M&�����Oj���Z������7<�h3� c]���ݼpɑ�Y4+��@��4ɬ�3Z���dj�z³�2���!�1%`���e�_��]J�r��PR|���H"E���	�@8�Lsm�+�k�{eX�G1�����i�VQr�]5q#��@�@T���[�Q��)���$���s�+���O�A��@ר2�3��
]�.H�6�eDڗ%6[�wq�&*�]v��������� �.V��	!\��x`|l�Q�$��b�Qf��ۍ>0���6��D��w*FB�I�x�.?�V���X���	6�����F�Ϛ`�1O�=���G��%��E�q��|2��Sĥ��{�
�������&��N�(����Ň =�Q�K���{z	��GJ8p�@�������swA��5����Ɔ�� BVD�`26�RǪ��h�����6�]����/m�i϶�a7%^	��,�À
��Q��KYT�9W��4��u-B2����1�I�:�y��ф�����SiKXnw�`Z>��f�{��#��ӕ��Qh\.�=��./^J���^���Ӡ0Q�����>��.�Z��$';(���0:8J�Uk����`G��z���;M�q��=%ҙ[�#�a?��#���h�b_�:�e��1g�Wt�J�"�ȇJ2�	T�z>� � 3T�<Y�B�ʸ���̮E�\����ʞ�OF~��Z�q�I,-2�%��d����$�v�V�7.`�R���Z{H>ȁ�W7��<zoO�����f&7�w�[�Uh�#Y���Oo��3�F+z�p>�B���Y��[��A��N�}�l4���)]zӱ�Ǵp7��]�fY#8p�&� u�j�ADTAO��#r�����TE%���Y�㷼����Y8!�}�X��wN^��a��ݘ��zr�;�c���<1-	7;^,"���I��G�<T�C�iQ�	x{a��/q��,�����d2����`��.�o�p&C�$}|ҕ@��I���@Xb���hZק(MFURh�f%��\���׵W�����H�m@:��(�
MϕxX�teucШe|e�X��:��Z��� �Y�֚;�U��Z��;c�^ �8�ꁲ���74��O·��j�λ��A���Bw��������4�VPB��j���㓑P�ȫ(R��;,{.�LY�+�$t��U�"���߉%I��>�4k��.�����x�E���ܰwo���pn�_h����
C��̶U9�)+eT_OKJ���2{䡽YL�����I/�g�?%�kE,q�YB@°L����?.�����B۝��Qv1�_��Lj͉T/iS��_O����I��A�7�
�ŷ�Ȗ&�����7��?�ZP�Q�Eõ:R��Ռ��x�|�����G|uJ;��d�EJ=��1g�&ӹ��c
�qn����/�z�.����=���bԭP��e�M9/c+R�q�!�U]��к����v��Gw�W�$�A����|��$d�=2�H˔p�j��O!�����>	���*S�=z��N��/���iT�E�
-%�v ���@��+;;)��Nۀ:�_TJ�{�	�	��9Sl�,�ũk24t�3��h��5g!��Zc-��5�xѽ��8K�I:t��|R�e6lio�P]��&p�u�w�D9��&i������1Tg���n_Y!t�Cbi�do���¢��9k4l�f�:X�ed���'�y��{���P܏$�^�O�G߈�m�v�{@܅���.S!7l�X�-.�Յ�
�X��vܷs�O%�~������������*����S� ;/�z=-Ct�L3�����>�<? 19Xd9���a����E��[�dR�b��=P�=����Q���5|iWY�Z�GࣈGX�R̷�T�%��FB���R�EF��ĪE���k�g�k����� ��d�_�9�$�s��� �h}�i���p�I.���y%�W�9ij�I���=�j�������Y~�]��y�d�R����٫��v�����B�55H�>U��Ak��%"��罠i�U����19?Dy�"~+��
���7���($d��/@����4 �|r(wY�f��1Eo���>,A\E�*�tՏ�t�J��=�����&1Y�G��A���L5Dme�:P.�F]�����Ol�!+@� �0���t�B?��3+��?#*T�F�6B��ǟ2c�������b�#R���a�ހ�;�$����/�ؽz�'o<a^~��?�q��Q�B���$�� A�ډ�^��R9Bo~�HW&�Ѱ}�~��er���@�Z=��K:�� `�ۙ*��d��S�r�͂�&t�]^�,���ނ�XDeɲ�W�;#���1c7�����M�~P��|sF��|UP�>gU&^�'���_�;������1���th�.	HO�E�	ړ��TA���PL24Tfn�.F��*ٲc@2�%�)�NrR�r�}�����<&if)p,�]!��Y�u��%vR-S
�
&��*��6a'�����gm#���&*�n�h�Og]������;9�1���m��uf�f��M=N��?�Z�-���0�s�I�#�~_��΢Ve������܊쌛�[_$&�o�$�c���V��gn��%�O�����Q~����y�s��1�x����'I�=GC��%5p@^ N��ͷt�o�^I&`�q�i0Rmt_8�(��A�����΋�;������ȚS�dә]Ow&.�-t�r!>b��+��Nh��G��R��]"��ű	0�����%��© u�J��,��f�8��W��"�4��z��3�ǜ�%,���롨s��*�6�^�b��s�E����}JN3ȧ������pe# v���k�%	�R����f��A¥Rx.���/1�t���N�ִw0��f�O_f�Ҥ�5%���r痫O�º���*KJ��p��.�V]���e����?��/�RT��܈EbCs�b�S;�9,� �d��>�����:��s�Y|-7�X�ڽP.T_4cԺ`�����([�a�>P��p-�A*.i���@�
��*�
�>p+�=�_��N2Û`��?cY��Ƶ'dC�[2������0���#/Oз�t���#�?�l���=}�`���[�^���p*O�������'UV���Vq�';���U�]W��7�� �QϘcj���ܐsp_��Ů�el=n_4�bT�0�u��̼���PЮ~�V�sq� &����@�$�i�s�dlTW����3/�w3M��Y�`�jI����W���6$T�IU�֗�х]�e��&b�z��-��h���gkE���MB��P\~]K� �ݐ3y�������f���p�\�,޵�V��5��Y 0�8�ɻ�E�f��f�I˅�K��z�V}�2��?/Þ��:"�A�B��l�-������P�v��#��Ȗ��ˠCO>��'�?�|�fF�L��������{B��&�+8Q%�(������K��b��T�}�>�E1G���qy�<�����Ki�ؑ�.h
���r��/�k�:�����Ͻ��� �D�N2�@��!]aj��g���U����l.b��������P��.�UĶ AS�����hE܊}Dbx�����ީ?���f6�$7�Np�Oؑ���>F�_:r@�ʼ����ޢJ�]�����5�x\-�B�FR��iU�D��������*;U6���0W�� ����\Fh�Q[�V�ɛ�(P�D�@M&�p*�(h9]"*�<Q���0)E`�&~9�%�ǝX./�2m������6��SY��G�T�G穑	XX��jݪ��K�T�Sj�#;-$X�6�����)8�eC�5������̨4\���k��ݕ'��D1ņ3r&��ۈ�>`��I��|tțC���-,v9�q��[[���R�3@�����c��*!���"��T��po��l�o'[aD�4��>0,��]
�oI��9�vtzt�*'j����]P���Ĵ���N���!�x�Z2�1�Vף��}W;b0�y1�	P��e&��}w&#K�HR2y��gKO7P�.CW&Wdab��F�70��ȱ�B��`(�;�8/
!�:�)�4I\7ʅ�Nh� �~E��N\�p�M�cR�{%*nt����k/c%7��Фu��:����,��;���Y��n"-mCPr{�<x�"��{|�q�0�NQ�	��Q�D6Ʋ�w�=��8O��4b}e�N�|���W.��k�`Z�]b3Q<���$L�>]�a�-וF�����!�jo�}�F���h�$��D�����I��l��,�Y��I0B��L��@�������D82��׵s���p����p[%�����	6g�i�n�Ƴ嘢o�Ãs�@"�J�+�*��OS��6��L�-9�mh5
�'@��5aY�^a�������פ+��/ˎ5�d5�1�R��t�
q�<hp�����AN�@4H=A���k9��FD�Q�`�5�1`deM���vrI�S�r�����,
T�ܳ�A���TΉ�-���߃��uw�� :��fG���%2���N�D�X�������o��,�7XFm��hJA!������h[��=�_a~��"X���NP����	�+���VZx6�3@���q�p uݶ���cS-D�Wq����� �`伶PLO�])�/�?:��3��X���;��l:q�[F̗��b��?��Nћ�P�&������%�	c	!'�6YU�k��b�����3�|[&=��^5o��`�R�f��I����ɨ��b�RpNO���z�F5��5o����p6�QSՀ���7��<ʹ�1�t���T�ZX��!�����KPov]y�J��t���8;oB7���I�u�G_K�u,l�,a���%{�����H�qq:������y`z�y�#�;�c��a
��^��Ӭ-=j�s�й�Z���M�R?��ل�Ba>kqƨ&:����[�l2��!Cӧ��� ��0*�S�<. @��8N3�2^ع�曆��u䵢�a(�&\!"Ko�Qw>��_�z>sي��m�_��-ޫ

��r�����Kil �`���^XW#��- ��$ޭ�3� dm�%�ެW9E.�ύLR@�3�X�����^@W	�ӑ !i'GO���Mܝ�$S�S� 5������Э9����Nlr����>��c��]�>:8d�IJ��z(=�t��i,���տ�� �=����؞5�|=�Y|s*V2C��f���=,:zϠ��'�0E|1��L��kom�0�S���f�#e��k�y;��ƫ�v�m�d+�a�|���7�bd`k���"�u�W��kv{��f�W���Y\�����'f$Pm�����X�9���o��jʝ�ݜ/6��ۣ$٘_&���B�n��G��F��!�5)�5��Q<_�١������C��v\`�ٙ:u�M�\�w�q\3~�G£��\�e������F�[���g�/��q~W�C�HV,�Y��"�cC�U�-�w(��~s)u�I�U,�e�^���]b>Ԩ��c7��.��%��*�P�Q'H':Wh��^�(�~E��O�D�hR��-)*`�gT�J�c���Q��T�u�� d �.A��n��K��A@��$J;U��\w��w$��"�I^�3��@��A0ݍ��T��9�5��ީ�-��%Yy�� m3�+ꑛ����.�2�ϩ�D$|���NM�w�h�o�����W,ܣ0H|&�5O�ޙU&�{�Ƌ�@
q��l��~����__��[�c0�s��]�����9�T{�Zݲ����_���j�BX�=t�l���D�wz�ԍ�:o?3�w�믠l�q��4�.D��'dA��ׯ���"̚yĶ���O�}Mi�TW�F�Py�|��������L)sB�b�X��ڇ�%Ӭ��U)$�=���O�4C��惔s�����('m+�p#6b��)A����>i���ːI��Iެ��R%��Ʃ��U�;]礙ދ�'�L�"�]:�R#ݸ)t3C$����͗gn�]�r��p̀�q�Dm��e�Zy��RFݰŻ/C,s�[�����OW��?�?��m��ZҒA�ڬ����N���w4J� |�e����=���Z�S��2���pΚ�:��;�A���%�eh�@j��tmNu��O����Y�6.5�j���e�7�@lZQs�uo�������u��$�`x>J%-D�؟����Ƃ��'�a�'�	-��aW[�B_G��-`�b�� v�1��������l��J�ϙ.x֤�
5?��ǀ#aT/-v��\����:��~%�(
��$�;�6L�XD��a��u(��8�,mS�ӈ\kOa<���W���]�󯌞ì�b��u�_?)��oK��cdP���voVV�1�_�޼A��;��������w5��P�Id8Q$�T��I0�2+�M9��Z�����rV�"8K��y��_]o�d��"�8��{|�X ����l ��.��6� ��򉌸J����텻�5nI!(�+�ER����M��jdE�fR�N����5�+a�^CZ=5#z�v=�@�6�vNp�P,j�XR���,{4�Z�AѕX4��~���8�w�8�9��R`F�ͭ����04�"i��V�K��1��ɪ��E�	�s���c갩����zH<2~-�����U和�s8N#X�bK%t����
��������0Ly�`�[sTG�2c*b�o���w��Y�U��<@R�a6�m���+��2�(����&k��F��t_�2_��`{J�=Xa�>D��;��-�QFv+��U�8i R�l�>l�S�2(����y\�OP�Ӌ��j�]w��7�H@d��e}2)�$��P���'Z��ӎe9��p{g���%U�#؟L���.���D&lk���r�Y�G�to�y6X���MYt��r���ԣ�K&K��j�۔+�{�7�!8�j�.$D��ȑE�w������6%F���n�n��a(\��=������w=��φ���+�%+�� ��,L'��ȡ�~l�c��H�w�Z49�$&� ����X�����덟�G�����N��H�!�<�5�0:��2�{����Q���S��tϛ��{Q���q[�.m��2������"�I�< ����{t��F����
Q1��Ba�����\����6Y�����-UB��۵,�>S�`%
�Jb���=���ξ2���H�xA�TLc�T�Za��9LQ�X��M�G�.F��-V����]���fCyn�W~�IL�s�(�;���1�A8XN^�q=����vÞ�J$Q�L�3}���lH�w���KB��t���l����ʹGGѳX���[m����GI��J���͔:�zV��Nͤ�Ie����<>��A�vC�c�.�WֲOf�6�hv6U�f ]��52ڡB��.>��U-��ǁ�g6��+V~I���8��|z4:�$z���Qm@�k#z�c����Y9>��<<��,^U�?Dq+��ND��e����>�ae_��C	݌�_�Q�#�v�2��z��	�Zhj��#T��,�P��SI�`��1DQr�I� �|x�Y�m�[sy��g���aȦ����������дf��*ͳ�OW�J��0�לI��Fb'S\�	�`u7rL��Ć�/�*��k�R(��G��ꭄ8�}�%�[�L 0�^&I�` y�-��[�=1m�՘)��.�^s�.I(�r ��T�y��Nb��[1��qH���`/�}�W&7y߿������Q01����tV:���
>�p��a \��7��x�'H�t���ɷ�B�UUL֔$�z�cxe���9���4�/r8�ܹ6:w8n|a��!��_M���f�	��.�K�E���8gk2+�J��?�-5ՃZ�ߍ��[u��ݑ|�x=É4�A�:0��)�V��Ь��b����o�u�k���i�8�M7A*U?��_ye*nb_�S���B�!��Ʃ[��j��S4���$�p:H��{H�pܼ�n����8�#��M��5a�UE���K��9���+�*	�����G�h��:٩P6�����*`o���k���H�o�A����0��6���A�4�s$^��a֤�R$$B�}yX�#Z7.F>�7I��#�Y˦������v�� ��.�9tO.ͼ�*�'�AZ��8"%���� �v��,�>��Vj�R����%����#�u��-��V���e��]8�W�F3��4-�hז �3i籄)��+����F}gp�?uJwW�r���oD;w�E-b�ö��SV��r�pL�&RM1 ɲb�]��&ԙ�I{�S������h�[
^����aA׻2X�g���!��HOqeԇL�~C��hc�2�ư�f�>���O��@1��\��1��x���<���v	�V:��o�h\\�X�k�T�X� W�4~��bR�muAA��]�=ja�,w�9S��@V3Z]����GƉX��'Sƪlֱ�x]U����<c�]�'
�����Wa/o��� 3|r�R�1��/ɷ�mM������IC>��~3|�:�/vWn�0�z�i��8e�M�%����d�(�Y�����Ʈ���K&��4��&0B��Ix�U]���']C��t:#(���\���R@�^�� �ck�aH�~�N��m��SN[G}C��u/��q�[�<׭��QB������!v��S����H��&���.�I:���҄E@v�j�qr�ث$�>���s	�,�G��B�='=o��k�����G��ո7�@{�Ez�w<vHF��&h�^��_��_�v=��%?m�t�������x�_����L�LY�ڝ�ӷR�4�s������K3���43"��Єߔs�� ��$��܍#�5�)^^-Bd���� ���g�[�48+n��������]y�x��j9+�gΏ�#�K�c��e5����cL"=�p�:�wdу������(Q.b��:�m)JFu�)��w�^u'xR��X�Eh/�dUx�G3�5��z�j��j}�RO�U 0�l\�u\���+J�C��6�CBc��XVL��WH�1��RN	D��� [��AM� �.%�<��KSiO�{ߛ�iVI��/:��4������������ws�n�96���A�d6\��^�i�5��Eǰ��!��H�xP3�\�Qۃ{�%����U��ؽ�����ٚᄉk�O՚d;O�O����ϩF+7�[X�O�Ȋ�3��	|g���X�����l5E�Y0%���a>�@A�mn=�7q�0�{�%�X����sQQ0��N~R9va��Ἧ�{�gs߂;�EC�N���g���U�����Mƨ���f�,�¯���,
$\S�(��8ݠt���a�+3�����v�������X5�=.�qq�k�`4Tht�/Vո�Ӎ=DXi����@ �F��ц�5� �K_����<v�QW+b��q�8}vxm�U�z0�e�je]�����.�Po���}��M�O�
��rQ�0����-��[�h�*�����z%��G܊r�=�l$@��]�H9?Ӱ6��h*>����F�3�F���G�2��n���f���Ch�v�j�1K�te�[Y.�/԰ě�?�J�`4B$)���]K��eh}���p�g4e�զLl�����C� ��W$��(��Hn��ك7V����c���h�o���DK�D<���L����$�&�
��mU:䘃6�����h�uv%�ҩ�"������ܶ�"�c|�l"Q�@J�b�Ea�'�*_���,�D�ži�q���&�Ƈ��y<��X~��FK�Y��as/u���3!�yc�^��D} �{ F�\xv�|ޣ����ef�e`��;~7w_�R���R8���S��L���X��0�)Ց�Fg���3�'�`�~|F´� i��A�}X�~���(4]� ���[�{����>",�s������ �$5ݪ�q��hk,��&�k=
����U��Y���� �b�P8rt>�AG�<�س����؈������M���=���]Zi\z��{w0T��0|5�WГ&�vɓ�N�A�5�yܸ�s�M;��H<��;�e9S��a�|���T�.8@?�a�������XM<��TV����f#3p��:�)��Ǩ� �^�U����Ap�B�&\Z;�.�' �f��?��
x����n�LZ����O4[��=@q<SI15�[9��V|�_�`����ٽ+h��#���8��2!5�p#w,@F�!*�|8�FE���$+�Z}E�W7�	6.-h�� �=Xg�ʅ.<%5�P$�Ҵ��=:e�,����AR��2'm%u��E��3�@�*A�,��ܵ���:����<�����x�G��>tV�y:��A�s��v x�mH�����3,%���Dzߵ^~�U~�2;�Q�*w.�U8����9/?�(� S['㜹4o���ŕ���=�wQ#�P��I	�Dq:������t��^xy�����jrNeؾ(�ql+ �!�*��_^��.�^����1A���2�1�m�L�	JvL��k$��RΒ�3��z�^R�$um��=���,*�Z�A���0���r�D�i�( ��㶎7,P�����,�JK��fj���K�����ΛC�rl`hrc����������JDU]�h�)���*ji�=���t�M�b��K�.7��i�cU�T;��%u�!���WR�>UV�-<��J0H55J�uʈQ����zXWD3��ؼ��/�-ÒG���Uh��䁇^I�Ϯ���J\�i
w�|�QCKOyv�xg�M#�@?s��yUQ��&V1/�����A�o��i��"��+��e&\���m��C���������G�w�73�&ᆺ	���(�=�J1}�³Ţs��ЇzP�T�Kt�O����
@,Y�$WG���z閩��Q�R��ߓ(QYު��A6|���(u�o큂��Y�]^�1��R�5ꑄ���J�^B�.�"�z:P u��v�<9�̑��������C3�"�7�[g	�z�����r��4?v"l� f�k��m�kc-7�}��G��m��Y��s��;v3����KC/�<�π��-��&�?-�9T�Ty���\"�8ך*+(J۰�^(��3�R���k#�>ZL�}��4Z��N�7Ύη���*�i�����փ?�/nX���/_⁢�	�^M�:G��,Q3x�я�H|���-�i�M@B@�m4��ri
��k��c~b���"Ø�����R�������=�"~|䁁-o+$�[�Mc��u��`���Ӟۧ�.�+@"�#�+��u�p�Po�|1�m8)��sUKV�B��07�_�r!��J�+0�+�G�;V����Mɀ
Յo�B����btw� 7��%�4���B\��sE7�y��@WI��K}Ä�i��Md?:cVg=���~`z�k:��a�'k�����Xy��}�j�F�g��rvv�#sG%Λ�6��CL��w3�H�zP�D&�)��ǥ�93N�w��0pY���_W-��Y!PkW޹Ȏ�Gޘ�s9���^���l����D�uZ���YჃ� �
tw�G�͙1 ʕ�������]d6�Q����
͠��
9�Z���Zf��@����{c\8�7
�� �]ܲ�ۓ�F��Lc���7�� 9���{�2lN�Ŋ�qIds��<�N���R�b8n�״2,R5��.� z����lb`���_�k�r��R{|�=ݵ�-��f��9�§?Q�Eo�:��¦�k
�6�/Sj�\`��;kXc�},��̞G��-?7�D�#g5z���"H�۸��ZY�.`��g�U�ժi\�oWsc�BmNw'� ��1��m'{L.?N��R��Ɉ6���M�<����_�h�x�5�W��P�\@:������*r��bV
N���Ih%���Id'��Ubhbֈ
U/D%� ���1���G���f�X
��aJ_`[B�u����օ	C�n�װU�%��CIc���cfI{�(9Nk]����}��8Kݨr�֪B�jb�8�}6��`��D����g��p���v�lMJRiH�oG{���'[�i�&RR���ʼ����"2�R�뛷m�ɕe�Q��v{!���]��L.
�� \Vװ ��'DQ�q��Dñ_x��L��4����*v9��J��s��~�h7��g�S��~Z�ża��(:�CL�6�{xHK5�2��k��b��ӱhN^�S6�[�P�|.O˺���H�;���g?�|ٷAGD�#�ܬB��
�v�o[��EPd^f|��E�|!�����şۙ��6P�*4��K&�-۲0�L�(
I��H�}������7]�r�EЋB1zr��3��c�9�7�qHB{iTf5n�uQ�\
����I�@ͷ;!��ʃ%\/�Oʟea�[�˺]`c6�0M`<��%P����������L����>���f�~b�ϩ$
�E�J%�p40�����u�������d���u6�Xy�qⒸ,&�Fu�~%��w~�A+Q��8��\��l|�C�9`5���Uv����BB�2Cpv&WĬ�*6�,�A�g���e1�P��Y2_��k"ɓo��2�츝uT��p��Ą}�)�z-�օ�8lVF����  hc��Ҋm[A��\E�+}R�nMA���e�*r�r�j^i<�B��쾹W�O�P�ʏ��>��;x�
�����̃D!�lr���/�>,[	��	�]q�
�qח��ĩى�h�����}�uS�1B	2B�j���$���ȑ�p}��1i�["�o:&m]r~�ٛBi� �j B6%/a�?��~���F*s��ߌwWI���%��3���5p������ٞY�ߜ��S���� _r����e-��k�h�d�K�����
D0@l}��pZy	�#�	�ƻ��q��P`��}���'dsN��b2�>�>�W�.@W�|1ע��1*@��$��nk��L'��X���2�Fρ{a8qt�y���o��}�:��[2��.�����r�J��.�U�H-�s��|�\�������3b5  ���OM˓���9�\���TA�,A$̉�亃�$i�R��o2�q�$�젉����!�8X��x�M�B�Z�k\l�L�o�=�X�^���!W:��uVL���]M#�+�|,ZV���#����ؒ1�n���b�A��<��a�^T�m!�����'����:�{/�+(���mˤ��"����1���]���UW��9C��Ml�R��.��R�_*	�-�*)�GoR�2_�ޑkU����u�Ŵ�w
��-37F�Ϩb�|vٙ6.��/�\,F��A����k~�U�QE��.�+8KGBOj�:J�K�rܻ��+$"�7b����W΂�\!��O��i�D���*E�tȧw��WE����4�@G��֥����u����h�v��w��K�I}
pO���Z�B�gFR��b%������v�.�ќ].�M�5ѻ�Ӑ鰕^ݫ$EZ?��N7Nt���w����_�ǔ�*K�4���� ��%�f����E��d���;�L��^m~U�9Q�`A\���"���bQ������BLX&x�~��J�܄~��NX���\��h���ȱi��t=�;t
�&e�p# ��d庎���Y��J,d��㪱��^�!s]�H��\t���C����43G�b��8nU��9;��p��Q�a��a�=�	��Y�g���{&��bI�2_�P�y\_=�}J�R����m�	0`�����SJ���;�W�O@�UD�7_���/@�<�={L�
>S�sd}���A����!)b�f�sQM7��4 A�=1�6�ל�lQ
V�$�Wk̆��4h�?��=I����r���1�$��X)0�]�~@7�vES��?q���D"x
[q�l��v�	���U�^j�5�zO]�w/F/��ߢD��q._��3M$ޏb�&)Ҏ���B���<�J�f�;^r9�r������b�f����)�x�8A~��2ֆ7a0��km�)�d�V���l*�#0��=.���~*���W�q�h���<N��ߜYw66:���0���I�r�kۭ
B���� ���ߏ�J������ɀ��_.�`f���/`��t�� �� 2���}��;}���V�����zp���%�%E��C�LHa�۩A0�ɻ6�� �ݵ��_C�	b�G��j��M��o�P�6�`r�(���:���2��ꗨ8]�3�s�9(״Q���֔�����9؈���J��|��}�KÒ��}Ԋ�-�4Q��L�$�r�9[�0YuO����ohfB�l-��b�J·s�a��m�y;;��܅U�3�zL�TD�>���U�Ui�@L ����J,�m�WO5���F�Z���d� ��0��Y"��P`�h*h���M���`UmJlQ�s��m�g�7�mp���N�N̚���)�>��pH�x$K��yV�������4!�9��R���.hI)r�b��R��FşLʧ���"�@��4�.��YЃ|�K��ߒ���[�sk +��Ҁmf��m��765�0 ���<��|�`�|�������z^��{�q���G�ѬoI�d��܍�Q���G��<ls��qr9�p�֡�VP�G"��^O�#�ͥ����~��<\!�[ȑ�V�p�K&�ה|�׃!E�x�I�Gu�2Gh��}�OW�}[���ܕq�����.9�ȣ�{��{S�9/�B��5��K�	+�� <��A�c�ҙ��>\N�,<��;(��?�2�]���6(i����&�,��L��X�7�x]Z�7Z��7D�L�����B  �t���5�Z��81�Q�ǒM�,������P� ��Y����6o�q�E��4�����ߣ���^�SQ��tX�b�yW@cȦ�|�N�� �u
baڕ��ܚ?V�t&�i*�Ά�k������?GJ�q9�%Z�"��b������G�2��:�Z��x+i[��~hy�L
_��]�5�{1�;�8���흡ѻ���!� �ex>�p�"���e9��٨2>~7�j�.bUR�s�g�f�t�����w����5\�T���0�K�L�{G�a���Y�1�)څ聃���݋���j���b쀞|}�G�/$xD��"e\�Eüꅲ4~<�V,�H}Ќ��+p�S��۾��ci�d���`�gP[�x0�[���T+�k�ʔ�ʞ�p�UZ�ԍ@')t��~-\��"��y"�(O�%�6_����� #�5����,��N��Bs�נ�8�XG�:X��D��Xȳ���i:qʐ��!=�lŝ�������w<S�f�N{�ON_��� ��E%A���>����}0�����v��L2-u|-gG��w����/~��f�сk�	�:޶܁F4���{@��l`�e�f���v���2��ĺWA����e���@:�ݪV
�fFI	C�4�7���7V�?R�Rq5�Ƕ.'1CJ��u�q���^�1?���=aOz�w�-���}�x��O���H�IK�)���;�1�JSW#��Չq�-36_q�m�'�n��~bWAo�a$�N�b��G;�1>�+�)�i֖A�W���spo��T/
����j!\����TX|ڋٗ
�ʫ�Ƀ�:j�x�x
�k���m��(��L�?zݨ/3��xפ���|�͔JL���}QIe����^�	�/sE�[�,���zi=t
D�E�XKhA[3��ޅfJ�H���c<#Q[��ە�o~�F��Z{�<L���2�,�n�K���`��RD�s�B\&|�9:Ϸ3x0?.��'�S�ކί��2=k��:��N�{��ڶ���Q�n������Y&~<'�ٵ�%��Q+-���)d�]";�ٰ�	�|&Ibl���?�2O�H?�i��7�G�s��U�cy�)7�?m�̸\wY��!�cӇ:��ֽD8!�҉����S
*��k�Yw��B��{��cZ�Ş�t��6�zD
��-/��Q�%:������pgC����U� � o��<:g�!ӽ�+���t��Z�����h�P�"M���1��т�@� 6�#*�0;�lR�"�'� ɰ�>;z��P��Aau��@�����i_��(�V��;�fٴL���j[�r���)�_��K�}Ə�߫b	���B.@�)W���(%�Æn%H��}ȭ�kˠ� ��`�eu�<]�qm��Ά��G0��.}���Ri�Q$���km1�e�t�wiO��<����j(���yfZፖ�st���}��h��>=ԟ���A8L��>H'����9\�R$��H��ć_���ŴL�GO�@7�˰�j@���ݰvhc�C�8��ݧVq�X�J��&��P�h\��V&<���-$*x�2�� �����g�ʵt�ޏq�aS��C I�{٭��]û���,��i�'[3���ַ�lNF�pC�>$�0�An�Ʌ<[K?�l��$Q�7���E1 j���BB� ���1S�?�{zVXc�
R� A�Y�մ��ad�gD��Y4Z�@�� %am����:k�k1d�A��r�R��f��x����~1�a�zu�T{JVZ�ڐB����L��!Q�3��4X/Np_C�hIקWU��01���%�A�nԔ�=�1����x������q�Xڻ�>��  ��hL���հLHB��%�P|Z�u2S@ۡ���/��+E�A;�kڳ��΋̧R�m�ɀ��/�w�l��YM,`�c�+6�PqZ�} yLR�փ���)�sKcQ�*�l�\qQl7x��D��P4��oL��Q���U���oC$��k��݋��Qk���Z���˴��F�_��>�
A�ﱃ�9*�ƪ����	���5��b��1�w;��˱v�V�K�d~sn�q�j�1S]����R���}{�5����6%�"�2d��ԌX�V��
�7mj7���'��ڬq)Y��o�$`]zZ0����J��yb�y5�rm����<1w�_�>a�n|��\0�ы��_���ߏ l�)�$�M#�7�8B�y-Q�r �����؎�)L�3$�	.��KU�
zr�,�L�Dq=�O��l3 �O��A_��T��G�jh�jm��Fڽ!^���)a��'>Y�)�
%�]s���W�M�q�%��)x�d[��`�u��u���=Ĳ�&]�T}� s�U�&f��� �F���8�Y�^�J��Ի?����Pcn��	�:0�j�@ؕ2��!i�nUz���ϭCk��1ұiz4'�av��!�LX��x9��u��q���?��b�`J���`e�R_�-���ӌ:zTv%5W�M+��I�U� ����\�*�ބº�������R��/���9�vꯕ�&K=2�,�Ơ�Ɛ����w�d���#�0��؝��},x]���'
���a���J��~�~����^��V�!хl�^��ƂN�^�v�R���Q(��.��`�y�L�����.ix!ᴨpI|p�7�i��+����ˆ�K�K��> H�X���d��d���G��9G�σ������	�|�ǹ����Q =CBȱ��B��%I�]ʶ������]�~��q3CU�f/3�#2��`�VWg,??��a@�_�����E\�QԲ]r�(+b�>���C]g)�����K
�&�N�g�T#�-{�K��bTg��@���&�����;�M�^�'���]"�]���s�k�S��rP���`x��yMM�y���n㿂8��|���]L?�e?���u���"�<��V�rd��Aj�{���n�	 {苘8�D������{��@���8�פ�/fZ0�\r�v���,�����R��_�2���C��!^�`��6�
D�X�k�^�/��45�e�0��"��d9'�]�� .pl}���S��M ����ݠ��#
^���_��C�9��oYj�A��ƂaLՒL�?4*T�@�)����[�u<j��r�3ϵ��q��'{p��]�z�qƴL�3T��zҨ����3��i�����eDF���i	��P�o-�'�W9{0RQb1��EF�Ls�@|�P2���u �������6���"���&6��C���p,]4 ?��k�`�����E{D�O��E;)�^�V(��6t��3a���q�!�����u��'ޙ~F]Tqƞ���S����Gg�����[k_\1I�3m�����|����Л�&�O(N�p:>�`%���a)������$��G�[l4� _T��e�nr���g3�G��W���ME׸6{p�&���+)w� �B�䢨���5�֩ͼ�-�[=�@@ZAj�����<������{�ᕩ�.O����lt�#�s6&�� �R��؁�1�*�ǿ)�	�wK|"��e����7.��Mg6��~�d�_ɡ�d6HGS�ӕ�Ŀ��i�UToc�zų�RY�Y��
��K�F�C�ECͩ
�V���F�> �15?T�~���8��+Q�������=o�\:�uuB�r��e�������E��d�e��%����${uR�S�3:u늨 �����RHB��	}+���}�-/Z��-j�+�0��L���[n؎�<䰮O�FH�3ؗv�1{�MLMM�/�#Y?�b��0��L_8	i��p	m3���F͑*'6>ã|�����M`+�KC�`����,	�B��dϢ��qP������}���ͺ���K�lFs�fY�݁�F���l�/
c��>��EnI+�.Hoa���/��_o�}�,pW)�kB��zuer+��E�8�<�K?���z
v��ː� ���I0.�"�"�Y�TS"q�|����ݍ�ɤ�X��W�ض�"	�9|8#�7�<2�6�(��^z4ʳ|��5�n�}��SQ	3ʤO�+l�&k�ArY�ꝟaP�̚$���i%S�һ<����"�H�@BT�E���z՟c��{�{+T�M�yY����m�l�)���"��%5�nW�<�K���\�Bi�C�bw�M�_���Ux�f)zbji&�TG���0�/�{�mH����%�����њ���nh�*A+�#���p�U���+P�� �Y�Eg�J_��?%�o��m> 4&�8�����)��"�bV��k=�6	�X YO?cw�ѓOL�Ձ���^�k�F�R}J�8�0U�G(�1#i큻ʃ>8�Jq!��`_��#�yM��
�Nv� ��P�9X����XX�"���	��F+�o7!h�1 �|�R�
�`x/�;`���Z�����Ӗ�S�Ŵ|t� ܾ�v��mMO7?l�h�b���_��o{��诓�x�6v*i�r������3�t�9 �E�;��~�5-%��`�rkÏj筁�UYq/%'�!���SL֧��(s;�%���:�e!<��y�Y�����۹1�����Oq�c���A�L��V�;ŭ����ՉI�e����o��	TV���t�v�\�Ff�.� ��y�i����8x3�9�'*���T�����)֦�M�wҧ�%���vFXN+��\���e�W�Fi�ͭ����x틣���]ˠsn�<�fh�Ji���Dm����u���^�to���%�
0��e�E;	��u8��%G�g��W��>���7]�X��n]�;(*���]eV5{|V�s�;o����	�����Z��P��s�}46�in��"*@���V�x��|lS}�C�ch�]Xs��c�=u��a:���֭q����L�*?v�LJ����,:�[˔Y�D�~.��c����Y䣸��a�x��ſ���zO��q���:lE��9� 7����-�C^�M��sŲ��YA3����쓭+��~���mT�`��*8he�U��������b�l�tUG���N�"wqNh���b�|Qc�d]�߫b��GՀ\WV
%c	$ԥ�7wWD����n��mX,�r��e<��P7r�ϟ�0��moݎ%�=j��Z��H	�o�u�H���4��P(�|B�￁�� �W9;� �B�΃<���@�͕zq�g�{��Vy*!����QXQE�{A/s��Zν��R�&��¶��_Z��_`���_��$�w;�7���ֹٮ��(	��>�
�u���,o�ڛ,�����g���<����\3���[���z��ˠK��غ��n�d�qz&ؖtD�.�pC��1��ɓ�n�G�|������_�Y�C�܏\����4�Ɗ0�����T���K;�^k{�t�ȍF�Cl-T�?_:��~�N�����BMa1�{�Ub`f7uU������
nF���>�fì��#�����Me��Ӱ���ʦ����:�Tkv-�Ĩx�n�ʔ�9[���HeQ/]{�w�WM��{�d�HL���L$P�2K��Pf�
��fX�}�ß����53�d���|wV�>rpM�L����j+|��+�J��Q!�У!z'���?EX�`< �kt8�s����}�p�<�nCm�)���y��Y��VfrKs�bC�� }��G/���Q�k�/7��0`Х��b�Sޟ�v6O�L��Yұ�I���t��Ph8��T��-�gLl��7��U����^.��RBk4���MSAJ���
I_��c�S2�a=m���>�KTXO�m<�2�l�<mpkevpU���y�^&��$��ͭt�Dc���o�^�[T��m�ۺV�j�Xi-��>L�0fY�����xư��z�+�g���U���ܘ֪F�}`��[��%p��C��R&:?U��8֗���h>���2�9��__���vC�-+V=gԓ2�V�57r��1�[�	Un����o�F:o�7�?,57/)����"�\�Qה9d�	��	ȃ��Db�P���g�i������j�T#�%�
+v�~�0$��� 
��aVh��tI��T��@55�[���`2}~LG�p*�w�z+?$Pn�d6��ۛ�!�T��#����CPxg���!p���s51��� l�Xa#^1!I�[g��ޣS6�����@v��/���b�iz e��V���N�yO��J,�[�?I�W-��\-���;@����֔
D�����:fhCLs]�V��׃�({��%�uoE�q4k�qi<ˏ`�F���z��D;�{��
���Un(�~��c	��y��E!!�}��ѧ{�.�&:��^���sE��"�G���A��2�e�\��j���Q wѬo�?<��;�$����m�Za�#j��6��i��Z�O<�{W�0f�Icm���a��WY�����=�X�h����=F��x�vz����;;�w��_Q�2��.۟Ǜ��zA���}P!���Q�K�V͉��-���+C�"��rp��Q��x�m<DS?��S{�Y�,�$�seO�ɹ�y*���P�m�d����I���[2���B�o��XHA�%g���Һ�Gw�Ղ��ߙ�hB{�=��K�(L�3q��X�у��G'd�@�mi�ֱ4�!1�l��Be�nD�v�y@��n��C�%ld��,u���[O�eՆ&U�c�Ađ������s3�j�ה���z���[��
4�q1���>����rf�_�wD�c�Qr*��lxq"dq�������M�.Y�kMAK�)A�V	�Ә<�GoBq9��(� E$���$��.)�eL�$�f�z���s'v8��!���h�GD��A#{`���Ż3ݹ�������)G�ۑ��M@ǘTÜX��!d{��|�h�G
�����y�t�W�O��!�m8�$u�&p� ��;�ƌ�z��+� �hE�i��JW��(UNk��1���N�㓵C���i	:�q�,�����J�QW< )P�\�˶���y�Oh_��n���������T�`:~��95�0�h,�P�#_�i�o��p嶗��
�1���Q��M��͒69{�y�;��4�#�br�������K���:Dvly�%v��|��Ù�,��[A%���0���K��Y�?�pEC>��J�:8	�ށ�P�̱1��Zٞa�N���\�bQa
��b�ƃ�:���3�;T��=���Az�i|����}12VR����3�g#�l����$F�ݤ�����kc��"�K�45���Ǚfwʙ��{�n�hE_��S�9T�Y��ry� ����%Y"�Ղ/�Md��1`f�u�i�7��r��ux��� 5���5I�BRc�
d�NBo����������t���8��B}	�n�Jl!�ʙ���I=�W�ڡ�o��?�l����}�8�;i�ـmX��i	0��u��^8U�Ρ�x<tZ�#�$������oѡ%�Q)�ԙ}~x�t�����X�s�`�+7���2��Q�'���C�}q�_o䀭��5.�>*��<O�P(�vEs[[o}�j�H6e͵������[�|�!;'���QQ�s|���s�^�@`]?ޒ/j]1qK#��%�pMa#B<J\6һ�J�CN�?
��	P1�.$�i)���`��� �h�g���l{j2�"{U����a�x�%J�B8�F��e����;e��UU��&}�=�	�Gc����cG�$¤��m=��X�7$n7�247�E�CVϴ�Yt��E�{?�%%�9@q���")��I�G�Dxr�}���E�~�m�.��il#\���O���!�M����x"Nq����C��́B��e��}�i�t�UC�����חs��[ې�IΙC9���HR�-J�ZYY�$�jZq���fg�%�.�̙�s2Ϩs7G����O��J�h��#����z��#���}	u�-�w����d4��黑ů��'Ι��9��l�${�"P4.�-ȓd1�A�ey�M�tcw�[47�&�b";����b` ��z����u�=�숼���A�W�t��v�V9f��硛c�̩ap$$lC��^+pu4�/�)�ԭ8jg�>sx���Q����^م������q�i�%�y��`��p��2fn���L�aZ���F�0���x��n%����^#��������)kh1�y�q2'��(k��3G�@wX��ɂ%��VRTor��L��zq|bD��@c׾��!f"����|:j3'ӣj����а�-C^�F��S�tPP{X$��%IR���VK����}�YUO����dc���uǴ*��ֆ�-�l"`]�=$s�!�m;�ɑ���W*����NCV�������z������|��^�ಥi�1i���UƼtn��V�%ϒ�*%������l'���,�@B�������˄^+��l�&s���	��̈��1�;W4|V߲��n2��J0!�
�7~��kX�TWL6sOx/>T&���v@S+�劣�>�N�}>�(�����
`���D����{�(:���HF>��&�B�{�m�D�^j�IW|������p{PK��#��������盥�Xw���\�P�h�p Y<�§��6��	ŝ���?�&E@�.Y��ą%䍍�a;8�\�ʗ_�zQ�3[����#^�^�ZDg�˶�|�����Q̿����܋k����@���dq��N�e6������;�?�ن�zU4Zi�<�Nǹ�g�q�&���;Σ/��Zup���s=^n�X�Ǻ�i<ڃ{�^�g�D���O��Zt���i,�	���Q^!q���p?e�ޱ`�~d��zD��bo�A��?8����]�>�@�����y�L�Y#�S��" 4��ik�s�1���o����!ȝS�"F�Y�'��]3ܾ�/�Y�:5��oD0��b�PJF�X�J��ze-�� �����G��á�;��M���T^�p��ذB���R+�h|�M���ޓX��L��^�W�.�$@?�Ey�ǋ��3\6��3ޝ����$�����;�ڱ�F��J���D�_�]�U���o��zuP�)Ǉ
F��[yƉZ�VH�j�;���^=uw�ݦ�1� ��	�u�`�M��l_��Z٧V"�R$��(��!ֿʥot>�����.Vy��@}P�?bz���|�>�\�y��ʛ�#���̬y
1�0>�?6�u�R��SI&_�me�ş�n���&���O���j�é,<1�˓����!����#4�5�QҞ��/=ϼ�YZh:�(��>M@[�|�N9�J��xn�|�.|���2}���:���2Ni��ߌzM�����RX�z��M�)���Ey!����FXa�n���%��>��y�A�Y�h�Q�E�u�vǶ^&��H$����ݞ�!�V@l�M���@�j㶰@C�>�R���G���І�Tt��//��AU�#;o� �-}ق�&�ꋮW�޿�a������slz�d=�0�'��(V���ฮ#��i6��E'ҍ����)�&S:�7�i��?G�p���t�3���W�@}�u��ȞO�ھ�)Ze�PO�����~]�(���8\Lu�)�e��g������⌤��L}kcJ�;Zn�z�2��]l�1ew��6K���-PK��jsJ���bt��*Q�����V."��%j��8��<tPlM��Ư߶a5x��+E��i�G���o�~eJɯ5��-�'6rI�݃6�U9ky�d$^1�r����x��CT����Ԯ��L&e-&w�%�E�(�e}z%W��b����k�Կ%���� �{�&^��g�)d�>�и�_h,0:���ݿh�������ppz�,��v������ /�K HS��hF���HB�2�&kR�k�8mr���"��8����6V<�₢� m��6����*ג�cH�H�XP�HG� ���U�KR�Pf�.��/L���Z�����Ql�ytP�m�G{�U��8�Vs�\$	��`_e�������Җ�f�m��8�sS���?��	�^9��f�~��a�z�1��T�a�hO�̓F�.Ξ"7�e�6�;P���,�~#=s�/I�O���.��0:�4s�w������I�t<-�Y%���U���P��n��^����\�"�L���f��#Z�̓��������W���8��?s�t���e 	B�Z��_*�׭༄�͒�+�-=��5���u��)6���7�� �O��V0�D�ak&!:4Z�-5�)�:�Au	q�J�5��]��YVěE�%�[��3�7/5�1&�t9@i��f���h��u�'4��'�V�>GƻH\�Ԥ[f�o��o�)7�W�\�c;W��v�Q�t��Z�ݍ��1"�C�2�>���h�4�&��%�	kw{��_.��߈�!s���3Q(��J:��{��?���{W/��a�T�P�-� �����P�P�.D��|�kV��8m$J|c�.�S
@f9k���o!^��f|��b���Po ����=&�6%k)f��o�y��=;�������VR�/�>��<�6��4�� Ff@~�Nmї�3���粉�8I�0��{{�o�Q�G�����lݺ%=�w1_�$���	i5o	y��G��O+F�l݋�hY�M�+�U{��әt��7a���Y�s���|���?Bq��2Y��񨻓��Ak���DW��t�7X�3�$6|�6�z��?t8��"n`��.���gYJW�Km7�� ~1��&���.����K��t�������o!M��i��y��n�Ht1���\�7K�WëZeB�(z���=�"
N�|W�,���qE P�5�`E&	����gY�4\!��'�FeH�;����\��Zx�?��]��Ǭ+C�V�ZgY������t�6�0��Xb͝')]M��~3�]�˙B���U��1q߆p�v����?6?����@��w��t��b����c0y�W�}>�۬a�I�>2\Fpа��0�[�4&�l&�N���4�6\���=�Ucx�2ɪ!�������s��p�D?�P����}��X���Kǣ����&�l*k"��j��{=�H�jUc1����篯J��q�{$h
�'K��� �<��$_��{ߺ�%0�"x2(iu1�tㆷL^����)�&7Ɖ��hh�r>�6�օ���?�"e�ף l�
yB�qj�5f| ��aX7}�o�y/؅�!��g��w�C�!���:!��J^�U����j ���H���uz�{��S��Q�2�1��9�ڕ�rk�(�8�@��	����n߶�-�z���%Wl�&G��%�l�񜄴D�>�?��������^�q�zN�����a>6&��kj"$�6�٤����Ir�e|x����t7EPA�$�RCf�k��V,!�T9�xo����T��޾G��g��2�k��O�[߫SL�t��o��_���%�z�y�;��(��h��l�S��D�:/�ht�N�,��4)�7¬q��6�K���
�$�ً��1c=�i�p}�x'Z��*#P��"���q�ک��BѲY��Ҧ���zl��,y��!�*�d�D�6(n��$VXNA��-��j�聍'5}�:"���p҅�#���`E>�L� �X�����>��o��TR��K�SxH!�ܣ���>L�mU�tw�3�b��/�Z <��+o)�Rb){�|G���N΁[�3�������%��ͥP����]���&�8�xna���ĕ��=N#⮠Lb�j,c��pdP�̊S���|��r��
ߺ^��(�u�A�n����	�Se(�O��M�3�������Y����/G�u��Aw8T���؆�s�1u�t9��=���<��(p��X�@>��\#��pK��������0hWچ&�?��������,k�ߵ;����ד����>N?�z�K,}J�`��O��|J���]�x[����	�$1L�K�Ȧ�=\p��0�y;c��_��]���O��6��$�96$����}!�)5��.7~�B��a�N�2CX�urH� ��f
��lJ+}�C���X�XՈ҈�����Л]ܖE�	�g�*�^T�,��Q<���jCr)ym�҅��O��|�*�$Wזv�m���?�n��S���ɉ�t	�΍�5L�G�97�hټtF��am�&Y�ZE�6L�~���B ^0F�ie`�!&��W:��D�貖�!L��N#.��k� iM��^�dPA53)�f4�L��
o��{<����a{4����بoC�w��S�m1�)TXg�HPU���� �AA�t�d�q�^d�Iz!c��ܭ?�Z0G�#���YEr�S�_nܟ��&h#<=���k�\�Ꝕ?4Dh�S��9m������k*˨���}h9�<w���+@L�J��}��p#�<�L������z�pK�����HA�ߨ�$8r]�^9t9��t=��J{�����,�P�����u:�^+�Oj�D�2�d5��g]N�p%Q��;�`[��a3�o��P��-�6_;)6��!����GKs�!+�Zl"�/����(g��k(0�"��a �ޢ'��1��..�U�S&U�X���j��!?>�!��B*������ԯFA��諶�\����_��t����-��r#�c��,�#5ֺT����=��V�h1Z�\8�c�;��.�)���Iޙ��O��8����s�$��sEp/H<lh����l�������%����A�M�'m+������ؘ��$n��P� &>-��s11�0v�P�[��a|��)H��6��kNw�j�?N�}�������;;x7�K�WAQ6S����3Hs0�;��?7
���6��~؍���mƤH�:v��<����p�\y��y�����Q�t`"�͈��R�S���GL�o��� �ճ)A�%��^��{Pu��#�Ö����ȼN[���$�a���iXKH4�2g����l���C)F�QYBoOtV��u[�rC�
�r���W���ok�U�fȡ.�AphL� |�P;�̖����#�̓v��3L���e�lrb���c���8N�<m�����M��E�tpL��Aƪ%�R�	���+�H[-�E�(Y�&3�0қ�z(Т�.�
��s��IZOn���ϟ����r"���d��gE��֛�Υ�o� �.~��cfk-����VZ2��R�<��<&.�zGV�}������>~���F���E��^��5�R9�������������}��u�4��z�aK���
s��l�:��i}�3�2��v�1~��1����8�9uLQ{u�2�,٥C�CD��>In��?	�/i�.�/)�x�W+w������
��Ut�־��u�s��9cP+R��ȽQ#�������V�
��f�qtk,V�3��X��h�9�`���E��@��ݻ1t�(��Ӡ�Cc�|"1�tm��'���4n[b�`���1���$
�Y�#7���}Z|���ʰ77?�|v�
;M�?���2��V|b0	�H�
���6���+�g��/��5-��]����lLC��GX��>0|p�3I_�w��Z���2=h�豨���C&0F^�3���%�=���ڻ�|�j|7�1ï�͓� �(��AG�d~;���N�x٨`��43RVmU����j�W�^�i�$ �*�69�ԛ4U���& �1��e�5P�,�;d��$Wq���!��7��z�z�[�������Yg�P�"�}W/���ʒp�99����d�؝�84�ҷ\K~۷�3
6E,ѩ�c��ثy��������FF����z���c�;�&̲G�v������\��G�.���v!�h6�5n�T�#��ZV���/!W�d,&{�ax�H8k�����o
��8���"�6º���_�,����)'�b�İ���b�M\>��:�d�\S�z�5G�ܬ���Ϲ�{j]����/�	5�ɋ0.́u_D��/���"�^��.������	�z�Ăfk� ,t�:}n؍�6H9�}B���>���L�D�|k2����%�����?�K�:_�y�i��T�Cf�@Bu�-	�k\�F�O��t�v�t˅��mZA����X�=�w�����(7����B�$}wE��E�$����3�7�F'O#2�՗���'���`�����I�����63�dPq=�����s`��J�9�Ļ�E}-��|�æ7���:{z��AWY�-���S�?�Ѽ��u�a�G+����.�� l�x��>��g��Ͷ�r�2b+Q�a���ٴ1�*,Q���x����Ϊ�v��ຂt��|e�#Z�鉙�w��Q�QQ�WQ�I%H�D�%�����4�?��C�������ap��o$+��{��aH�[E�Ԛ��������`�d��n/U	� =iѲa:�x�;D@F�ML��\��D
�b��E6��:�@�5��p%���.�bK8�`��6�ZyJ�#��*H��<�@
A�$����h������&g�ܪ2 K�a�F�ZkF�l���OL��:���#�%����I�;�}B����_rk��FG+����q��\�r� ����`�Y܀�e����}WE�������&�m�*�tv7	5�������%w�L1!�,\TD���j*���&�*��T1�%������>8t��^m�|� ZSQ�����M,M��8���#fɷ��ſ����]������I����Ox�D��������h&E���J�/��O��C����L�݋��EF����j�����?��`�ѯ-q�]��N�݃��$�PҪM�I�}˥F�숏�2�X}�=մ��Wa�)	��w��$��Ss�D�z����L�t<�4�hފ�U/�œ�ͪQ�{�b�ާܘ���U[O�j�M��h)���z.�4��Ӝ�[�(m��@b�dϽL3����N��=L�7S-��
�/��vr4Ut#���SH���åΟ�/B�O���|	��h� 8����U�����*�㌾D�6��5�Ōm�k�j0g�|8��+�O�b���,�S�E��<� Й��C���S��WHv��Vqe�Y�|�	-�hr�e��8
���>6�e��:%�_�X�}��.y!o��[��9F���ߕ�eNྤ\n�\qX���U�.�߉��3�G�Z��Ɠ��G���B�^v����nB����.�t�T��\�uy�*�t�����]�>�E. :���)-k��9��ԭ�A{�V䍛��cMQ^k��0�T�LP4����)M'����T}K?���
���;�`{j��hˎt
�C���|����fmy�F�L��"mߖ�=���	�Rno-�M��
ļ�:3_���Y$�,��ᒬ��?%�?k�ӿ�p������9�NxU�8�.p����k�v�o�؋qOlf��J�{����u�1(ɫ-{|������k��� ����;v���΁)�7�&��Y��ݰ����?S0�셷��6�y��W�_{���VCn�h#��x� �a�����y��F"r34+=-�@��_�ϟ�L��eG�-=����	�� �#�m�Y����m��u&�b���?�i�����ғ�.t��{����{/
��Iǽگ��E]���7�ǻg+d1�Ue]LL�{]��Ř�/��m=O�獞6�k�?�Rڝ�N����Ѕ���+��ab�:�q��b'�����i!�m\�Siqꨙ�ym?!Q	�˚�}�C�c薳5��J�~�������?����ͅb�۝J��t�)���gd��������� �0s�� �˃����p������
f���k�B+<�?Fal
������W���;���Ni���@���4�	d�$e�G*�'�A��.[6�*]b�c
,b��!$��C
=81��1�=���1�%v3� 3~�T�
��D�VU�,�B I�۟�"$�Ux��?b��~��z��&�x��r�L�񸚟�X}�:m�)���)��2��ӵ#O\>�|�O0�x�o}U_I�Qp�΁7��~زD9%d%ir��E�B5jN��	ӽaY�A�a">[����w�?ë�SY�/gF�qD=�������<E<sP+����[��i�k;��l��v=%��_��C!I��$u���{R�b��]��__�_?�L��~ҭ**�q�-��c5�<�Y