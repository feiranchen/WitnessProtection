��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX���6��E'r-"A�ײD�M�����G<G�=����9�qYq�~�x	zK6�L
�I`	/�*�!�"��nM���t�0lV��eɅI�Yz�l�i���И0�f��G��=2�����46Y"o��X,Y�U��Z>5NX
�apV����8��Ӕt�-͑z���ޚ�D�
H���[��-��>/�G��s�%8��X�-��c�?D�����r�_-E>�%�-�Te��/��ĸ�[���p��DA��WO��Dߤ!�~�e03�4�?M���k����-{������탾����\�긐ox$��.�O��������,(Y����gf�E�=���y傉`�P���i
`j��RW]��K����B�K�`(�y�R=�>p����R��>>Ň�y���ă+|k+�s�8+h��X�V`��K��+g����s�T]KG*Ϙ�O�P"JNB�BJ �w`à����9rڵ����#�ӌ.�] �hS�}���ʽ����ńD���� ��휡UM�4�=}�%oZEv=FiPx�K�0�/qR3{4d"z�V�e6����1�Q&B�g:b��4EE#��I�r�0�b��V�l`����5�y�� =�oP�]Ɍ�:�o�"����.�C�O�����z䕡�lF�~1���$
@�2�+�K��Ԛr(rc���[��/�hw|�Zi��9�|~$JL��j�#�oI�s{`��{�.�g��*3���z�#N@��w�J�cU�}����zc��e�!�bƟ����X �p��jJ�������3�a��WE�P����Ft���pmp�Ø@c�k��m������F#!P1�h�Z��!'�>�(�'Eɥ\���7��Y-���M{G&/ �1�9h�\`ë�թ�'�.�w��]�Y?85.�J~'X	c굺��CH����eĸT����# �������K��}]���<L~}L�Lم��:�
X\�H]����w�gM��(Iϖ|.k�x:=<��Â/!�I���S�{;���^<ʆy�;��+��ʐ5b	vo=�Pn�������6[�g/�����_q���O�8��pj���]�vg�0C�帱����>���-�$+,�C8�Y�:�O�T9�����y��'�!���4���:���]�!���^���yo	��G*
�'���S��eVG�%�\#>nqx�nE����l�T?>%-~=�۶�0$ui��h�/`�t��mG��?"B��0�� �c������� #��WV�H�ph�Y�,�5?�LQ�
���;���N$yJ�zL�E{CC��G8S	�Քɛ;���ޝ}�e�'�b��Gb�sbL�0u*�7nM�xWr�}�K�-D���T����i�[Q�-��J��D¬X(�aTB���B��^�'�Q���$i�x�b����6N��$u���r?�$D��z��[�.5KV,���i~��0ݮ���i��8�r�`Ʉ�/1��7�u�W:"��3���X^�����x/B�,��A�w%�7�>�5�{�(y����$j �ϥ��W_-�q��s�����#{/yk�Ҷed+�A��*�r�i6מ(Xd�`BiWW؇�����G��f���[�x��ܚ##2�����}w%� �nwΕ�/��β_%�t�A$��wYvs��O"Z�a�,��Z�t�{����8+�	����ĢʹNA=L�ό��]JS+�d��a��y�^*T^N\�X�E���`�ܠ6�E���Y�	����|#��Ϩ֯�^�蛈.\�Ʉ���������XT��iO@"Ϗ�^'^@=�u��[''�쐹��Kp�R�x�-,F �F�|u�����nş�(���Ϲ�T4!��2_�j�`~9/V+[
�%�Y�� ������QW5����GB %�
���s��G
1\�˺%n�dSe��Ht�q|Ӻj_�������μycV�%����K*�;}��t!�ָ�,��S����%�L��sp��z�c��'l=w�p���(S�zp�:��Q�K�y�1�a�d��vq�蝀G:w@g�sD�F�3�p&FNlS��#�ΝO��rp~� ̠ʎ�c�뙤T��ó�%�>Y{���P�_ү�	�����D{N'
��='�^}N��H\]���6���Y�(���t�|Ыc�l�O+g��(��H���G͍|?���t��2U��c[�T�F9�/�䳓�V9_w����ߛp�#ae�uah����L<Bz��1�,5ɕ�������^�[��
�<)펣�\�]wWJ�dl婑��:i~��qNM��*N}�s��H�{��	���-t��j��s&�tk����*����T0n�����Z?���UĀ�F�Q��w'����Mr{�C�e)��cؔ���bn�r�\?.pM1�u
4���}S��D44�*�i��v*H�8��C8H���f�h3���]A:�L�y>~�����Zb�V����C����vU�,Hc�l3��@0�S�_�$fǱ�#���-�$��X���Xx�!��P���;F��"-����ɏ�_^ԣ��+���X@1�2|�x3���R�l��ɑH �G���Q��ݟ��(�Z�2^�m������!��.
c9������Y���Ԗ��2d��+�2�X2���!��]%�a`�'�SednAGL9��0�V�fW	�ǧ�,�N����oƚ/�X#U�'�s�73����d������B6vFoo|Ý��ǃ�TO��K�N�c;��c����9��9+e{O���]�҂	n�x�h8�����%�+!� �g��U@s#"s��·��N�����Л����@ˑ3F��%��u?Ɇ���ݧ�h7�Q���$fJ���n���}��ɛ��7�r��0K�e��{D�0.*�_Fj��G�����p6 ���\Zc��K,����[�X����hz?igz����o�~�)A�4;���P:(���A���f��/�C��|34��Y��|���1*I8�V5�Gn�!��V���s��<X�e���M�jd�.�/M��S�K$��_#���.ϋe������"�dR�a|{}��XH�Ma`��"G�m%<6S�P�z��D䴈��L/�6Eg���C!.yG��ر0uV���bc��L_1���
�()��{���3Gif�w]��O����0I�lbO�]�@�^�0B���2]l+�T�D��M�D�&L/Ir�"��D���|�܋����rb�<�^k5������� �P��]2����p��IQ����� j�G�d�� �璦�$^)������
%J��$��--r
�
�x?<!��Ä���~9�sq�.I��utr�[�X��0�_y�|������1�
�j2��z#�T�Ԕ��GU���vV$���P���m��sY=|xi�]|!p�M�h���2#ã�1|�ᎯLZ~���d��M�F�;�o�B߂/�K_ze��@$oe���˯�#+��-�-���?���Z�L��d�>��K�<>�x�0N��kL�7$�c�����?�ҝ�h�m�'����7T����/s���]�f^��´��c=�3�(��1ɴ�>��rS).�&Nԣ}N�]S����I�����C�[���.+}n�� �a[��Y���T��@|�m-My\���D���Q�$��-�y��i�A|���R�T����}x�*݈5#~xo�P��^��b�J��#��9�0�36���{�͜���r�ѯ�i�E1�\���r����,�PF	j�.��c~F@o�g�ɨ����-�M�bֻ��X{p�[�Z�$��
��qìyJ�}W�+�s	a�c�71a﬒KZRnp��V�yp�R��ʠ�\b�X&�Ac�B�}���#T/��J�v��J\�����n&���E�I`��(����k�D0l�1��>
�؉��?�Gn:l 4�C٫�ID���\�`��_W��K��}k���QP� �����e�V7�sy�*,�^i�Y_?+���F0raB]F�b՘0��ws�l���1��,X��-�-�G_dm]���=�L�3kȖ� O�Q=�]�_�|[-���JZ{�����!ne�U��x��y̆^]ͦ���5���`���]։���#\���G:	Ձ6�v�:|��N���y�����^�8�����!5���i��ׯO� ���VcȘ��>7�*ke��]�~U��M+ӿ��.� ��*Ã|Ӹ�t�kr����$eJ0�b6����-ǀm�nU�]���T�e2���D��>=d��L�QM�D�g<�l�	#�X������!��^4�M
�r����vJ��FGX8J��FÚ���?�Q��t��k|mޑ����tz4�}���S`,�@U�/l��5�#�HQal���D�2Ǳ�:lx��2�h�/���n�;�^^is�+�v���>�I<P�G}�D�Ě����t�����Z�Ԭm�J�����߾Т־��scM�����G���}lH713!I*m#�4_?WQ�%q���V��-IXW96qf���Ci�4�9v���k_�MF����%ߠ�|h�����5�\��M4e��`��'C�>VI�e$��x"'V�Xʙ\j"U���wʧS9�g.�Z_�'R4+C,:ƅN�A/���h/��C,"fի�G�u��'� 
w����s��o@Td��[�]Y巾�A�\�l�����}�C���փD�!�1R��p=�Aʠb�v�8�U;�`��%8^�~�NB��TGL���ԐR�E��F�C12çoKm����ˈ�U� -KB�j�������SJ��ZD
 ή���..��n^���l��
�#%J��)[n���S����|���cCΑVC���z�6\C:/�U�[ooE�E�Ąn����X��v��37��q��+K���3c�χ:�󘧿�(�@��|��SHY'�u'B�m,c"��wkO���i���\�	�\�6�?�	0Ή���%�)Lå<s_��@U�|��c�|���|��E�R��P�ۀ���`����q�Ą�7��z�Z�?E��`�M"��`d�Hh3a+�n9�7E���'c�xR	�=��1ԅ���n�?�%��ᧄ���[I+k}Gfr�'i]�V
��	��W�}���'�X��GE����
��q9q��d������1HPd��m&h �'�Ro3
ا�3߹a=� ���a���$`��|W���&0�PZR��Ԑ�
�5O�y���'qe0�
��}�[��=�/-��^Z$*�E��A{5�e�cYAE�W+�P^�6����ݯS[��Qn`�E�rf.	"<�4Υ�6����N�Z��t"�w���M�oġ"-���,vm�>q�c���/}�����C7�Yd�ý{!jn�z�'&G�>�(p�.]��I�B)V�c���ȶ���_�W�o �z7����r�M��&���V�eb���8ʭ�_@d7;@&Xy\�ݞ*�*Q��A��}����\WƩ��Rq�@P����N`�:�Z�7����|N��,1z�h[J��q��k}9-�o�;"*=s�0t�pƔ��벾J���N�/�{b�Xv�f�D��E=���(yQ������Kn��uE�]֍��Շ�i��Lۋ�RG�T���WD�V��	@�6>��S�F�bИ�z����(Y��Lu2,�b��-`��/mMyܧ8�h^٢�!�2BuO� 9p�O[ԻR �.�;Ᏻ&c�)����7���B�z���M���\�2�Ń.6�b^�\�R,7J�|�ExGY^{� �O�1{Yj
�m��>T��h���mU��p�` )��/�H#d&�ir���r�y��Fc,���b-�?�`�}e��hy��@��6� &���9,q��?�G"�Iش��2��='ی cypFdY�5�V�A��HZV����(�Ê����0҃@�+�&�y�Sw�SD�.���s�aL��)8���������nڂ�BY|��u��&�t�D�o� �.�c�d6$K�b�[�T[Md�@�G����KI5h����ێ�����Y���
�5�xj����f\�ء��Tό!���ˊWŰ�┒��w�!N��;~Gc�6�T��dn�+,6[�~�
)�k�*��Q�#�$��a@MN#��ɵ͙Q*�S��q+彔W�c!@�=\D^;�G��.��f��ɓ���n�GJ_W&�21�5,�r]4��dH� _���OE�(%V���W�/>K�T�q-n��� �z\�jNg�j�t��C�Y��i૵��D�Q`(mKD��cXz1������0>V*�M�
���>ǳa�A�ҥ������=Mh"Ml4��-�k�mk;��>����وl%L�z�_{!qtx
��U5��w���R&�������ϕ��)<�j����Sv<��g��ry9�g�E=[8������æ����` �A͐_�Ǵ�o�&5Ty��4���栖�4!v���A�����o���A���R��S�n�-J^W��g��\�GHnqѵ%��p�8�c୤�=�P���Qa��S!P�����<�@Hl��XlS���`p舨�{��;Y�Zi�:q���Zۊ$��nq�ժ��<��K��a�?6wr�y܋�+W��(3��z���;�d+���u��%�<��R��@�0[�	]u��nB	P������Y ��\:����px�+o��J�/s�EQclk���`��R�K#%���p1�c`���[�jF��A!�2�6~;��`��iQOa�\�R�m�X=�s����BmE���1�X�m�.�{�*۴`����*��Dҝ�L��e�.qP���7��St����1��N������^�%��.p�7ɂpY�q�?�n���kbu��ۓ��G�W!�v�0��Q��;hu��̈��:��fI�Q����J�Hxҕ.)�Jx$�E�lUOx�a�M��&���}�G"ŝ"�8"���Ku���e?3,�N��� "%su�1�W2�_\f0&�!�3FX����K�Ĩ��fY%�з�ٸ�)�ϐR]�Xs�vI�b�	Vw����}�)I�T�K���H�^�b-uo�f��E��+�<�!��D�j�c*e!TE����s83-v�g�����,b����(�cY,m��q^�-q�iTJA@�V%���?,h��HW�)��p�̂e�b��>u�G�~vڷ�'I
ً0E#y7�(LzH^KB��7�#&���q���gG�~]��Wb�˥�8+���<U�[���^FI`����jf݆����N��u������a�t;����S�y"��,�p���JNӯ�֖X�F�ԧ��M����(��*n+�Ʉ����X2�P"�*�:.���'�\{����ARER[b`
��A�D�g�`���(";~������K��"��3�.�h�9gAgE�`61�?%)PI�z��' ����1n��J��q&�@�M*XU4մT;o~/p�s�Bk�����t���&�c��调�������5
[c�"7O��fc��g�"m��@�B��E1rn���/�Zn(���'�U: ��h%��
wAF�fK��c�g��:A�57P6�t��e�=�,�	�@�o[�w�����Y���o�|��D��N����K�&��-��/~�n�@9��5���'*�,���?Wm�3��a g/�-"��
���f�	e�,[���8��4A?΄Q+�^!���p��|��ھ��\]�Zӥxe_.,U���	M�{l�p���M�L1� ������
h"a��'
����ܤ�õ$��:�z	�VA��a���|�ZR��n��4�:�I�4:Y9�R�6�ǭ���=lԘt�`΂GJ�vnĲL������}H&g'�0ӋI��AT�;7�G��ʩiƘPV������|�U����8�A���:�c��)j�s���;��
U{���
�1aK}$h˹	t�w�Vnԍ�uP����Óu����uW�W�Sj�/zQ��abY	�ه!�>W���8�Q������{|�2�Uک��9�����H�!��f	h�jJӇ,�O+�s\;���V���z]mT�*q��$�
�b�����8���Z�>=�Lu�����I�J�<���L@�uéݡF�i*ؠ�'�8IB��Za�.��(��m��0/F�9��#��O�m>+JjP�F�9u�������v%���8�]����"�B��� �͗ͿU�cL۫�	W�/l��&��؏��#NK�$��i.��C4��������lE��~�9�A;=w]:;`6���n��RV4`$q��Վ}֮���ƥK��}UC�O�nY�M]؈��~�G�!=�Kcz��h�7(���G�n���Jf�qBI@}8f��<�bK.��y�:�!��J��Z��ﵼ9u56�E