��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX���̓&P����6�O���iU�?jz�Gm�'�Y�Z�G���&���λ�]U5�x%�*���b�>��%1&^c���n�R����~�_�L	���Ǚ�k�a%E�������/���cT�1n#�$�"l��5H���$�]�g H�����.��*q%��Ԧ�]:�_���-M4z֕�q�5m�$�FK
FJEL�A���4v�JUJ�U]W�4@�;��v�n�"s��v-N��C!M�QO��Pr��"�w�K0�����E,݊+f}\*��Pa{%�K��g�v�싼#Q� [��R�R���w�����a��� !e�*eP�o���$�,�{8�YH��+T�u�kI�R����*'��,��[��q�=�$�F��w�o>QV���;G����>�3�{��zN��^%3ԫ�~ܿ��-�]}�OĻlYM͐+�
��)2���A���cxќ�\�nA��� y凸��e�<ț�<J�T=���Y90�b�-����4]��o!,臕<����) }�D��Ӣj﬩���^ښw|S�b�Z4>u�v��i��]��������Sجx|��u7I7v*%bT�^6���\���m�͕8�p`7����7%�q�f�X�f5j7�^�jf�s%�ge�0D�6,�޲�	P%�4���I��q���0jď[�F=!�hVS�,4�ӬL����4�n> �o`�L�h�$���^�[sM�,�aA��`��[���,���Co�K0��� ��#F���4�Lܲ&�����R���������,�F�u�<_����EQ���!2̋6�k�8�Il,�DID�D
 ����� *�a8�o9�v�~%����U�eB�j*�̜�&D~3����h�� ?G�	�� LN���\(�z�";NK#�mY�&�M�;�,�/�0m�v���TZ��#��/��/����]�v�!�v�Ts9s��>�oX���֠���vJٌc0�A}n�Z~�B:���A��#���2����6q�?F�-�1�W��i��I�#yI�w*�U��U� �b�4Ȱd��==�KU2�i�:��n7}�؊�����$�5��,X�+�+(�����GX�1?-,�+�>W����W;��\�KKh�k��l�G�ɥ:���	}�鄕�״+�"�V!���;�rY�c��Y��RKZ�6��GG�%���F�����a��t�/�<sT�NpV$nS�d���[{pOXȆ��p�'bɶT�M0z1͋�X����<�`s6�}�1N�����0$n���3��@gft�?0Z��'ǥ9���]������	٢6��vio��޿(�W���I	��)N�JB,0D���|���_jxtȭą�5�_�t���u��ӑ2�K��Lrڱk�s�Òi�e{�(M�`�u
���w�ΐ8GT݋��D�ސ5V�}@�����`X{��}����A)з�-;�n�mH'C
�Q�䑩�����7Z�����n�<5&/z/���1*Ȟ�7�,Aj��C�3إO�N9tS���c��T�Dc��a��BP�ރP��N�h#��ׯ �u]ut�Z,����7֣�zb��Ͽ�ӽ
���:+�2�=x¼���\9��R�;���1�����&C!�5:��DO�ޭ�!ä��&M��c���k� F/��U�gd1�[P���4H��˵��Cm�TM�W9�y��|/��/z���gbHt3p�C��NkH�Lg}�0�3�u3��;/�j\|��œ�2��|�_�J�I<�i>:k�b�.観�u(��A�|�q��Ѓ Y\��(��1�?����eL��W5U!1�4n�)*���d���}��u�k>��v0e�mtyLr��'��}	�E�����d��O���M3v�Buz@,·�iF(M4�iF���x)���/�e��1m�JW۟AM���Mkm`"�����Y�tb�,sd23�>�em2Kb��`�f��� ϥ��٧�Y�fW��"=��Rd:�C�����v���9���[�{^�Y2W�ɨ[f����9q�	������1� ����5���kō�>�1\��E�]�k�t<�9�ѵ��}!m�:�N�z�o���?v�z����]6ńjo�=Y��!�g�);��bW�Щ��X��p�hb7�1�G�2+co�Ӹ�D\PN=�X�(!UN��	�=�����r�v��(%�5��­�ָ��q`�{��|����ޙљ�/�D���Mz�蚹��x�r���Q��jr#X9�ɭ�8�1�����8�B{P~�9|+Ǆ�T�I�{ei��M��݁]���j�����Jp=T�D9 <'��T���c'BO܄��
����K�ǒ��c��WU^�6�@w�}���][u0�Ai�YޓD��%��W� bnl&�_�W�:����������<�wq˼�E��hV���@�Fb���$+_�#���L��_1r��<[/�v�l�TZ�U�f���cV%�I���N�1�L�?z�Q�"�����8}�S� =�{[M�[2��t��ԡ4es��u-ݧ���ulE�� �wA�K�@����i�L{kœq\�q�;��Y�8��u�}�����ɦ�����)�JR�/z����.O:�ZY�w�ܸ������3��Hן#�L���g�Ta�}�����wM����e�fi����1��8@Ph�H��-4C�`Gl/�E���"����A���J;�z�D�л�	��H�3t�s.��Q��2	X��4t���}kע\1�Ჹ.�ٯ^G�t�/���.�7��2�����US��%�D0�,���5=F�h��'"�L��Q��W�u�؉�k��랜hxu�_���;~'���Z��Lo;�oE)�91tb��
P��h�=Q% �����h�&΋���aJ�D�J������;~���RRB�O�\�q�B�����:�J���[d5���	�����	�,%��0�sV��Qܒ��|��[�k�^|?����kf��NG��Ťi�͖G��V!��S~����d�-`�l�����4�:�䗄�"
��܈������\��cf��w�Nr]h���1ஸ���ZF;�*�6u��>~prЁ�9"L�W���)�u!`4#S�����w��}�?�&~�)XǼ�>�=<�M���!�J+s�x�O�/�&��Z�KH<�V�S/�<�(�IVrP����yG]u��n�Գ��bpA��W��Vg>.��{�7� �V�1��ۖ���d1˸C�}�T)w�v>s�QuϢ!�zg8�C[D�yp��DZC�~c�R��+�!����\5�.����M�B��[5N�7��f��;�g·��g��+
��V��sq�fNc7��VN�޻Y�Օf��f)\CD�B@���5E�S0�m�=��SN���R����C���&]�g��C5�����%E��@\��׉$\U.Ǭ?�S]_����/��-�f��v�<�<Y���: ����~7lĠ�}���C�c�#4	���:3�S�̟b{�5袊��3>�p��p�����ė��/��|�P	
����E�{f8w�2��$����g&_�bԧ0{�Q�G�>�߆o�%Q��@���l3*L��!�&cA���=;�(�E�z��;�O�>��w3��<
y�yRk�Z�7�ƈUKl����[�Q��H�ȝj\MܤL��5��a�N������
�Yb��톌�rG�����-=+�ZH(
dU��z�3ZV�G����fy��#�8����	j��8%(�AЃ�5��P�kZ@ᮅ9��f%
iz��>�u��������Qg�2�P'QZ����p��Q��u��͡�|���
����8>�!��QIxJs��+cޢ��9���+no�j�V���g��:`UΔպC�z��L(��"n�#�k���yĶMZ�g�!�eԽ�!u����.��/�8����})�F�:'��-<X��Lq��[շ_w0�Wn�-ܶB� ��1�|�'bYK�k�t�d����
�="���|mzJ�9�<���N徰*�.��$��"��?Pϼ���_�"�Nl���YD��gJu�2b=8��Vl��ܻ����w��i�� 4z��*iذ�6MܖXC+��*���m;�W��;���@�{�"�DE�5�#=�T�ʿ�v8/�� �(0ĿAolـ�4���
ږ�v��1nn���[lQ�q�̥�'6���vW��N����;��TnC	ȋ���O1�}Vt	%�ue���0�}���ϖ��[n9}�Νh���+�V�������-W3�9��UwM=P�*Y���%��[���[����$�%��|;ȁ+a9\_���J��+���{)I�x�����YF��ѵ�t+��s�V��]����#��C���/]�/ ��Y��Q,�����&n+��S��7��Q�4&�A-��LDS?�iƔ�g�6�dO���r���ykE����gcb���!8�0�9�<?���W�ɀ(�}T���[�[?�(����`�7�U+�L����S�L#�O�
H���o�,�l�S��&���!�}��x픽��z��J�~��Jv���cM~PW�����%�2�5��[�H��`s7Ȯ�1��-�.���<Rx>��3f4�j��G�Y��v�QU���FH�3��#�C�bPS��*���Tp6l�N��Xf��Q���}c#|ڼ��-���'j@�~��I[o�?:�a�J�Lb����P�O��O+�	��"�J�����y��ʛ��C>١��{99�Z�s�Th,,�?�J�7��B�]%(���[�BbDjI�ҏ�2�:d���t�7�na1�SH;�fT_p�s�` ��%���p�����<s|�����<���EQ~�D�.�
�++,h�������41��������#K+���9J��R�g���{<O{���_��q�So���X�e4���q}�D���l��@"��U�(`2nn���O%ǩ3ڡ1;��1$$V��!�!�и�������PE�΢[)ղHW��P`��&R��H�-�gnn�R�{�$�����G�X�_C�"��۠�ǟ�x�}���y ¼@=J����
�BUH�`��v�`~nFu�țt[֝ݾP�U.�6m(s,%ZDF����B��e���R�����$NugO�	M�f��0>��x�\�e����.0�5�ѓ���BH��X�#�q��R�%O�'�MQk[�E���N �VQM���C/$��~�!I��)G�Q���,j��ߟ%�)���זX�&��m8V	p���&�s��T/�P �e�!T~N��~�`E[�����$���W��㞒C�ܭY��@���E�-2��#u( T�R�+Y�Y6�5T;*$u����梨���B�\
�;F��^��"���PJ,S5oV(���S��q��b����t��K�I��R���+�zU���!�O��6�!��_�+�!�\�T��-�x���ڀ P�w��l3\y,� ���#t�ѧP* �]�8\���z���95�#>�$3Iѝ���{�4X�Ճ�%��Hj���֜je���6����}kSqHj�M�M�`1]�#2f��HY����O`��[�V{�K�h��NƠgvB�%��
�`��Z�tݑgٿH���C��餫�>��z)� 3G��@^�{p���jp݉��}�]RQ*��S��u���h盼�Jm�Ͻ朑�| �A>J+]L�ZkխO���ιϝE������s������(��!�?g��CE��{�&8��P��� ���SE :�k��[��?M@����Y�S���+�Qg�j�K�^)z��A�e@��8�X1ΰȟ��o���i��7
!鶩XW%k�+s��b��
�5lL�{mV�L<C��BU���X�i|��=�6gXw���V W��&^
D�'�:�ģ��m��rf8{?f���Tɡ��Q���h,,��B�q��,3��������|Ϛf��B@`��К�fes��١�1(�q&�,ᖩD=�{FKZ��cK��01\A���T���P3���v�I�Ț��)l���������0ćw�(Ӆ���_���yt/W'�.��T���:]:<�(��8X��&��נTx���E�~�£V���jtq��0��A@�ml��\���ad���F�WK���V��w�`�^�f���!m���|�C���`���)��.���ߘvPw����@�ܺ%�[-��:e���FN��IU�7L��j��O��Xv�Tn֌�nzh�*��`��������K&m�����Jۓ�+�YW&�	g).�7�Z���G&P����)'��X�r�Ϧ0�ڻN�,�g�b���A)�z��Ma�j2:)T�(�~�%�4�q�fh�,�@��0��?iI�卐t�{(����:?�!ңe�H�0t�\���y]��	
�Z�k\!��{��"�-���!eGȬ��2���W�Z��^�����`V�@\�Tb��m�W��έ9iz��oe�X@ҷdJL�`�گ��y?���p������� :��AG=[�\�.�85��o���ç%��Hq�-�L2\Ո�� �QH\.�:�]���D����2"Qs���4u%?�\�Dc��y��C��qv %��>���5W���O�}`�N/ˏ�e�� Q����s��̀���WL9d���FN萱����{�K���W�]Xʄo��by:Ա$�a�_K����2k��]�[���s�vN<�'���~��I�u>�07�;�,dP��n��k�P�H*��=T&?�}�3��;]�z5�:'9a��'����	�B�7Ę�|e�7g�|y���t<���Ow�� �����Sng�C��� kL�װ?����\晤�;�Ll�`d�)�G4�!����i#�#zOg��S�K�#���Yk���2.1r�"�.�ܥ��Cfbx�C����]3	����V�0��@�j9��Ï�"�_������?i�f=��|.T���?��c�S�(1?�>������zUu+�P�.��6TI� �'T�[�����FXv�̼X5Tv?���fQ*)�������� ��Ւ� �Q>Ye��񓃊`�ꯗ�FS�0����3Y:R������� Qupq�G��(�v�8���y����ɘ�{��l`�1�;?�'6�Q-��u�HN�.y��	n�!W��y����ٛ�#"SzbR�C��-Ʒ�/+�+q� Žr�����߼�0�+����	g2]��kQ�Pv<�V���۰�5�j��	h�����c<*b)W��<�[���J��^N��������pU1��g-��� ��
��+%�-Kj�e��N�	��>f�2B*p��p�u�A�f���K���-t�CcU*�h((}1I����F�\GS���D�z�l����@HuHY_��ϝj�ěq�2���I��S����H�T��At�G㢶�2��7��
{4j,�tF���{��b��+�������1M"���@#���c�F��ק��=LT�!�6I&-6�U����~Ⱥ�H]��Jo�_�i�'f	}�sG��Db3�VI�F�v�����6'�ȭ�;�!^2�Wr���,��Fa�M��OG���B
�Ï���s�Mj	ǃ� �/ 7�M�v�O�+<��m3d��{�
83��(2�����P����Р��n�NN5T��[�NP���o}T���M^�Rˎu�9��S��|Ko����ó8���knv7�r��Q�´�K����Nu����!�X�	IX����z�n���z��`Y��w���n�k�v��U4	�ym�JP�4G;Ldd�M᧋��^_�Bu��(�����#2�`g�ht�:���ܧJ�.�Mfʫ�A�w�)�5M*݋9v%	*b��H���A3� B��\��>A&�]��h4��*Zh��YX�uY�X��	j�L���c�xb�K�\�V�L����Z�=��4�B�bi��SF��wpz
���=4-��:n�����v��I )v���"r����	�̟C�Ӓ�ܤYeѨ���$y$�C���Ϳ@r�E){�@�lD�
P�{0'O �7RG����p���Ә�4q���NX��[�!�>��uaM�5g��A�Zt`s��\9 �l.:jҩ�EK,Y�"ڍS]̰�a�~#��w��sN�uGz���fX��_鄵����ť	w���s��}���ɞ58{�p�զ�
�(<l{����z��V(\�a�(�Nn	��7|9���9a.Ғ��!�⎾�J9��ĆRƲ�G��0/��K5q�O~8��[�=���8�}C�Ӎ�K�D����_��s���!�R�Y�N�^Y���2.S�`5,L�֖�w�X���Æd�Ag��Մ}����/Y�u0V�+�
��LE�u�g�q\}��x��(���Yclu�!g��7�ǅ:�-�ź7��ׂ��>�s)�5�!�ۭ�U_R�9!h0��@F;`&�B���`m={>ma�0MFx��c�H��%Wvt#QVt� ��� )��M�'=������['�e�$=��=���\���1V"���ܓ���DsQ&�]#�ѹ�Jb�K�$quM�����S_�]Fw��<_�m/4 Ij/k�y!���hh�$U����:�EHR�M�1�������}�H��W��(Kwro���H������0��%�;L��0��R�Ə��k�ӗ"Q|�+�����9���"ѽ�}E�[���z%�'�ӡ�6|�72�m��<���*���O���1¨���<YE���F�K�K�Wjl6���H=� �<����Բ�e��P�B�_XъKA'G5�MS�]P?H�p��u���e�x�n��)�I��y3�x.W ����W0`t� �]���ߦ��F��.�v��C�|�$�Ŀ��� ��<�C����,� /����!lI�rb5o�g��.������2���� 3�A��<^����ǭ}�~%Xn��E����G��ft�xl�"ţ{�͔�q(A�y,��>�T��H�yhϧ,ģ0������Z�P �V��4Ώ�c�Iݛ �TNۑ9��Nfnbl��!��� ��SsH^r�����0<R�^-�t�nBEo2k���v�̕%���T��
��%D�P1lO#2�A�] \5G����8&��L���\�K��Xw�R�����p,�^bO�T4VN�kU��}�6�;��m���_��>��Ŕspx�����c������/����i6�����:,q0_D�A���Sd���*V��˧�qg�B�/��:�'_-!L&�M,Nwר���i��DpRE��3}$��j;��:�T��9�G�~N�u��KsN�f��#��⿓1��f��K\��?T6���[0��)bq���� Y�޽a��P�@'ͫ�E��Ǿ��,z%�x���*��28CgL��;t�� �?1�;!+��[��GQ2��o�-�q���.�M_��n��,���w�笍9��jA�)><,�0�����Ai��J�,q|��I�:�����<�����N�E�ozE �!
fLΌ��P$r3#A}�������z���oY4��Hm�"3}~cG�\�Ll��
O=�_��&���Pq����@\J�ٛ_�;�S;@�FL�k��]���;��C����K?�* ����q�2����U�Țr�ҙA����g|ӧA�ة6i�Q3CT�b�d����mcD �1�@�6sz���|-�b�[V ���:��y���a�d�8�4�#�4��p{�D��Ե51@e&��?�"���4_��XS���1����Rq(v-p�hV>S�-����P�ꨍ���\�rp�k���-����������0ԯ�.�L�K���V��X�����Ү���m�v�_,�̊���B�)�J|��kS����5��P��LRq��9v��Ì����=h���O,ˈҩ@@�{�K<���s�]������g����bm��&�L�y�'���~�q~:����y�"��ȫ�kbHH��4I���,���uU��Άh�3��;W�!JZ|F�~}�%��Ζg֪C��ș�H����Ҽ*�����Y��d��6�h��t��n���͚��1E� B2�U�q��7���^~(�_�A�x��_�ί���b/O��>���������Q#�Xꌨ� ��,�u,�@���ȓ�C6Z���u�Wl]��W���{���M�u�(�(�+h&;����8�=���KE&�HXLK��K@�uo�-N�Ӟ�N�Q�d�#<P�'�}��y����bTh�N2��a�L�#��X";�����0Ǆ�Ji*�Nsn�s�_��	���'�W~����48[�^�7�·����P?VI�! IMd�GVڐ��â͓��Z���� ���BT�KLM����dE��s6���{)g1� 6�*�/;�:n	���>��P�?�acȱm�I37Z�A�Zef¦�0�K�B:u���B8�!�ټ���>�T���2(�T��)����v��F�/�#տ�q�hP>�sl�j��L����� �5�Ŋ|��:���b$�̩�v�=�c��9A��vf��J.�E�S�M$���}w�az*���Prw��,�_ay߷��q9x~��Tŝ�*�J���8�ֹ!Zk�f�u�%o��Y�ܔ�F���}�~s�������Qh�3q�&uʄ�	�C� 6W�N�|M����5 ���6('�$g��">D�G?�3�ߐ;{nU�R�t`�,�Vm�'����Js�R�悘��֓�V��g����f��߯�V?��
&�R��|��+Vc����1�\��#/���֑g6�h")s床�&��0c��׶	�q�+�_JUF��ۖ�}$���t̵K�t��J�ף)zw�� ̦#K�_�	�Pc�6m
Җ�Va4�@~� ���P�Q��U%\Ťh�k���.��?��%���ѵ�Q3��Ū�9�Ɩ]����Q��W�<�L�]f��T�2�a����m�Q��ዀާ��ӵ9�T*g�9��S#�X�!�����?�m�k�@|����W�����>�yN�J�w��oC�����ΜDO$��w%�	��=��!�E�LP�kyq/Lս�р��puez�!�/J`�E��	�@�qj��wκ�fT'����5�c�o�� �~�FO�K�	x���!�h���JA2�7��Mh��:\���T��g-R�$z��}4ߧ�������)�U�Qo^�XK�v�>r3�ä?��PD���Q 1�L�e܍���a�zR����H�T�̀�r1�?�Q�_��.�ހ��^�2��6��s6�����
W����֚�8��=��A���B �]� �Nr�]]ض��,>UHg�M1�Ξ�I%�a����)~���,:���`�����6�/a,�D������>"M���ՊP��D����g���(B�ʆzAB��M��*es����������C5����R|������h_��J��E����"�!(�)I�T���Y����{�(R�1�{#T}�U�|�C,M�r��^y��j�z�>��+th�5�r�WQL��ݡ2��]F����'v,�W.�m���Rvǃ��nBv��y�m�`�0���L����	��e )�d<��w����!�":8F���@Ć�}����
�"���1e�0�ƾ�`t+u�S@_b�x�a��2�&z jT[
�-��l��x�7��h���w7�}F��+�"yқc��n��*0�6�JG�y?^iE!o7�J{�i���k��_�n�����X<�4��_��ޢ�@ǩ|�'#��m�y ʏ#��<&$L�LBs��6�@�w�v�(yq���
V
�s��=�=���Ö�K��R�o�����CFBª�F{JI�ߪs7+y��_���ؓ�/�R��:h8����h���i�x#if��o���7nk�ה'�uL�B��ft��*�0h��0����$�ǎ�Ȼ�{�[͓�xR�oN�D�|��� �lK����P-z$H�k��rۿ'�a��w��S}��vَKt93�y�VM��V5�U�)�)����$�Ӈ�9jV�ʕ3��7ni����UN��u����MN��g~q�С��U6;���n��Ԑ ���68Rދ�mn*k���cW[�ٹn�:��'N�	�2��������K�2rᎮ����Z�T0����}*�#���S��!T���/4��do�B��Ǹ���U���֍�s�'�pZ��m��* ��s�v�Ǹ!?�h���d�8wI�eOBلO��󡒔i�db]N;�~5���V�ŧ��3=<�M}Q%^1B�⡀	�D+�ʺ��U|�;1�l�Tqq��gY�G��'�i���Ejjg��(uR�gN�qB>T����^�.g�3:��'$~L��U>9�Nd�RR:�:�� ��K�(�����H#��W�Yޏ�y\Go�@�k��B��x}t��H bh4R�5���%�x��Z1:f����hc�0��[�%t�
B0=Z�x&�}�i�K�
Nfnl��hn�)4��ʹҮXثna�I��H�4�Y���n�f�j*օ�pi H��2�Ub��e"��/�&jK��ڢ��-����>�6�N��E ��*�Q���J�7I��Ìhb������T,���TtQAJ&�����7���a�J1��I���k@�����a:��&�4�y�6����;r��o��9��e�Y�����( 92F�r L���%%M+5�5NY��DA�+n�2k������C{jʴ@����3(�CPb�|���rz�_���RtO(��H��<���%�#9������!�x*�gv>�*��|[p4���M���(�����=L��n��4S��]�=��u0�߇T����3�F�Po��K�z�p���u�R�Hmb�jؠ�4=��f�DmdQ?j�|��7hRv�X�����@`��,��mg'�&o�hN�B�ky�"���/Vu�:&���,��_�.n�?�ȺR�KXҷ����: �o�rݐ���ؠ]�L�ݴ�^���U9`�3X�+��m��9����@�h�"�eU�+��7'y��̋�u�����H����#��C-r��xIΰ�V=D� 
���$א���,��]u[���׀G=�j�k��޽`oU�j�& �J ��|�sa�7�;�C��Xc��^�����U2�W�����U�#���\:��-1�=�ь���&�;~s%W��t��͉o��7���$��>J`%bI.�䓒��2u��� pc��1��̵��M���:���
����˽+�>�<Rb����<�I^KY9�R��qc-l4}�d>?�}(l�?��R(i�g=��]M;��g^��h�d-P��!W����	�_�|�v��=��Y�{����,//�;��?2`�B�(^ڼn%/�;�@��o]b�Z�.7Pu������)@�R�+&/���l�S/�� ���9��nV���tG���X ��!�"E�Wh�/Á��_�#w0�Ҥ�9۝ӹ��w�R����?~��G��?%�T��X�B�:����r����F�N����h��G!��_yCll.��t���7z6T�嶱�*�Y=���FL�fq;A�홝��
�H�w�A�s �$��2̉UIlY����.^�\4���~L�r{��u7~��w��>�]��&�����$۽��&5o)�,5D��K6��i�,y���Q�ؾ���7�@Iڟj�V;}'�if���o�B���_[��B��?��B��>芷�^��GtVОl<�7+P�3[���|'j�f���_c/j���Ma��� �7)���;�T7�fW�Ne���\�28���	�^U��Y����n�X]�n0�Y,�	�G쬬%R%�^@����O5��C+�9��
�t]�GGD�������B����SP5�\�������)�UB�$i
�#��T������L�u�H:p���4����ai�RA��'�������_��Z-��K�(��A�%Ec$[ʞq'���I�Z���3jkhdj�x�ſL��4��RGh�?���W �����j�FU����51�|����ygH�^%���2B4�#վ�8��,��B%�Y\�q>���6:��7�'t�����M~�{"}�LX�H��g�ܦZ&*��S[yg9�I�k�`�sF��*�x����³��i��i��Ȯ6#��x���>g�I G�#%V8�����r4���q�<��T]QV�W+�w�B�uv(�>�Y�Uӕ'{���*tneC|cy��.Gm�4x%C���@딙̴�,�w���Q!DgM���hr�Yl�Jn{��kqZd������6�ך!#<g7�4�ԯ��y:���A��k��2��P酺���+����n�h����ƞ<j��[񉼏���B�����~1�V�)T�R�ӑ��Q
Dby�\�kbc	�.�c�#3��|K?G^ﶘs�A^���w�t���&+uM�H��W��oB<���A����邾�ԅ��ey"��2���ԋ����O����N�z(�
�P���boC�N�oS[��t
9Ŏt2v�M��ň�v�kA�e��T�J�'e��Qs̝*Dм��{��O�!s�ؒ������#�?�[9�x�!�Fnǰ���?����1��O�\x��q{�	�Vhn��*�bD)���WK.5��b5�nv9�L&S$�0�F�/0��4�Ò%��hF�2~����rN��	e�$�F�ZAfG�䆚�^nJ�� �2�
����QO���^�e��˖�O\�7�
��`��xY3��p�"�'Cn�#}�G3���J��~��� �ܮL�=Tv�/t������:x��*����¤h"���)�`���&�t���XW�ķ���P��rqTU�z#AC�oRH�ʈDwK���biZ��c�戒�,��ڜ����g��K��*	=�ޅe�l/`���~��F��ӱ���A`���o�@�� � �r�Za�x�W_CF}^Z�ɱ���4��b�����w;��}�2��eת��f¸��D�g�-Sœ��]c���/5JI1����y1M����������~7:�r����H 7��(���r-mngӷ9�f=��2�����Xt5���M�ʅE��_C�hh�T�����iR�w���
6�ɰ_PDEg�8�ͨ)zGmF|q�={�z�IS��S��!��"��8]�"�č����	��+O|���h��֋�ӈ���֕������T#������ ���*֚]*�ɒr���C=�2���A\~;w���Wf@`����`}�=NR��e4/��m�������, ��OC_��f����󥠙�9ͷ,f�irx�c�K����:�^��}�bM�~}Z�2nJ����[��ޓrc�b��D-�jv����U�۰������t��92�y���)�����^�̤� ��5ZLxC� ��Nһ���Cj���R@�����}���|��&ԜcR��!45�Z�^\��*59�)pR�t� ���������A��Є�c"i�dM
\A']O��5ә6eo��XF%^Sq�
s�!+��X��n'	��6�0~���4h'8������n���77v�9tˤ���,�M~z�����r�����ĺ�4�����U2~1?����ǁ���+&�J�O�5W�1-��	㙳`���q�Ts�I�HaǨy�9Y�����l:��Ix���h���͘p���=b�Ģ0��Q�+9Ȋ�E�|.�XC�g���2;1���X�@W��mg�#t��%Ej�T�_m�5����*�B�F�~�?"f�>���k�aU빲��a���䢷|��;�$�r��,��#*vS@uV~� �a|H��4Y�� ��ت���Wl�VCx,׮>��8P����-'9���2A��	<������d�g<{��l�D�
W+�poU�b�쇝���`�"��Qv�.�!-4��ه^��W�|*���Aߖ�^��M�_��EnH����e����4�����[^��xlP�H�HC,?��P��a��}�
P�2S�~��Uz�|�PmL0m\�3SE�ޅ���@W��'��*\E�)w�]�(.,o��K1�UR�������E�C�ux�5qK�8/�-����z�l����r�#¸|�J�9�xH�{%�#�u�m�do�~�-�7��iq�P]1�O�n�
�[0��%� h|:�
>�c�Ӳ�3Q34�����#�1�9JlЊJ��2Tޛi	��ˣ �x��x�/�IY�^��b��#�k���Wb�Yͽ��������E#:��ֿ�O���+9��x�L�+WR?P�$0�(z�_V�0�Y�/��b����������9�=�#D4l#��/�e��N[	d�Y�*Uנ�~} U�X���F��f���/Zk.*%����ո���%��g���UUˌ�,��t��B����S�F}L���+;H�
��]Q��U5�'��� �4�j�Z���,�>�uy�.SxTD��~��I��V��搵����}f�p(e��4h]4��+���OP���M���0� �_{M#4���h3`��g��a���Oo��;B�ND��jd�Ƥk T�Mr֘�L)�U�'iMSzJ���a�2Y�Ɛ}���c����2嬏so��Ț�Ȧڊ>�ZJ5EY���3��L�nbzkfP*�oH��.?�ߠ*�3���43�R�:��f�:���7 #.L�k���o�hT��LA���M�h���#�S�b!����Qx��c���m֍Ѐ�SJ�ٹϖY�>_[�!�h
Q��"!6F״�I��.�*NA����S��Fn�����&��$�8�	+4�*��`��l�]bhQV}�j'���uh��ĉ��{a�h�wr�OGi�U�]�T��U^o�I�� `�ӆ��`Rn�m��/�V���
-�ꆓ�a�"���I+��G��jf�VB���z�^�DgZ�}Q���A@�y��kR�a�;0��!���@~}8.}H�r|���s[j����$�ڕ������$~�'��(k����5��z�"d���ߗ���L���uŁ>�Z���H hK����Ø��{8]���y���y�Y�Z��H:
׶z��i��i�I!�˧Tg}:e��r�!�?
���Q�ꄷ�*I`!,��FT-�᪬��S5��Y�ě�������(ʭ%�^�ӣ7bEBy�w��sn�#T%�zj�h �(0G\-�VP#�	4�+�U���$]��ĮUF�o�^����}�'0�cCL���e��;�W �B���`'�h[nv�
�O���¹�zS�������X��Z�I�<��=������i�QoE�#�=֐!n���`O�%x-�οE�W{U��?�$������~T��M��P�O�*+]��Ztu�(;7��!����JL��h���Z��Cr����O,�.�AI�F�ׇ�>�R������N-2>8J��>��i�y2���w�_o2��.`=\WJ�m��}p�u����vI4���H��4%Lوq������QD3!��AşhM9S l�;�M(Q܁9Ыzd腱�F�Q����{Ct䒘�x�7�ې��}j����E'Qu�9�t�T�ˈ^(�Q�P�B�%Te#�~o�lQU�;&D7�)Yp��T�M��<۰��{n�ި-�֩BZ�5�!� c},��p�5�
 ���� \>�.�M��(]Ly�x�,I`�Ƿ���b�����jfk�;�nS1]��
ĿA'�?��8�Q��%� 1A�^"w^��s�#۫wOFM�,�v������d}$#�WLE��$�\"�� �����H������r����OC>���ĉ��I;YH�%����7�9a(���u��I��ӚH K�y&�Η�?�+Y��[��?�Q��O)9�w�k�gi�Y�qg[��SYhƅr�j�{D�����\�G&O-�t����p�c�S�WT�3� �y�=��a^a�	�)a�$� ��t�&��P����]a����ƺ�ƭ��W�Qݙ& �1(-z�u�QW��Ϩ���V�0������/-�"�z�(��OL��!g'V2���>�O�H��RR2�I�)ƭ{v����a�CS��N����l�!�����5K����l̶����;���Yf�մ�63�(@^ɽV���ko��^Ǐ�]��Ե����}���	�t�a ���.�唤:��j6`]��� Ǚ����	,V����>����fw�`@y+��ڙd2�ܞ8k#�b|�H�W�d��%��ڠ�D{�hO����L2rն=z�rC�9�j��*^�~ަa�0Qfk̐L�bh�XW�������/�u:[�l��^sJ������7 	�Zn+H���C� �7mWo}ә��g�q:= q���L�k��S�ں�����.%!#8��< n0`<�0�x2'j�?�7�j8!��������Q�8������貮�GVx�{��3pc�U&�d�σ����b�da�-1ć�D�qO�6�	�(�<�N+AP�1���x�ud�%���Xm�0fC[^��v�4j���c��r��_�e�[f.#3�4���D���k��`8�� ��i>w�Y�s�yEx^�x�Nv�u�a�Z�%��i�������������1�phO��{h����#yKJ��T�m��.ZM�i&&�u�����Z���;]�d���e�Y	[T�D�O�b��gT�8e�#ӯ)ձ������5� "sX�h;���s�'��Ά�mAp����8y��.���J�ݩ�8�?�rQ2�E��ܣ�b`޷|&��Q�ڡ��^b��~l�:{
|ӻ;#��-T���v��U����Tp�{�0���Kc �������.�퀠�A�S�"S�O�(����S�J�8��ɣG���qXp���$-X7�>�`x�b�po�-}]^�jW�C�:�V����o�T.�Z�	ei��[ �{aj����?�$k��:u1�7����v���L��v&$c[~�?�Y�&��7����-�'�;٘� r%i�g�n��ߌW���m�<O;�P��c9�zA��y��2WH��a�qEs�-�����aD< |�z�V�{�ܸ^�2����B���r���([�rQE����jW��-���Ђ"��p��*���U�`K���n04ʉ�������?�D ��vHl˹��-�V�^���U�2r���-t��ݳ��_�m9��ĪBxk]� Ӊ��ξ%iB��>�'��^r�gh�32�1(�DF�L�f�������|@����-	5�GH@O�������r�����i.�BCܑ�)[8�~cc��؀�G�̲Cb2���M?h�J�&�Z���"w@c�=�j�� �:휴ޗ����OCM1�P83q�L&��>��t S����:x�j<�����UM��"���"�T�;��u�«��@9K���)�@���=l���8唭i�vUBIn
 W9��Jv��b.W�R�����Q��A'3[~�.�c�̢*8S������2�B���(�J�v��=D��ᯙ
q�X�{�{���(�cL�}v ��p�e�o0u�G��=]�۩[$�aꛜ������x�K@��ߪ/�q�*9c��dTY���s��3)`R��I?��,VS�&�fh�sDx����Wܒc^e��QȔG|�D��p�vAe�NaY���W_~���B�/s�,�G��(�X��>�Y '�;<3�L�n�Ds^*����G�x�a�[��n�a��B��*>ZD��d�X�HĞ|(��������k���`�vH;��9>��.;buh\O[��+�A�����Y��Hϫ���{=�ŵ�V����������瀤�j���
`��8!��/��~_|S߈L��@W��XN�s-x;���h�?qu$
�&XC>l��Tb�T�m��:�͜���[z�-��є�Ћ�b�1-�h}�PilM~HޙQ�)a-��A����F��=��W����4��Wp,�-)�Ƥ��Ҟ_*�\���GD�|HRz�!��a8:�MP�'k�U����G�"���޽{�k��CE�&���k���6?-D�c���*&ظކ�o�ic
�(�T���7�a�c�3��G:7"^���0�m�XF~IR롫�J�,�*zj��٣yG9#_:>�1��Q����GI[�Tm[W�����AV��TvPEZ|Ƴ�г�]?+����9�)ô�`3�JFс�]/v��R�j�A�SU��f�h�_�r�oŔs}_4�u� ��d�	ބ���V�(L��mQT�UV|����ZP��%�Ƨ�s�l�� �̀�0q5#�B#�m�iUc$�|�ܭ�D��5'	Q�uǢh���T-dv+$�y�w\���b朶ڪ
��9�[����h�S.$z�����/�SO.�D�x��Pml���?$M���}���;S����7%�ؗc�C�kJV�����UL�c��F�_l,j�������ݺѣ�@��d9�]�{$������}����V2 /���&�*Q���0�74)�5Ǳ�-�񠤾� t{4��V�;�8��&���=�uUq��+1��_Z�ˁ�p�h;h�~�dl��n��շ �T��7��a?�x]U3���b2���f8�U�G�p��ϟ��ump�ol��) e�ܩ�3"V�p�e�eg�E �T���s�>=ga=�h�z1��+"�4���l����ZO�Z����媷br)� ���i�`UY4=O�>�Jb����K��7�G����Rw�x�I��i��~Rs>(�b��K^Q�WL���9������� �_��i0q�*�5�a�l�?�V��n����V��i�1��ϥ�%�d.�Uq�5���4��9����>{���
���Й�
���c��ڇ��Lv���HZ/��x��:w���u:o��'.�וSq�_��>�m)�-WC�1q�ۖ�:y|�)���T�s�	<A]l$$�-�o��Ҳ��1�T�)��x�Q��POH���������
#I�24"��գ��A��$��A��Q�7�[V������t�� Ϋv?���3��R�ȷA;��qUz�e��>���z;�PC+Z�[�(Gp&�6���q;�qJ���!-<�h��^��X�4ʍc�k몡�P�uM{���b!M����-Ұ��p����Τ���TPZ4s=�~��>b�:FZ����D�~S$ޫ�Ʌ��'����_�Jc���Mx�����_M���8�{.��+�Q����3���]x`O��A9��;�����X��Kk��"���4W�X�|�����+�Ր(K�e25j�+Yk�W�DD`K�J����Q~-hN��ӇVɦ�����ȗ��Չ���'1��f�([N�"6��\%��"�\��5I��m*k�s#�o��)l�� ��b+���(�l� ���ww��eځ8��``�y͒�im�d�|R�7�+���:c!�a(�4�ﳀ���������w{��,�I���E|��F�����Q���r��@Bae�c(ftv���uޏ��A��߬��gE�p�1٦��C)<-������#���4��T�Vr���.o-d�r���p�\mZ0}�z���]j���ѕ�C%+�>����	��z,��i!�	Ǭ�,s\�h�x��ju��.�{R�l�Ek��!�ri���Oij��C����g�|�'��,���G�fH��"�3]�avQ�lS}X4�����*ѻLol�#�T<� )��c��σ�������0���k^,es�˫��Y �&�uOM	�O��X��֕0SAt4k]w�C���2aJ9#8⑾P�b�K$I:�۴��q3��Ȯ-�:���}�n(3@5e���.�D���1����I�Mӝ.(i��������E�b���B�h�{N��ɺ�a��Xy����E�<bR:�; ����#�@�&�d;D��ar��
V���?�.S�n;�?�ղ�^UdA��l����\`;���=�㞾8��T{�`�$���Hy��Z6	Vr�W����^Ў�PN��� �a�ºGY� ��#=0P¡_�ED�w�Ө��ƜAs���@WJZf_Rf���@_y��aα�N�<���ٶ����(�ᇦ�L$���l����?#7�g$�� �~�uO��u�.ƣ��_��it�v�^^G
����=��pj�g������S��B���;)����WIFNB��{N��]���(���M^u?��|?����b�f�Ai ��|���EZ%��.��QA3O��j;�>'���*$�}x�q���7ID�MGH����s�U4�m*�� �T�f�G�L'���n�@x���i/U�i*#�L~�4C�G_��l�ՙg@~j�ے ^��ҭ�h�gӨ���za���=��2�UW�!^:����_�9��WtLa�Z{�S@6!k�7v�c�E'��&�]+�!�9q�5Y�g��ֶ,�MJ��b�[ݓ�F�'Y�B�����c.s�1��l���J�y-l�B��m�`�! ��gS��L)�X����
{P3١��B1�c<�]m�i���H�9D�R$�r��c㶲XPr7��80Y>T�8~��r���lQ��h�b��BW��x|j��Z�٨� �V9��w�<Ķ�k��h��e�X�8%�X����v�ڲ>zs��&��iFc^�̖��6/.[��������L�@)\)��,h��
%��
�Lf��[&��g�g�-�ׇ��K�	7�JWfS\��(��*�<e��G�_��/#�));���BG�Ʊ��*7���3�8�\��T�ӆ�_�R�/�U�����������D�y	�׸�'��(��s�;�;�^;/*�j�0��=�$%W����Z
I2��&�Rl���BU� ԓ#X�̺�C�+n��s�=�����p6��9����3*h͖�^ֽ.H�Zi?H�i�y?�d^�3ƅ!sC(n+�i7{&��;摸�F�U8
N�*j�rtc>���8�V!	.��%e0	-�EM��ab�!���TT��1�y�Y#ި���`btK�K�W�d흆�� #1�����)~�h�&����D���)lXF7V, �5����:m4�jVE�J�E'L<���'~
$��>����yP��/���M��N=��Tm�T��e,��L3Ŀ.1>�S����n�}���<s��k��g���ڬ^����7)����'á���m���`�_b1ǰ�� 
e�
z��$�X��1,_.I>P��G��$95BU3�R[紧��	����-�?�WkV����Qky�*� '��\�n)%�x\_LϬ��E���GD����W(�_"EbY}�T��k+p��D�l�@�I��!W�u#�(�UO�h�O�����4w���_�ILf���]�N�-�����6���o�j,Bw�&R���`�������g7g��b�%��Z�曈*���V_�0��y��g������=���@���a��\�f��� �4���~�ae�������81�$=�b^��k!\���U���>����ۜF�)͌�cr��\CE���-�J��W�2�`w�ܳ�b��E]��0d�Ae�p�Q�M�WJi1~k#���U�����I�/,�#V;fU3��ʫ����caۖc��
-g}��΍U[�����H[��kn�m20QQ�0�Q�<�{�����	��-���C*�5�aDgFh�L�;d`!�:�Z��S�;�����ͨ�_��e(�b�\��e�帒��O��?��X���l7���CN
"�{8"J�!�����U�]^����%#]V8n7�|��|fNC������>0;4?+�-�F�S|LYU�NPD=�.��G���IC�F2�Nä�G����SQ��0ze2��$��}����ˊ���>����a���8��ԼO(Z{�"
���V�aY���� ݘ�8 �Y)�t%ӧ��5��4┎�P��%�^@��2[����ͻy��3�￷M�� �IH�=b��g^���g��L�h9�6��C�[�V��f�+"���_Ŋ �D�M&'+�p�+`D��N7�y�&D��E�+Ӓ�H��	ҡ,��p��^LI,� ����yObz7��N@���@���n����z�dw�h�Dr�ؚ��|��͢�l���*�@���t10%R-[��T"߄�2�$�\E�O��般7M�}M�&e2r񗁒�bv�R�)�0�5���`]�n�e*���|�4�����휠�Q��*�	��ͻfE�T�!T���C��Ϋ�L�b���J�^$9������ۗN�1,��)������wȱ��eU%rM�O?��6�ߍ1l-�K��<B%�D�^�aZ^�_�"B�ސ��)�8 )��YJ���Y��	r��bP�ӯ�����_�S��"?��?�l����yujP�j��%�M�4V�#6��T����tD� 4��l3������eɑްX�� =�\樺�ul��D|����땉dN��$H-,�`�m�J�����"�q6�Q�Ԇ��Mk��\a�"���ސ��/��k�FY�9�
d���blh��y2��Y�$w����$dl|�p6�	�h��?�Ȥ�\`�V?�
ŵl��-�_�g$r-["���n�����UC{ck�Cs=�M��er�y��<����Я�DY�����E]|�e��ޚ����~�=��`ق�/��A�}�c3�He�pi��b�2�eH!_�q��B�!�0�,��ץ��_�<�@���ל��z�&l�KR\��x�N�ʮ�b�\�MP;%��祿�vAP�dM��5��j��岘����>E��FZ�D�G}Ҡ��O(�q�:P|�<�����[�c�Ei0�>�Z����j��K�)c�ST
�aa)L��M�����W��rKk�&^|y� �#!�z=��i����'����K*6FV�{.h��4�385`�|�[�V�����:�=K'���A�e�
�vO�v����2�r�^�# 1t�4��D�?�Ds��6��N�T�04E��+�O��f.�������+�[f����7	S3��n���>k�dw��KOxF��^`����)��±�M/֤��y��	� �s
@����kb�)�W1���8{����59�{����7Z������̨�4�)��o�s$�����*G��C\�l�̈�	��n��CE�ht+���H�F����{Ev�%�t��@���He�� |4�S��29��c狰f�~���Z�:����)�t�2vb��ꤐ-q�/Ƌm�]��Lwz�����0vV�mt�HJs%Y��P�n�c��=�<����/�kuX�٣#�n���a��;��쯩�M�A(!5��|2NOUo�HE������;�w-��ϔ���Z;�%�G��ڟ
��ՎIIN���������vo��<_�
�:��kB�,R�F?���r4��$o���+�y���Тw���z���n��� ���T���R!���~g��MC���b>Qު���`��؃�b��P�p��p�5Z�ŞB��J���^1�Z��8D���-�,�����T�A|�@�Bk��uՑ�A�����Ey�?N~*�W/\Ud��
i�<�B�Lk�_��57�&\>�	�"t�5LNc��i<q�Jò���{JK&i����6+�A���u/�-JL4<�PD�@�B��u���Q�E����fj�,�'���qT����/]�giE���
�°g���*�/�*=���mb~���ͤ��ӪHWUƼ��Bҩ�#�1��Su�w�dT�ϡ�鞪?�|�:(L�W?�Q��&`��?׏TO�/����^�"��q���%'���J�8��nJWf��=�JC|d�.�b�� �����V�-��rh;�:��/�)(q��$�)u���w	YzR�U:Θ������-�~�^j#I%4�<&��~�&����ՠ��>�1�o�i�5<�h��9S'�J���MM8��	�S�����5�ͼ{ˤ���G@��XEGh<@h��9�kH���[%Fh������1㏆��������{��?����@�X�S�oW�C����6�G飐�u+:DIR;;%I%;nV�&�)�.�s�c7�B[��|�3��P�������]"��7��/�.Y�_��=�[v���
c���p�Y������d�1@̩p���9�M��(W!I�<��?�CZ��K0�rT�dv� �G^���'�����>�3���#wfq��O�*�Eho�]��d��rH0�Ԋ�"* ��qh���S��$Q���Sઊ5��"�X0�֢�3xǱ�S�t`���彜d��ԑT3�95Xַ]BP�V���r?�F H�[�ۄ4�hh����Mob���Q�l�Doz�ô&���h+���88�7
�?Ṕ�]� �qk#��ȃ 9�L/��m_O����\��G��	��	��m�!��'�3�r7Z��z����U�=����ߍz\�/FgĐ�MdM���f����0���7���b+���@q��m���鐾X�2�W�����΂&(u~!=~o�`R7�K~��iX�Sۙ�p� ��MLd�f��n
���W���i8��;s�9���^`�3-�z֎�s���ۆ���a�UPGu���PH�\k��đoP��e��}��j�7?g/.�!�;� �t4O�- l�E*
�8;Q(�� !纒��&�4�M"�;����3g�O� ���@4�pq�7�E��5�r�@��|Exe�%�ZD�b�e�?��!�o@���9�*��h'�MI��� ]�ΚY��o� H�Ta��2:��%[iI��&[=�V!gz�u�Z�$�5K���e;׏o+Z��� D�wj����3�
�,��}�h�+:������Y0��~�`�;�@<ԴR֟&_�G�>1�N:"�y�]���<mG.����?l=ڊhx&��:r�_�'T�u�/1>x�c&���P���n^(�G ��n7���h�4�4�W;�ۏ{����g����o��9zGۏ��ImpEu)k4�k��ۚ\�qQ�����ѫXc�3/C��V�;j�ӵ���e1_GWTH�~<��l�����#L��ݱ�	A���2�=�>�u�'�ȟ���9�)yt��tbYT�4�����r��ʘ�k����qV��J�{��V��u�A�8Ю�M����DK����Yt���F.�Y)�Ȅ0a?���w'3V��d�����|��M��.CDr�̽_4� ħsE����td��j)�Et����ֹ	3a�?�ߗ�>��sta�+D�3�D��uj/Y�I.��#�|!��}��Cİ��MH��X �n�t�}.|�tا�k�ǆ�����P���|�H
���}���:?�dh��j۰��5g�(��u��5~A<�9�.�s�ǂ�S��!��g�V�`�����,ZW��(3֜��ǩ���J�)�Z�J�=����r�rPK"�%����Z\���?y����Pq�{��\p����KH0Ј_tY�(.������ D��TTINqG��"p��B�E?����s��nvt45�
����d`�ٸ⋲��W4�B��x�~FŃ�y��msv)W�����N�6�{��џ_�-�6��&��&�n�2\ͦ��F�~�}�� � ƅ��ј�;ڭThnk��l.&{�
����6Mk'H�x���6L����4��e\�f��Mnz8،�u�\Y���xZ��݉Κ����yۆxG����ְrY�������������%��gv�PҮ=�rq�{���^}��z�t�G`�U����.�����,��%‮/&C/�$IC)����"��F���?��A3�Oi)y2������|r̘��M���(x���SS>��Bk}j��IN�w�a˒*{��R�Y�>�hMV"v�nI,�6����J&�2�d����ml�E>���Jn�;�+��qKv�I�-�x�s	�oo���3Mh�����Ė���OCR޷� �|F���0��Q䩱��y"h�n6|~�f�)�E�Wc�g��+���&����6�rm:Ctb�����<�Y��`�We�g�J����!��
��ȇG�q���kǫ}�į��VX�r�j��*4������1���\�H}8֋�̪'qi�m��yT��F�vl�s��,�XK�������[bY��m ��~JH>��m����3a�-
|J���J��6�j$+�_�e/���q�]$kӴ�V�9�X�mG���*.Ў���X�Dz^ ��rx�&�d�<K�+�/љ�{��*��}���H6��;�{3��YG�$0�,�ӳ�����ɀ{7�"L:h��E��B�%�u�V׬��[.���q��X�}�3k�މQ9��^*�Vl`	�����)���*ND��q�G�.�q�'!B}�	�o��JӿL��DK�M�mFfu���:���_�[�J��O��a�����A5^>����ܡ�H��j��0:ZŬPr�mi�\�D◇TM1���g%��
g���펋cs�����"yhP�B��z�>�[L��*;T���b=ћ�W��d�pY���{0n1���f�¿�"�:�0�7�(��$��5V �?�XT�
���sJ"x~��u�F�G$T�g1ҩ~� :�xڸ2&IXdr��ZGu4�$;�^�h:{�[��V-�+�m�؇�u�S��n�-+�*Q����N�y���\	Z�bj$�����Fw�R_����"��d�6{?!�i�h1}A�ج2���.�䯕�ˮ�����9�A��	֑�r���l�& *��Q��\���u����ߡ�GO���
�X4���"�$�I�����O�j[�@�@���W2����\��៸�*��Da�D/>y��^*�^y@�l��5����g�_S1I�tӃx���<��Z�����0�T�H��L��$�r���u��Z���䧭�Rw�LBt�2��'�Ȕ�v�vOu�SA,B ���6��n�h��㮪�����d�uMJ\
��$B�kv�kDwN�]v/f�q�߅���.���h����tQ��"��9��W�r�FH���c}�k��a'zi �j�"���"����D��HΖ�"j5o0��a:qv�1�kj��ڣji���QsQX��L"ur��4�t�;���nGOFl�y�`�ST��S-vx�7��Pl�|a�TPۑ�����q�;��;	<t熋�r/����-�z>�a��IH{KM�ѫ�]v5[)�W����t`��'���	��]h9��hY_�W.	/�ҋK���D�1�!m�7B�N�/.�j~ ��lu���f���j5o=�c��q�[�ypP��Zj}���k����ckY"w�#]�_^��)y+rw��F����GCMZ+g��Xo�h�zG�hƺ��6?��'��)=RM�&Γ4�����/�s��x�4=/�LQ�mN>�³�ff��F�t2;r�̾$e���
���g�,���ؔ5J��Y��c��-��J�/hl�^��r����א��<�8*����Ϟ�Y'.�g��+��N��"�i�ٚ��f�n�BO^�k-"�%zI@B�ի�W�g�����c��b9�7��y�6n�:�/m_/o;�Ui;�c�{�5c�)�|{O٠��ɃIH@�$�|Pr���Տf��<rz B0ʟ�m�v(�a�+/S��c��4�U/e"c�d�_��V�{���nn.�Dt�?�.s��@�&-�Dw��AEu��鞋���=�c�^ϴ �["gc[}�EaI�禉wKo:�_^k�5���;���T��vw����r�
%�3����3��NZ�L�8�kU1��9�̚g����B6��
�#��Ά��э����5j/����x�[�Ȝ�����b��P�����MXM����B�]��v����Kb�+��z�H?��+b/�{S�ѽ��/�M6�
7h���2�[`�|����i�w�Ӄ�C�rI�.t��tY�L�,����Ès�i=�b�H*\��Z��/��v�O���IgU��W�Uw_��A��C�|"��%���TԴ���й��!P/�s�F�c���mX+��9�f�TČ���f�&��{��'�A����'����嬍FE�ŌT	��>�_h� '��Q�p�$E��r�"�u��3�;;o��f����mMw�����)v�_�O��Ly$�}�J��[���{Ξ���%�JM :���n�l����\�J�y�=���Lsu ���oG�uxS^}�h�9���ʔ7/�
�MJ���Ҩ�ʩ�>6�Ԥ�"���s��ٳ� �4�Ėni1��	ш95��v
C��}�\7L�ҏ�+Bh�K�n�����ز�61nH��p���S;��7h��Ӝ�h�\��|�O�f�s5�j.�Ы�B�&��j�4���0�̿BE)���qdMnD�-Ga��9�Yn6b����> 9�*�1A�A��s��uC�S&سQ��D�	��P��KТD\�6��щ��r�Qơ�l�W�8r�X!�.B�	�٘VE�dE|B/UH*�t���"r^@$M��u��5_e���4Q�W�p��<�,47�h���L�ȭ3�J�@\΢~	N/����Q9K�Pu8�������	�}E��Yt7��+t�A�h��u>ޓz5�!���U�S?������TO�뤣9P!��n�D�DnM�
��@H$LB/ΤIFс��j�.8AR�Z�B1z�n��6OY�u�dl�����=�t��oe�нN���ƫp�d!�J��bP_�?�
zzk30�_�|U���Q�����!�E �n����W[��0�S3�,,��0��648�`��&���c�zC����������H�v>?�{����J�N#Mqi����b��V@��Q+�#Z�䨧�s�ѿ`��|D"�S�'�87��&����`�L�1�G�5 �����G뱣TDԟ�tD��Bo��BU@O�d̅{H�lc��o�d�\��	�Q$m�d��g)��)~��bQ,0ؔ�D��[�q8d�������+�\��/	N�P��ΟJ�������1 �ѫ�1�㬘*9���c#:�b�@	�`����:L��
��[�"#�:���>�4�p��;VJ��鮟�6-��� ���w�m8���P�����A��Kh8>I����r� S+�;o�3��G���I�+Y�۾�H8(�~�!����
��#ʠEy}-bK3]�:
͵��tЕ�<i9�q4�/���$UB8wxO	���Wۃ�&�C�פ��s�S�Jű&�Vu��C�D�غ1���6x�L�_.��|��C=���7\���d�����E.�e5�:�r�SF&�J�.}��ϓ���\�6bn�j=�{�Yah@2�X��nEao�`Ԝ��|���w[u�.���Ip�bʳ^E�}�����\�;I�&�nF�˭A�Y�:�e��ۇ^�zl�u�C�/�H_N���~�A%/օ-N�\�mĐ�9��s�*�r� E�|��C�{8�����*���
���5�/��:�k��A����	���@]ASH;���Wtv�j�⥈�@q�,a�-e5Td�ӏ���-��Ժ,xU���p,�G�)����\�����rW^�9�*
��w�.�gf<�_o�T����֑���A^7�$���H.��N˞��,+�
@l�n�V�6L�@�
ܬ/Ǳ�4���>Ӫg�ʹ�k��=|�+:eqJ�0�&yV�~T~�k-�=-'C���h�~4ʈ�c򧚪�7&��wb8x�x@��cK����1A�_&�S�>sN�\6��Bĭ�%��cFX�`%�>����K���5e��A˟��O!��[\�����$����q��;.��`>�Wa2���x�����@<$�>��ms���G� m�7vU��Ο�A��#���2�Zs>vq6��h��v��~�Uen@����I��h;��YZs��AN}(��<�i��oV����b��i�H��;$:cH��xJU�0�����Bm�-%|6���7[�^�N n�d��(�F)ȡ���}��	�4�énc�9�=�HlS\"E}��0iD��Ce$嚎��?��3�b��L���d�~��iJe���8T�#@^��^�rm�7!7��Q��+ 9�\�Ke��c��9�
����	���rj֡H���C��7o)��;"�����	�sD��bt���.��t��le�����ǔ��qK"�f?�M��˲N�
�<Հ :�O�k��|ܠ4��Yӓ\���|JS{@���Ԑ����5H
�V!�1]]_=�*�J����ؐw�^��&�b��?����iD�SkHp�aw�10���@�`1u�O���֒�Aͷ4{l%N�o����\�����g&�<6&����5{�_S
 �����S_������2�'� ����� *�(2�})���vH��eʛ3���_����@v�a��qz_7�T�h���i	������> ��3b�ҭ�G�C!1�E��U)��굎�U�ôr/�^-q-���f�a�T��;y�	�ʅ�ĝTBs3�r��j	eeO$ΫveXwI���+ԇD`��HX�o��������zR^�9�-R�ü`\W��dN�&v$uy���)�@.+�UR{l��A�W��ġ��-˜�dDp8��o}l}9���rh����j�b3Gz�7S��Sk.��|5�s*�v�םDO}����p�7TK��/�2)�4��z�!�9��)��uJjU�ٵ�$��-�"�;�����y���.Et�*�d�8���
a�H&tF��o���Ѹ� 0��Rm�@��TwgG�;��6#�qk?��47!�E�����&2�H>"�[��A�i��iM�f.����j7�5ëoX�'RNv��w y]�eLK��p��'Ħ�*��1fo_X��?򑗒�e�T˪M/?��؀�m���T;L>;!��K0��&�|�?�C;%� '�,,�06���!M|�y��h�F�r��" �+B��j��6 '�x��*�8�� )؋�(w�#�7�j�M���)B�A�YwA!���N�60��<��V�K��uF�[���q�>�eN$k&���bO:{h4�r�s�k��8��¾�5h'�f"r9�BB���P��0W�s��_�����hhI�+ڄ��^���L햹�A�ޟ���{��m�	��,��Y�\��K���<�U�dIb�~�ß�M�l=<B�5J`�!�Q�'�p,Y�$�� ]�p	gC@��&�=�\1f�"(�7��*�����c|�&ǌ��� �If&	����{L���0b���N��w�
�}*)��_B�ϵ�js�f@�uzChE#�X��^q���:���}��� lz����Xp0q��GJ��>��]��-e^����T/����Q�}�٤1��6?#?�����(�Qq�2N5R�ke{��_rʞ=5�ִ�C���<�V�-�u������V�_XO_���b����N���V9��8�cH�ߨ��
d�T�6�y����MUE!��J/m���[���Z-�UB�b�Dj5H�z�4��?�,>dϳ�L�%1���>���|��|����I,���J�M��j���1�拃�Š�	�e�j����&W,�m�Q�}`��W,$/�k��_"E�F�1� ����h��hS��\?mQ(A��y,�N���l����W�{L7���f�ر������`ԯ�&�;��4M���E=+h�L;�8c2=ңл���'���sO�d'#O�3�=(�U��ՅO�(*��B���B���ċ��q�Gq7�kg�I�_�K��iH<�v��o��'��Y��e��`LמI�lO�Ɠ���Z<��!�R���ɯ7��FEqn1�����i���
|4�8M��1�[��WFi��ݯ)�Z�	K�_\a��I����rN�����)������-����|�����s���{��XI��NAJ�*��g�^9��%��T��v]��F��g��i�f�����Ӑ7�W�꼨M��]��&�HK�Y�Mt���^��e� �T�D@���-	��Y*�� e��?�V�ЧAT%V�7w^��D5�I�Iw�nܑ�a�p��_J汢�TWk^R��A=��B�8�p�X�E+��\�R0n&���h
_p?�>�a���0�=2�"4�� *y���F{��ul5����R�+=�����ȅ�ݽ��^Z��*� >�o������;@�� �ɐD<�\'Sd0�"��5݉��3�S��������ȕ�K짞�"*�N��U?O"�����I��AW�'�0:Z���i`��M�ʡ&Q1��w7���l���=}��ĵ�(tz��^&�E���Q��BM�8���Vro��M�_��6Vؓ1�ۉ�I|��M���=8���eHz]N��&��N��E@�^�����	B0<��0�(\�oЬWi���Z��H�'Y���搆FC5J�ZI�2+����/6N�	B��sn�]U'Q�v��3������Qsi� "r{;����>�㋭?�{��3R��q���yf�ղ��-�� �k6�<'���k�e,���zT�\/��~#L5�|�Y�0�lH3x/�c�k�K%�]���~�B� 	5�.�C�"F\�+]X���w��gK�<�X��a�l^;������|�ޔ�t�"',w��t+kf��b�$��|����.���Z��myΦ>X$�?=Z-�@�;h,\����Y�^�EF'vc}��·��3�n�#�'��Ș��]6�{�?��woB%C��Wv��@�Aܰ����'-�O"�3&�X�0��O��_(f��$��0-n�n���_��?���d�o��K
5j���Z8QB�I?�w�/��8���3lu��Y��CUİ�%ʰ�* [���*#2sh/��;*���TU���V'?ݾ������y��ird�~��)P�͛�\)��T܍	S1ǀ�Y��E�MU������<'�����4+���-yu�!�Q�e��d�q�Us�͵���^?�5r�F�,��v�t��
v�u�x'�QX7�ɥe����p�E2
��g83|D��.��uUu�7�,&x�Y�X��Tȏ�nl��J�������v������� �ӄF*9B���#����~Y%�ogz�u�K��zw�kc����򦓈Y��q���E4�Si��.��F��.�	e#5������Z��(t���1�3���Jlzc���*��Xtk?gO��,�[��7^t1ZS
a�;l=?*���Tg�a�F�z\󐡀Lkr�r��_����|� 5w�$��MC�8^�q-J���ʒ���O���$�Y5*$�#��UJ�-��Y����o�����vo&�Ⳬ�8c["��vtM��*��U H�M���*mU�� �+�2�����������_B=�^�;X�.�(�ద�C��ߣ�X ygIJ�Oe�~i�&�|.��o�n�k9��վ\�����d����q����F9���ޓ%�R��,�dR#��	ٹ�
ת�a)��IZ2R�B��Np��r��d�j?w��,:\L��R�ϯH������-v����y~@�Ϻ#>�>ke���>�r6t���T�*Q��^�]�]�B�O/���ǅs�"R�lB�k�W,"��bOm�n����	n,�p/�Z���̝����pA���h��	'#��Պ'I�l
U���KX|���L��߂�R�#2�r�s��cgv�uչYğ����Dm�A�p`58�g�y�z
��&��x��C
<vG|�rBQ9���5�bo�Fh�YAO�@V�6B��}y�C�F������t�:�k��$����d����� �|�[@������CQB���)ء�>�w&]Xn�W��/������y�ϱQ��ƫ���<�N0A��b�vp��p0�q�h��Ʈ��s��Š����6��
���뗥��s�xӚ�+���*P�"�Re�`v�|��t��r=Ι"�mh�p�g��f���ɢ|����s�^~�+-����^7����>�~|i��Ћ�ƽ�e=��z���a�Y�2��(,ō�9m��:u^'sH�o������Y"+CS>T;�e����l"4��;�	G�I�.ن`W���G�{�}f���ԅ:����b�GE�L�G���~9<n��WJ1UcZ6|>% Im�ge��`������T���Eq��܇\�(�{}H8ٽ�fkP��+ ���x�:�F�v�ͦ�{��Y���>;` mѬ�s�ݷ#ikps�����t�,-,�?�eF��\:�|�I�_��ui��;�돢��;��M���:M4���o6�т���:���7;ǣ��M�����)�������9=p�����\C2&�*)R��`mh^�(E�PK���Bv+���F�ǳMH���(���"6[�d{ �c��o�<(d@f�����Y~:�n�mn� >~�sl��l����h3Y���ܮ;��,��a(�`9jV�L�x9-�m'�~<�[��c�r���pڢ%c��D�^�*�IJӧ:� ��p
N�Emm��{���Ȉ8
i��ncu��O�tx�ǈ��P�_��T���+'�K�č�|A�p�z~��lж����q��$�����Y�ko�<��:У����ˑ��.���,�j�B���.MB�?;�gͥ٠�Ɵ���Bj���E�������.�K��$��9������������=� �x� _y�X~�>��c>O����'��ب~ߍ�0�[>���j9mdƦ-Lr(�{���BC�O���7 $�}�j�4�����#��nfKXd��1�1��W��6/�D��K}�x;$�װQr 9-����ϗk
��N��@.��,��ܻ2r��Y+���M�&����t_�.�r�����D�˴b���F���|L�����NZ��D�z��j]?�O;Q���c(M�-D��K0,�Σ8�LE�G:J����ƛ��\�|��r�����h�/��)�z�d�I�iM�	 �/5�i�4�=!�=o�]�Q�:#Y17/)�<�O�LQ�������r{�("s�P؎R�*P����#Ӫ?U��T�'�=cR�5�O�P��~A�"���+A��P�}�Q�O{�Dt��B��z��9Q -�vu,f'D����^ �p�rLݻ�U�2��xI��TT*��� �H������N\��\�
����/����R6�e�{�c��4������1�X���9��)�EF���p���.F���G��Ff� ��_���j�!r��%��, ��֙3���X�h㕅;����}Ă�+��FQ,��ZOa%��f�P&]Tl�8����	� H�Sͫ��5ѭ� �[�f�ˠ��B�^e�ŋ��\����r�iI3��Y���VVQ̕R�:�'S�La�'��H��@D���/��[Dx�l{�)_Ж�9��|4j�6t"��oy�7rm�����uj''����,���#��������{;.��k�e��Il�a�X`�+m #�VZ�Lc.�݉&}������>�
$8Q��M�;@c���S�q	u���,�4ˍam�׼4i����lw2G�U�t�ֻ�`�&��/�@$��@��n�" � ���8���7-��|l����2�EJ�H'����<�%�H�Q��G���GTUc��j�d��$`Ta0�i�eL+Z�?�2s���������r�e�|��_�u��X^�nᨃ�a6�9�M�#{ԝ��9@4	���W
�n����hFIg#���.�������eͼ�qpa�
���8l6�t��,id��6����L<�(�M��`����6_l0\�ݼ�R�g�?�͛�k�bQ2 ��V���q/Z��h��`4v�h�y�n �-�X$�.����C�OV������|�V�Fx�p&V)J"Sg��gFi_��Ƃ�?��c	�y� �0Lti��3����
KYq�xb���șv_����(>���-�*����-����1�@�=�S�%iCb����BC�x��Kx�4b�3��S�d�U�ԑep���+��Ԟ3G�w`�7Z�3ߙ#�at�:^�����4��"���@Qf�%��t���1��4{R�ZM�*��d�O5n7j���^�����Y�5�N+R����3�8����(���wT�p��4EU�=��*Ф���f�v��D�A|=~t7�V��ii����.]��2^}qn�g�hd@�ۑ.���W�J?�nsB+��`�DvX�}!;͗%���#{'��169A+vʓ���r�б��7�W�ٹ�P��ȏ�D)_����� I����l&�p#���[��9M6���M,%��)�t��x`�Ŭo:�M�Wa�%2�����94F��>��U�a������玕�-ff� �Ҽ������q�$��W������k�B/���Z��1�:Z�Mo�lU_r��d��>���9�K�}E ��"�P
�=jx�Q��q���K���ʼUݵ馠��R�c_�#�ՎOףE ��~�3#�)ԗ��i�P�b������U�����M��7���Exm�=c��TEF�v����z^�$!a����d�:��������js�V�.;t�����g��������cG�dv�!ا��q���K�,?P�
��"v�'�7k��V��cy酓���
�C�b%��-�%ai��v��E�����47��ݮ�KB
��n���7�]���?���9�HT�z�����H�Br�f�[��[n����pZ?��3�d�!�2H	�>��q����H(j�Ƨ��U��)��"�TF17B�j�{e����/]¨�}pNJ��}_{�rA�_
�j���~� Sx���OI����3�[���E�9�vf!U��m�%�o�*�_�&Q7 ��E�?�^9�O�?�'�7iaH�dr��G�h�r9�y�%Cj�輣�����2-��F&�hY��\5cX���A�%㔬�X���\�``��G�}�8��R�G�W{�� ��{E�斠W�����=�hO"+0|�1E��Q���o�v-����A�}��+���q�7Hf�J���(锄=峄E�vB%�|D8�xd�O0����1���6��Q s���چ�+d�� ��`��#��w=^Q'�f�}�͆ 8��X����Btɨ����冨��K�>�s2��Xb�)|hJ�2����$	b�eR�V�y��&hG�� 3�&Z;I�g�A�ʚ[��;I�ݽ�2l�򏂔.�66��g�-aPA��Y�(��Q2�-�7U�V����k?;��<�p�%���1�+