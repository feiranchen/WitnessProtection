��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��=u��*QZȗ�/�fig��v@�g�v��9��~��=]b͆�XN�i�����N�hDX�`�9ƚ�$X� �H���>��}�@�lp�Pc7 ����3�lc\���R0��HG�[��/d	�7��T:v+ȑa	0�>��t�����F�}<�д�scزg�L�~����'��t��]N��R/�m��ٌr�"}ۇ��dYrN�%��S�����v��\k�O_�*1!�U4(k!m+��$��s���Z7�W"����/7��8r`v��v��8Ua���/�Bߋ"h���5�Yz`��p���=�PZC��U���J����0WP��@;��9M�Z�_z;��tO�J�J}�^Qz�yD6�&�6���!q���9:Oę�Gu]KQ���d��oG��{;�oY�-��>t["嚤�y�v�Z,f���&�ml\��#j�y_�\N,X1-�kf�����ߔ+ڼG=��{ٚĉ�d}�E#�.v��G�B9��2�Hm/�2B ng�:�,�Ϟ�NR-���;w����.�}�\�lj	�w<����,�B����y��e����L2���,	��bw�0%'�|���\"�!"����$2�Sg�mlxc}/uƙJZ��Bg�_đr=' �lN����H��b{��
�ԡk�]��<@�?O\��w)��9�/#�Tz��n�-UB�� �p�)���H[ɬDT��������#�
�D%�&�z�s��J������� C�b��s�j���/�|��vI+���=pL]�A���o��N���ѷ^���hj3M��_���I���t��2�+���p�PF�¤Mk$jf��D��B-�g����:완�[�U�\9HǗ�J�#B(xI�s�θL];�����lQ�֑�.�^��l�#�	�>1(�D���\�s{�(6�a)��/}�3���c�h�!ŴG3y��6����Zz��ɯ^@y�r��Kk��D�.��@`�Fi����|x��R��8���k��:� �]#&��V����j��%���x�����`2HԽ��g�r����g�1��������φ��u��v&�+T(��K�GO���v�9�ۯ������>�#��� �F��Ȧ��ە-�K���l���o|bġ�9KO���'G�D��V��{�2�2�F��Pt���H���Yj7��8�>�k�F�.�C�����+W�8�域��F��Z�V �3{d��ũ��8��,SS�JxUXMv��L���r߭�'�&2Qð��b)�X�͚��ui�n^`��Uh�P���z
�e!���̯T��<��]P*�e��;���5x�\��9�q!�Yמ��0p��:��j"}�0��02f�ln�hT���$����ZW3�]f=:G�V�gP��"�
��V�
v����KՕ�I����mėz�H��qI��Z�PV�9���8�Zc]-*}�i;��b={e����:���x���s/}����
<��vn@�r�����୚�)�1�2d���<uy��[y(��r=\�Yj�{�����C'kIR(]�@w8��|�I
ʾK���m���$��,h��Q�Ja�����)-�p8�H���NO���U��D�{�+�k
~�Q������'`�p:��B �aW�q^�_�0��-�>���6G��*J ���n(�}1��g
e��˘+�t;�ep�\Q�����Z(�H-7e��
�e��T�y���m�v'�[r��R��N�K=b�(�ୁ��%,����pB�����S�K:�v�{�h����'�6�)��H<UՕ,���	_������̎HQ�~��ng���������;�%��:����!F�T���i<Z}������J&���Jc��[�)]E�,yc��Fc,@��	�p��I��g6ǵB\R����e������#8��̿�_.k�>������*��Nw��f[��N����mM��g�c�k��\�����!4˾$ie������t�Z��P1ܨƗ�*(©0�Sb<t�����W4$V�m΁?\�
���1����ԇ�j �;�_��% o���
&�5�<��������a�-�R�����1�	}!c��/N�vWeMM��45��������. �0,�t<)&T��0��!���ŇK�:��3�}���Z��RN�J>R�1:y�x���ʫ�0�qV���ɢ|���h��_帬�=d��������e�AC��z-.]4s@_����C�n��ZY�g�w�,�P�q:W:������yv�y{����bM����������#>�_���D�3�A�e�}@�nANZ�^��1���(3�7�s__P�*�ϱ_#՚�Bx4z�s�C��P���\��IZ��QW�j#&���O����jd��G(��bh���.����~0���k�Ve!�O�a�yf��tq�G�z:P��E�n=�a��������tፙ�i*�)�����D������cf��+o!.e�!���\RU�y�_2z�m�2P��t���+���������<��s
�r�z����$R��A{�U����5-���G�e��z�_�(�?��l�M3"*S�I賧�;'�>e?�W"�IL?�x{[�Һ���1_3���ŵ�T��V�WBf>5�j���]�F��d�e���
�;���ZXE��&J:57���7��ˊ�� �q��L-���1��%�>}Љ�/hL���0 T஝���uq��o�Up�mQg�Y�����LV���C��C&��k�s�.ʬ�d��t�tn�<���m����5�Ř3��`��%��]����K+)^��%��[�{(�� �La���F�͘�d��"_G0�_�1����=;�'�[�c�I&�kʥ
x}<w�W(����%��2d�r�b�,�`���4"ۏ�l��pO�m��H5�Ѽo�i+�U�8�Uyp2e�@-`��2����p��F�
3i_�|s� ���c���W�0,�����q�nm��É��M����!�fgK�F"&�*&��T�g�+�]tV��lF�	hW~��!՚=ƿ����m�0J6�)���*�Ql�o��D�% w@&��D��[�$��WÄ�93�!~v�wʟﻢ�F>h����<��uN�*\��O��>�;+��f]�j�X��d�A�#пx����oT,��.�uk�' '~�hYM��o���2v%e�&p�򥻑|x�BѲFm`��d��������S�1��J���&2�͒۝T�x0���qS:�r↏�/��8��j�697êh��3�Aa���(��u�+ɲ3M)q��;�>qi�71�.�=(CX��7�q
�v����<����3h��Rb=A��� ���|ėnL\�r����r�?���l��X�(�5�%	�����9���˪���*@����j�MiC[n�h�)�GEμ���o�
֯vMAƠ>RNn*��)w-���D�Νz�3�J"��������&�U���9?��h�ar4V��bɾw�81y�W�L�鑙����j`���HK��֣�O����VF�H++�l�ꚙ�,�7�8��'v ��Py�ǈ+���ڧ����
`O�L8xBvw��H_��\7��<��lg\Ó�H��ɹ*�L�%яK�ba�ɐ0��a3]7�Zx�p��RX��Sa�Ã'{,�RA��ݼ̀�ߗɏ��߳�%������[����_Q��Z�1u���r����9boE���a��Z7|�O��l�G�.�$��Ƹ���US��kmc�P�G%ˣd+��Aks^L3J���?"U�E���{� >^Xy�W��ZK ��M���l���WѦ�~v���^��ɚѪ��3���ֽUν�Vq�8��R����ŐA�w1�O����R��#�y�v� ��O�q?
T�]�1 !�P�B����5B�F���r0x �6��l��l�PS ��ލ�V�h�w��T�uGoX��E�/�z�6�|7ߴ1����I�t�ћJ�i�sJ�3LЂ���T�S��Jd8�a�6�11̏c��hϏ���Ħ��'�p�.u3|󝷥�ߠ,Ո ۔-}>_2)��_������!�9�����A�~Bꂙ�{P�MD���j]���c�X{F�K�ވ��Vh+�4F�\7�6CP�,�p!��zk| {��C�sh��S�1�,OU���Yźv��DK4[R1��ξ���V�[�����jfM��?�ԉ���A)$�U}��ha����Dp���K�4�t��*���k�31`��ΰE����_L��6)��� ��	�h��[���ϙޘ?�w'4�4�k�(<�m���>�Aڲ%�~����F6�M����Y祆0�0oTD��8�}�ن�~��(Zt%%j�H�FsC����GT�F��Hsc_	U(/ݙ���ǐ�m�)6�5lf��@/PxT߂�ʽk,//Y�øK��yF�y� ݲ�~l�����٨�8O��z��R���[���\A<�"���a�k�\+܌.��o�ilGC��v�/>ku����Jdi�[������t	95���� ~X�3̺!'�c�ߟ���Iv��Q�D�� ��3��,�B}�{GZp������er���nQ�@@(�\.�qS�P����2���$�5g�Q�إ����>�³��OVU�IĕZM��V-eg`�GC���'��o-��iŕ��r�*��ɘ����S��k�� ?)D�
��>�v�i���d 9���d�[�:�
V��CR�820B�7�W��`�n3�V��pc_��0��fxж�?K��tm������״�,��g�onҫ&px2�=s����������硼:��Jˈ
�4��?îE�A���MIw��2��������=u���f���ۿg���������Z���N�_ӥ�{1�_�L#���U���Q�%C���Z\2�
OE9�����D/�V����cQ�T�Xf�XWiWr{�䬃�����G�+���V �:��*��a��!��I`�~[F|�[`'�ʮ���M��y��4��m���F��錎 �p�zw�|1|VLVoȜS���Q��W�"�P[Sn`)6���^I�'�ȝ�p�� �{���v�8qgu�H�Jf�f!��W��|�9�}g�����B��dρ.B	�V�EG0}�3<։�j�Qe�ڻ%�	r�b�b*0��:�*�en��g#�X>��uC�D�?)W�����&�cS(o~�C��aO�JB�ꭉC_�T�Q�DDʥ4� R�)�d��A݁Z{�N���=��9dT�:r6֐�}l�#��k�%�e�[�ܥq�Z��Q~m]>�K͏��hL�x�ֳUf�vsL�)+��(?x�))��~)�
^��������\�͖*
mU�=��P�̱<Ey����{;�j1]�9Xl�S�@��v���+�j�!+����q~��|q�~��������) U��ӛ�]2��լ'��1�c}_gf���t�"�b�,��J`���Ӽ��HFi�+��y�9�K �7�� M��1�!|�OMUN02'4P���fқW��_	��f�"hT&�%xtŚH��HY��DE�%�K-��?�5���iz�Z\54n���>�J�,Iw����e#���3a{��0����lfw7\�ˠ�J���0��m`�mU����a_
��F7:�e��ͭ�6��"ót;bn����˦�	y����q[�>�2e]��Tg_��V�����{���D���ڽ ��'R�M�竘��EE�4�Z�*��Hd�U_�)��ל�9 T���o�,� ��q.者p�4u�S�������#SDg��[z%0�� ࠰�4����>��y=ۅM{�p�{�ܣ#�*:��c:�L�@��ϑ�R,G�69Om�����Q�m�z�5p�l�]����؜:�F(b����ݎ���z�n�� �d_�����;n�Zк�����gZ��o)�h��yuA�#$&����.?��U.cZ-���^�g�a�>�G�l.����wz���EgET46NS���K��f^�(�n���x����ULC.7��Q�����*�U��+�&#��ZGS�(��F�E�L��|�f�~�uA�f��g���τW	�
���;7�w���m�"��R�rF�3\{wo�)e4���+�p���N�6.&�+Su��$��ю�����~ɅE�"UC5��(�?_#�>��'�ESG%:�秜��鷀^�͓dE],6ê�yn�K��O�c���ס���^�-5��y9b�db%�Zf���J���E�loD+�)��
ʵ�6�N� �`ې�]!��<�[@��2 �R��	{�W׍H�No�Q�I1\�0x�G6 };T�_mJ�nW�(6��l��Η�c��6ڒ%��+|.����uTq�cOC�
�� �6>J���~ޖ�9����R �'�`2� QH�ٖ�)z|�`� Xw!u�8�k���ɣ��P�sz�����O������e7�y�bN��@�{F���h*��!�Rozne�������¹Vk&!p���8����W��<w�/����\��	
\u�!�������
�s��׻����,\���Ո� @D��B�.���n���H�'m��vP7��]���o��g Tb�~h)�g�N��H�5��`� N�w����ʗ`�㠄u��ԚBL(wH��S��֏n5j���dp�HRr7bT6�+D�U<���-� �!н��8�_�0�+X2;�����o�"���[����;b�_T���W�Eщ>�mbs�N�b�z���mё��Q����O�����`Z.�� �n�4�2�a���4�~+�����r:���Qb!U�E�+��	G��l�h�j�5����CR���P��]��?e��ܫ�8;�i;۠~��}{�=��|!\@dK�Q/c�Z8.�>4� �y�c�,cE�*k�[^��{M8�[�ko�-Q����j���,^n�_H�ʕ���&8{2�#=E�O��o�oLw/5!%ZP�M�v�=�5!ԧ3p|�_C�h
R�6��I:���	�޶���S��r�bx\Q��uh v�~܀�
�+n�k4�d�R�����s��(�Չ7S
P��A8IP���TJ7I�gژ�ld3�/au�IM^r?�zN��`!N��Ym����д2��[٢u�������nR*#�ĹǨ�#,/��P���%�/v���J���
"~a�W4֒Է��S��\!"thL3���d����@�ǫ�8Ũ��x���>Ʈ�0r��R�9�Y��%��6��|رE�@t;ڟ'��Л�����II��}�sH.����E�q� ����'�_2?���&�t�c���*K�>W��2^瓞�K��ֻ�;2���3����G%�'�����6�|rvM�C�v�0iU)���}0�Π�^#|�Ik����W��eCݱ �@?� �n�݀�(��'�\Q��RJ2��9�u[�fuV�w8
�?v�:%�	NAO(תCp��P���Y�ۛ�>�S���eg��c#�+d7�a�ݤ��� ,m�܋>f��R����Ԝ�n�`g�VWO0�i�%��x�mS���u�L�AҪ	�|�.'��������Q�X�U�V�"�����i�j�p��D`8��^x��\�+���L񿕺VGJ?;���I�ƊJ����(���p�M���v{~�j��)�6���h-�$B�xm�:�]�8�G�B���%� ���)\��^������bX�kgŐ��a=���c��|"�jKx����EzR�dLCt�e3A����I�X0�<f]bH��]���M8@�iFp%'T�8����BM/������ĹD��njH|n���i\r�-��N�j��h�]X"���?�dMo� ����L�;�tp6>�I,CS��R9��`:<&κhDb6v��$<���[:�X-����m�1-�s�}-1�7��r!
�k���[fߊ�\�V������)�����HT�P:D�Or��+A9y�'��:���jqy�[H�W�R_ZHP,:��;�*�h/Y��"}I�E��1�2&��H��k;��)��ڼ]��S	فgr�L���;��������M��C2�2���*W��J�C.yc"�Ҁ��A6��ԙS&U�n՝��4� � F��`��sꦍJ6�y��3&ƿ�N��r"C\���	m�J�> D����7b4g��ܤ�n�e�H�1>��]0��@_�`+زK(0���12k���!�.�3��D���[o�$�$[9����tm=
��`O�؍ԓ�@ҷ�(���ݳ����x�U�����+��7}y�<�^S���:ȅO�?���E,e�̧j�� r�����Pi!u��`} ����R}i0Ł�Pf+\�4a�ō�f����[}�P=��}5���C�ߩ�5t�����D> �2q�+�LK�_�'���;�A�/*��
�d��V����n��r�u��=Ҥ��ǐxb�W,�i��Mz�6-3֖�RsF�J����ˊ^f���%�@S���}4�E��M|u���̻����pkg.֓�Ѽ�%��i��XEL-�7���0�K5�1:إ���5u�O?%�
���bP>�/�rL�"*��I{iF�
:��JHF@�0�е�0.�K8��+���E{W��.EM��3�3��3b��m�ם0F�a�-0Վxl�My�P�(*�C�I_P��>37�@���]a仰��'���d� {��3^��S���n�+ܕB��Q�Uw��ojS�^�&{��e��Q���ȩ(M�RQj���Q�O�b{�i5f^���&���|e<}cPp"���{�2��s\�6���G�fp3���!�y�q�OY-#�91Tu��'������h�3@�\jB�`�@�p����=�]�%��O�aT��0k�ޅ���Zn��'�;�.�<i ����.��@���p� �w�ヲ���)_���0 ��r�N� �02<�}���9�TrqN�fk, �:LZ;D��+�x��tq)Y *F�䈓�|��I���T��ͭ�4<6&��mR�x���le]��}A�M�&5����_	H@��r&�����@z��j�yz�n6)�n��XP��iϝ�JDߪ�(ڜMr�b��ɍ} ߔ��Y�XlD����ZT�Q0�dkP-�#hj�O�y�7�0�Ax�L>���(Gp�
�7�$����;����[���6��;��/��#BX����\�&J��?�=����~���w���Bձ�&�~y��'����wQ>L��#7��S(�c�y���i�U����4*n��-��z��x������c�9�bD���z
�A@����{P�
9S]!;�@�dq�ȑ�%fL�H���BIɊ<[��p������Ȗ�H�b��k��m�/1kVL�T�j�����_�D���t��V�����OO���o4d�q����|���:�ܜ������%d��e�!F���옙�Y�\�Ǝ'{Ѽ��CR���s���tV+��c������T��,~�J�o��8E�?z�k	�|��|ҿ�D��\��0����ԁ%�и�T�5U����_99՛��:Ə��q�倖x ����>(x�h�������)>!��!��I�5'������;�U�*y�,SHhb�)�!���չ�^�Q���D�,|ۄJ�oLb�-!>Tʜ�3M�
����O7��$`��HI<q�o=�f[΍8�MW����� 2�8Q0DJ�:�?�Q<��Z �#��Q{���DG�0#�B~bib���^���磬��$}�{����ڤ#x�� )d��HH����1�D�C8���Y�ߦ���A��j=�k�d������>�N`������ذ(�O�r�>�4�R��� ,$��1֝��%��[��Y4�Ж�mt`����'?��s�|�ѱ,��^RC�=�}S�;�+�A-Λ���ߓ��%��s]-r�ɣ�9F�V%X��u���
ݍX$�x
��e��3�R�����4�j,���:���f:��C%���>��B�_�X����R�[Mg����Jy�P|��_��^!8�.<N��Q�f-O�W`�=��tm�K��i�	F*�l���N@ �u"�l�
EZ���[��+-���	!\gC��~��<.TZ@wt�_�4��A���i@�өZF�����M��#C���`���ڍB����PZ�O0Q�f`;ۧ�k|��ߗb5Go�:	���{�;�b:?/h3D��4/ehe�T�rX�f�"�ex��US����
j��H~�A��E΂�6�3�?�&��v\Ϥ#���$Y��T��#1d���o�/��DJ1�U3`MhcA/0h�����v��jD���>�\#� $��\R�A�=���� �S�T^o��p2P��BA��l����y4p&�N�+�3X�]����\eI������K����"a�e��� �ӋG�k��EZ����SecP��:�I���U3 9۰;=l�<,͵"ŝ�
Fy(�}��4�92$������Ez��r�LM��<7E}U@��boL�`�����|eu�[nH4�9}ԙ� mI����,�tJ��錨ƢFPa� :��0��
��X����چчr^4{�ev�%��q2���;��(����Mlk7'J�w�������U�<���I��D��(�Λ�a�)����n1��w껺�=s��7�Z%�<��GI�,���PI@����~6�,�@��L�(5G��i��_Ô [�����I��ѣ�F��I�=��L]��Z�>���7��S3i�S�:���� �{A���OdU�T]�&Z���e��"n��FĥO��R��҈]�_�: Abl��G��>�)�U�����ƴj|j8������@�D��6���Z�[%p�{�x��=��X�u"9��F�����v���S�7k�\�*u<[%���ym4��HV�O�H<&K�9�̮��׼��	Jo��F�U�0g���!U|���"g��d¤^=�@K�l�%$���t����a�E�gt+��lt�����ދ�f�\����� �I�3�t���|�.�(����[�BF)�]�Έ;AG&���Io*&�V*� E+λIJ ��^�O��W&�כY{��H��F�
f�<��k|`�{�S��p|���l����*���1aH�;"���8��xw�6���&�R8���"�L�{�SԴQi�O)�)n�f��������I�m��2uX��%ISSS�����WG O�5C�j�]iX��Ն�bb�1��r�r���%L�7��iy��h�����Q~B����4-���v�n~�F�z��|�n8[|ܟ��X��a.ƚڱ�h�B�	,�]Q��9wT$f����, ���T�V����=����ߔ9DlF�ִ��+H�B�����l�țЎ3Uj��m�ɲHK2�3�2�*FZl*#��bڝ`�ؠ�`�vl���d�����΁4�X��%��(ԟx�IBIB�g�*8��PTpp�Qpz���?W�M���p�k���9ㇲoMk�!�gP�� ����RI�̩ǿ�2����(�Ėę(0Hm�!^�`�K�
�� uE~�C������$�@`���8n
@;~���(�E�7�h=����Nm���z�0��ڔ�}�s��z��	D'�gkE׵6�絊�#g(]��s������5���ٿ�R�u���6v�\��+NL%����y��wk{�;��%ލD*�gХ/h�"7-�-��?�,e���Ue$�L?b��n���6����s�����H�Mʍ?�u���e$]��m�n�7S> �c�������?i!m�?F��J�j9�n�g�.uX���>��X\�.��jSl|�IX�o�dv�yJ݈�Ѻ�_O֓��Ǉ����	�0���Ka$��T���;<��!R>0��˜���g���S��A�F� 1���O�B��Gi%���]��q8��a�KY^�H����S*��ne��D�U���h{��H���w�5x@� ��6|�H�?݉�1U�O������a�_2A���]3Ue7h��m��JM3(�j�c�h���@~�]������~*{6A��ZBFG�P��/��z{�e�u��2�^̿��������4����g4���6�N'M��鳡�r�K�k1w�&����;k��خ���b�f4�tNj��+�Lڙ6YY��W4�O�D���:*��w2Un~"ܩ+�]Ş�],i��&~?�S/�%%�Sܗ�l2�:���ٟCfV�Ԁb���0G$�*�T����ˎ����p��:ZYg�S�g�joK�u���#�Cz}�;E:��b�����mja�������y�Y�&̎�{�\~��Fe=�Z����f��oe%��bW�|sՅ��ק� ��@:0��z��|
�M��i�JP�6�լ���;�+=RB[�pG#��J%ψ� U���"gm\�x�O7}_}�>�뺄�'�"/�_:8�soO����a�?Sʼ���kKEsg�蜱����?� �(b�9����� �p�-�0�,��GUQ1ޗ�٢�W��<|UA��"�1��4��`qS>�Nh�#�("ż�׬T�)����ʠ O���q�R�xp���8�TssN�c�;����u�2��">�Lk�,��ABۊ0�E��Q�	v��(	-G:s��RRP���%���L3�aۻ�����؝�6�:Eq��)��t��W��3?��+���4t��7w���u��:@)�b� �8�]����_=9���ެ�e��s�4��U`Qi����̨�vx��|�h�Օ��݃����Sߧn8^�=,�{�5w��rH`��[��'�����[w{ޫޅ����W����j�@Ξ�3ȡ��P�I�V��NmV&� �'YAJ��$k��M���v�j��ߒ���NL�KKֺ}H���2\�i���8�tB��R<��V��iEO]��T�"���b'��v��O"zM��~s�����`���A7f�]��Dv9��y��_�H�#VX5t�S�FbkG�+�G��_V�0�X`���8t�������Ѧ�� T^��aW���=�l;�y�5�=�{x^N0�sP��'��;�p���;31cG�ש� ��>��n��֚}��q(����<�����	�Y�疅?!�C��v:?:!���J�M�����gl5�[�F�%�_򦴻$��c��N��P\8;�]UN!�K`y�������nn'�ҳ���d ,&�~Q�8h��	�	l�5�������lWG��z��G������wڐe�4����YzucO?X�΢��l����I�X]���4��6X��p���a�k�c��1R�b��c��HK�� �����M���kd�o$���H�*�j���һߋ�7[>�S
Ore��P��O�A�&��!���?�}Gl[(X�A0�S�b�8���`�����,�g����}Ƽ����a��5Z�a_QNd��юq1 P=�"xA��?��'_���}p���,��j_y"��!-\���L�u}����D=A�ο���凲�������% k���N�
���a�t��,3��C��戆Ƈ�@?�o��j���Ǣd�F���\��Lc����+������Y @mE��[��j�� Y�D/��]��(�o�xA����֍L���o�d�?V�������<����]?wɮb>�J)	]��Ȕ��;?% H�f���5N�=���+�qV�T����������"��a=��(^Yx���j�|�)��En�B.�[v�Z���X^��Wq%���N��]*�K}�uMۻ��tLj^_��U��y�͖����\d�����FW���I��K1R�24��q�y��aC�	������GM,��y��<WSm�h�')!	��؍i��l�V��kō���c���F"�ן�����U�N��:m�t_
��*}�_�"p�-��6�ٽE[Y�� �hΝt�XM��cK��D�*�( C"��5�d���;���CU����vd7��j��i��b�}�#��<��J�4�&��-M��Ίz�uX�����XG���I+�7D/�k�Mx%����T��ފ,3��뀼e-��d�/9.�d�쬱r,�@`��S �KO�V���X%�!����6�>l����w���;��i��nH�w3�_!���۷@����*�ս8�SF^�h�NA�]��+�͡wyg$�����v�"HSu�0l�Me�6э��)W!X��2�ahֶ�0TP���/]���T7�!�ʜa���®?������~7�Q; �Ѣ��2b��4Xv�V�}U�)f�i8U㡉�+6򱰚i�'k�sڬ�t����ot��Cض.)���By�X,g�Y��*n>d'�d���R����L�ގ�?�'��m��f�03���?|�>%4�5�c�%��(N�q:M�ߔ�*@�_�2,`�G~>�(�����N1�qޭ�z��xN�ߦ�Y���]ׯ�7-�L���a ���	����dG,o���-qQ��"T1	��X>$��o��ɤI?#���g=�jTtB��ZdwY���D�Ow�z9��-� �ɟ�3���o��X�ʢ�~��=�y��W�~�t:�kY��:��W����K�6��c»�K{��~Z���?j�v��nr֭�cD^d��iۅ��HW�x��
-��������P���v�u���!+�g���0e�t#��ިM�M6� �x���}:OK@��ix��Y����9�������=,z�����E���`�RVқ`���a�9����Nlu�����5�Nyh�/.�ð��qI��u�����\|�3a�d���c)�4�7%�9��i�;RL@��`���4��I:8 ���'[��I�wx1;��H�8=$]��8���OAPvgEX/��a�M�����\
������Mֲln?��_�2^����ZH%�~�W^�8>K�Pȼ������0�q$-c�Mz������N�88��f2R_U��"����ۥf�bX��i���R�m����Y:�#}�bt-hIy�x�|�ZZG��m/"p�͢��dF�0��{���&y;u����;l������J}yU���&�����]1��	Q}z��,N�
C�Kg��.6:��.�[��^X��H�P����`a��p�V쳍-�GS��+��aOa��k�����C�twx�%����4~������Z+����F.�w����;�V�$�u�*���Q�o���fY�_��`�����z�:�-�S�B0N�0�&��{n�	���c�娀$�ךx��0��g8%ض�E���D�8�{ّ���VG5�(� C	:L���/i���L;�����U&obt\��箌7��	��Hr%C[�4I;y���6��1ҡ�����u���DΏ���S�z~"�h;{-�w$�,���4�[�'��sq��A�aR��jh��_��Dy:x�ē������~&
&>R���%鑏��wE��R1�*+< �-m��0�sB�]!yL4����;-�g�@I^��z���;�R'��M�J���;|��Ѿ>-�:a�c��!��k���*�fK5L�N��3C�.�����6J��_�!gãϧ���Kz�=< �.U
d�g�yI�SBM�����;�tя�#
�l��&�q�U=nbĖ�wbY�˼ղ�?ɾ��On�?Q�Ar��E����o)n�"�!���P�s�ߟ�r��,�f��s$��>P�����:z�_�'؏���՞C���m�81�h_���<���^�htc.�|���\*DBY���#Ji��,m��Ъ);��#��+�ʣ(c	�� 2Jr,���s�(Im�×��oT�E�-.���G�)� 혿�e�$<�x��$S�ٝ��j�� ݼ��݌�<�*�'�Z��t',����J�6ܖ�:%.�P����!d�rD6���Ě�q��Ĭ��9k&�����R�����Y��<�^S';�گRv:���>�I5�"�Adj�W�o>l�Ռ���%�V���k��h(��@4�C�H�H^�j=��
�y�)ٟ:����%;�\(�����1�<���{ջ-�E��������{��@X�I��~���Z�,Ap�m��(@/�&9J��衽/d���������j_�?�ɜ���;^:������2e�zh)4(�(�J�.�R�+�c[������̞@О��з�,��姞���r<ø̚ �JB�R�q�p��wAc���e�|H���O�����օL���0�H"�xcq�G�Z���X��Us���i�K'�>����1\�]DO�u�h%YS�
F��W��=��`�d�s_���~jgcZ�vpHъ[�?U�R��7� Hsh����R�~a��
�Ғ7q�X��wn��,c�Vg����Շ�^8
����I`S[��c�ӝ0E�J#�81rd�gƎ��bp5,94/�/)qI�\�" h^�8��U��{�[W�"�y�Q�e�6�7��8%� �2Q.�[C� *x�x	F�Ǣ��t�iw3WL���:#��pѬ9�S?B
��¾��t8%n�,=�Z$��&4J�p��-���S�ܠ�����j����,C��G�g�n�k��y?��,�hͬɋ�»���۔ #b�9���jN§FƗ���0w~C��~%��D��+j_���3U
�Am����Ʌ>��|/ �!�Oj����x��T�X�&tN�ΉM,�M��W��BoXu��4ֈ!L�s���� �XxPV�M�v¶�p��I����Y�Q �k~��`���M ��.�<Z�Q�q�p�\C$G���n�8���'��!�1�C�̼�H�Z��9��8!�5oAD��'0p����i���R�݋����"��?����X��L�'������Bl�/���m�N��C=�<���{�9�u{���l�vy��[�|��!�� �ЎΞ���K���ʞ�n5:�X��� wy�H�}9#����a��_��#�� �GO��1�.�r*���u��䩽S��ՠ�[
����t;Ap3�Y�H��8� �>�Ȁ_���yN���&9��G�f�'�E��kY�m�hzv1�6{�uP�F�~K�^�Vα���Vz�ƟB0���n|���ꎑ�X�^Z7ҽ(r/�9�N�������S��}Cӣ��+ks���f��:�\���+9Ri{B��w	�8	.1�C�#Yv�T�P��9�;��VM1�j�IO��m�����+4AP�Q��n�������#v�A��xg�b>��vp�M�Xk����Y��1�IBX���W�Ez|�@V��c� ������f�k�N 0� W����s%C9�s�����+�G����%�Q�@P_��=��
.��Ȗ�L���������X}����Ý�'�rs��+%In��lu���c�'��Sn��	�L^�ĉ'n�k��Qn�L_�l���m���u������b���̇��[��nK���D��kP��7P��3=�ӔG6��g�=���ҩ��1���ֽȌ:�@�O�·�I.^����C����X���EA. �(Z'7�fI���Ҭ������΁� R��lFB}4��j��J�g ��{�].�
����^h��c �6��2��.��4�&�/QF���~�����^�s��{��U�x��dJ^t��F@�Щ�#�e�AT�ɋI'�ձ$~�[5w�3��x`5(8^A�`Aj� k4q~�T�t�]l�ȝ啞�S�Rh����{MK�K �����:��\6g�X��=���)9�F_/�;�~P��f&2��A�g�+���a v��Ɓ;�(t7��Eg�ߖ������r�π�	v܇V�H�B��#��|��E���Jq�H�~��/m�|IH%�H�@mSL��ۡ;���:�����:���OO�r�c>"m[c5]�Ϊ~j���x5��no���F�(trً&��["������E%oG��:�5_ώ4_�̍Tˌ�����HƳr4����s�K�I�j|&�����\-H3w�P`�$�dh�6tɾ$�ք1�)8��t�6"��k�M�]�o M�d|L��_�.�Xm�`i��/q�B_�
q���������|I����=�q��3��ӹwkW����,8)�}J��>�_g�8�3�ؾAv�N��'�w���B�8P���߮�q���q.�I�������!	7+}�i�A?��V_C��g퍂��Qu��F88���ou|x5�������%~87r�o��b�7Q���i*[7&���ܕ���#DK8_���RX�Y�Cz�Ω2�;�����
DD	Ä�w��N�$� ��72e���%�0�u�8y:G��L��?M
�4���Vr�
4�1NB+��G��-�<�73-7r�he����q1��l�&G�lw�&����!��A�<pʙ�s��5�U� m�yQw�CA`7xo���7�S���Y K��5<��K��'�hJŤ���je������in�q,�N�2/2�ώ0y��y�S7UT�H�)�+��*���{O��?� o2���j���r���i?o۶���� ������Q��:�T�����%�"�G4��>����"������<���E]�V�|'�gF�,fGߟ��|�`W��X��c�.�Nk��#�,���۫���A_�0:ڔѓL�|�eV��s�8 �HC*>pC�y���ևj��倣퐃b6�X.#}�Y�����	t�4e�FW�#�/j��H�W�g������((�:\$�1g�S�����ֵ �Ϗ6Op(�VI1�H�'n�j�TFz���N*F9LZn�Q�(�@�(����$-�e8�R�~y�2�W��h��6���<2t������d����N]�me�?���e��
o���`���qBt��E�fj�S"H��<����5��l(��J�'�<;�I/�	�NK�"�?�l�����K^�������	?(�{��:ԡXn/�Sfy�ˏ��h
0-���dȰN��&���-:_�c��7tMh>㲢�v�!\s4u�ډ9;�>����%��`�_��̪��4�_�O��a����p'M�s�éOg�����N�7�P�Q?y���!qG�&	�/�����z����hN8y,�#���9����Gt�A�ȹ�b�P��e�~c����I6m8}<�
o�0g��H@i0� -gҎ�ؤ�l	C��e�����`	��q�j�@2�;���e�&�����|UNf�ܱ�c��p5)r)ඒx��~TbU��n ��N�MF`B�x����ǈ7�@�U���KiZ�q�F����^Zh_�[�|�`b�Σ�tp=���ϟ���N�����><ED��_��F�'c�R
��v�=��H�וD��ܖj~3#`\�`4�S[^�%ѝ��p���p���wʮ`��t�Wߍa��P3�v#�	Wa�����qR��!ѭ<����|:��ݼ������������f�ܽp��Px��P2iE�ٹ#��)�}ܼ����u��6u����@���y�s�~�e�E�/��T���J]��x��O 1�����.�d�|?��:����1��CfGq�X�Dp����['f��������_t_�*X�0H=y�'5�{�:S�m/��|��}�����B8���,�d�m,�ڀ��>k{�<�O���k����@1*�t�*Z8��
�`�/�	��8�0���R���?��2���۠�b�3N]�64��2��(��[�i=��n���(|L��l�*:�-]�ĪhO{�fؓǉB*6LW~��c�b�� �Y���<ՙi~�W=�O��|�Hg�Ƶ)��Ӊ`���g�L�#����S�j�V�Q���eZ$[j����@)Z��@�&v�;�'�fo���&=���	N+I���)^�q��� ��l�m}cĹ���C����8ӃW��fhsRG<_�pk�y�z��<<�d�,��qM���q�$&�H�DНRy��0���2��L�.Z4��� ��&��`5 :IK63�мVmQh5��gx?����g,��)�@SFf���!����C�D�n�M\y'
DQ`n2���b-����r�����ӕ(q����b@8��:��9v�'<L�`\@��b4Pл�\�`�%xJ&o����"]��g>;�a�p�E��"�&���:�>��7��
�'#P<�X�	���,R�*Tp�-Dr���hc����8�
�-������P4� @�q,���� �����γ
`�����
�W��f�sg��Ks�F��˘haL�(�;�[[mwk<�F�bf�y�ar0/&��4Q��;��x��۲p�`X�m�%#��G���3�R�F��?}�@\�y}��x$u����P��2]��v���(�9�Sa��ɯ�3�	OJ��푹W�(�+����x-K�3v��{��=c;�1T�R}�w�(˓�D$�weE�)g8P�:�Nk>�y�׊+�v���{��1*�n�	?�_W;�\w�筊q��+_����߫�����T���r��"��f���.0�i ^�J&�����8R�K�E�T������2��F=�(@FF���~3���;D����	K]��^uD�����r�`�|�r�nD�yd��bmoQ�}�� c o��n�|������ ���{6O�8�o2����w�H���LԀU]�m��2V����ŗ��c���SM���G\ط3��
e#�r۲�Fk��l��#����z-��C�E8�bYp]B�ע�f�@UG�N,D�GJ��68���xP���I]�Z�y˾���`�$��n��C�����W�}T�˄���a�ƤL�����l�O!|b�ϓ^4Mϧs@K�h�<��\J,�kZ%�<�{4��fjDG4����?N�d��=���r�'��<�Z��P�鵂ԧ�=6�.��pc�|QJ'�� 5E®׆5 mގ�.hH�τ�¢ߤ ��+F�E�nW3�q��٩�6��R�5Y(�1س��qN�����`�2��s���`@��lV�d�H�~'��\���č��j��tӃ.�3+�������FW�����T�Sցz����<yΡ�t�n�v�b��s��1+c�%�i$ 7��=僂$�;�e�0�jn���0�"�b����S�hW}v�]ֈQ���9�:cIO��]��0{�Q�ލ�L��j��" �\r���u���|`��GֺN���%Gm�nJ�xV5_���P���x���J�H�EQ
�;�$9=�ש���+?���kP*��_���H��\�P������q�W�-r2n�����P�n94�7 �r�g���0�I���[�T�v#����֟����"$�`ڣ� ���`�|Me?F���϶�<1#Xga�%��@ۗ�5�%u��o�b�w��e<:��B�I�ζ��H㏖�xg)�s:Viw�ς(FqX;b�C�/-� �����.�Lnay+T���L��� �U����.߳�v������8��R�:��{~q�j��ϴŢE��vĆ�:�I�����+�S0��`�!��u~�yv���+�Bx�ͤ$;�ܷ��D�7�pɴ��)�i�w�h�c.�$��}"5�9�KT���N |��󜼙T�����!�4u���_������*�R�7����+���]�"�J�n��9Q�,�Q>�˝��XkJf����iY��RPc��Y�B=�X�__r����D��1q����	�Q����R+���G���X1�U�[���`6d�'A�n����v��Ɛ��lk1d�4ݍF	Kג�����c�X�!�����]l T�<�� D H����CT��)��>����\��!��9ť�XT1����_�ү��=�sN`+�0m�x�y�r�!���R@��_���x�`��r� (w��*��=�O����ao�48AO�9�B$���$�n凸�\��;�:NH�&��Ul�w��,�'�r���I|�_-�dD�so�h�	/�$T��b������s�t��"t3&(��3���4Cx���eK~?�[�p��sl�����`W�I�mU7]OAA7��������$wdy����n�� ����ב3���Y�*Ff>��/�Ӎ,����-��?*����^��@� d|6�F�Z�l `q�F!%��?��7�<���K�"��Z�0<�)ti��J{)3�=�,N;qZ�;��x�tCk&�1R�4�sS	�R���V�E_%�lC�CVF��32��,��?6Fj�e����D�7����{v����S�=���H|b[��e���[�z����K=���﷛0[ ��Wc�Ue3Gʏ���P�|4��Y��FT��(Қ�=h������f@G�s�b�� 	���T�>'ܧt+�F,I���$RjQs���p�<Y�R9��K�,pHA��{p��
)�\����ν�Z	t����+ͷ��2j5���X����|�<RB��D{w��~]��dV:H1�~�]m�Q��ջ=hw��<��@�3�L�5*fS�|�J�ǡ����]���4oG?��)�];�$�
=5����	���P�be�m��k�2:&��ç��Z��oB���x1�ڈT�JD�F�M��یλCb5|d�hM(�{��[R�������l��8)HC	�N�Ą�&��%���A��!�T,?��Y�gj��� cϺ(Yq�ʊ�Tx�Ϗ�bL�����e�;��ij��{��/�09.�ӹ/��q�-~_���#��G�P_XH�Ė�{���	�H+��������i��)���3vw�#�ќ6M�X�u.�z��?�E�����9~1�h�������X�k�}�e>��#�ʞ�6�c�t��V�lFO,,�w�<����V"8���\g_sI�T���4�.t���Y03�<���~�2@:����i�@�cQ����_�E���"��[�k�oDH�ǫ`4��D1��LG$κ^���M�L�c}�F���Պb�h[Q��U��jmCq/��͸Kep��t(��y�Id��D#�f�/�Z7�����`*��,:k��5��L9n3�-8��!V��lusS`��I?7u�/��6GXm��qf��ΏF�L@����\)�9\��PgM�tԩ� Y�R�����4(��s��������#.�s�����
�#ݍ..�;:�����9ɪk�� K���>lA��&5�sdt3��X[%�Ob��4�ߴ	?��L	��A�9�����I`�9���u��Bzx��S�I�8)%���YN2�<�Iu��Jo
X,⪓l��q��l�\���KPc<�T�C��2��g�����X�Aq*�f�����\���R��z_`:��9EnZ5��0���Ӄ��=���)նa�p�Ն���D�l���Ϛ<�$R�o�.BG�v}��Y�oj��9F<+�����iS'�f+R�a���^����"��|��]̐��|�e�E)�f��},(0r��=Lrn!x$(E�y��'I�S��&u�U�98ŧ�(��P���&
��-���Y�3�gɠ���ځ(���H��V��E�͕kiݸ��pӦ38|Q� �`'F;�IQ^�����8��ʆ?|ڞ |��YS{kT�},�ً;޹��A��bU��j����f/��;�V`��2�Q���,��[�k�s^㠉�!�Z�$�0� "|oe�4#��&������T◇_C�R��O��Sa�Q�em�xo���ivtz��I֎_4��d�S���4%���Ҧ�}W�o��R�	G���_[�nWLv0'��{=�qe ۘhȵ��DO/��/B�M �l�c�m]�MiĿ��Kuw�>��ɍ��z���ܛa/��
]izW�hXAf���q�k߸�9�m�Ƙ�i�v���p\�V��'��4>S)b��sǁ*7H�h$�6�Vq���wY��&� !	9o������Ǔ2�J�����My�_U=���c��^>��ظIBEP��3� A���4����Z��G�Gd,�b	�QHj�U/h���R�
�^�@�A˚��3�t9w�-ĴJ�*��ֹ�(R܀�?Λ�HJj��탦�<�=L�q9�@��V�� �?�5��ZLP0i�Òem��Ϝ��$?�%C��w-��ZR`4��f�1�N���D�܇�>%�dVp�;����hl2��ң�M;��L��xY�XFi�g�O���k� 'l9��%��$9nP�F;K�tobZ�~��QE(�`��B�dy׏���)4��1��b����J�nN������b�A�nq��P��6Y{���{
z�lEZ�}9h���z�$�gM���E���ޅ�	�)p&���<YGK%/������i���iD�}�`k5����N~Vy��DZտ�?o�����rT�3f�<*9V�3�s�Jf�Ծ*���b��j��u��N�I�qZ}a�r|���6s,v`�f,Z�=Wl�ґ��_�O��מ|'1��]���;�$�d�9�l��4c��*�*���PeG�Rgf7Fc/LE@0�+0���w�^N�G�|�����Ӹ���{94w<�g�Z�:wkh�v�]t��`w�x�z��<�XT��2�ܾ�?�6�`XNܹH��p<�lK�1�O���,�Hb�{�ζ�4��T��"&̂�HI�ÂdX���N��]dPc���"��{�]z���^���O�'�OK���4���	��(	uRlv��[�5���?�!nC����:�-A�Mj�BH��2�1�"�(z��7�����l�;.{�Vą�7S-�z�B��c!xp�#J��Sޙ���*�KY�"��Yk����(%���.�H�{al�ҫ�纃@���ߛ�=3SO)-��T�F�1R7.����J(J�2$�����XfےӌW����@s����`Y�<�}Eӽ,��1#�L!����Nf�/�%l��	������
h��"�ݧ��'t}@�8y�tY�>�����x��C����O�s��%�� {��!��x�G?��qV�0������rm���m{�G���������Qs��0�w�ck�h��*���`��NE���ٖ�D���0\X�p�:+����+1d���/�ғ�jw��?,�Ч�gՊ,������5ICk1�u�i�QQ�	o�^�����m��ES����|��oZ�E=��A�m�A��99/�Z)-w䣁Vt��3� ��X���4�W7pfYn��X)�����9������7�3�MIm>��� 2TvXH��25�_�^�ޓ}�N���d�]���yC_�[h���=H�����Ϡ�ƗE���;=Nw�����[��R��ݲ2%�X�
��A��B`_���.����[F�@fZ�N�Ѹ�!�
Fރ-[oŧ���	��`3;0�U�x�j�]H���V4�N���D��PR�&eR��\#�7����W�)*o��u��o�
z�ؾ�f집J�d���Z9���	�3W���P�e��D�G�t����%������u��_� V�]���E�ۖ�����0����}�AX�~�)�,���P���p0���a�{'���͙�L��v�Ɔ�+�èY���n���\,�P"��� 27A�?�e
��o����HuR��������pC,���w]�`P�?��h��A����hy%ۜ%��. f�5Į���鎗�T�h�eKF���UlU�_|��r��G	���p�+|��FԖ��n't���[�Q�ޜ��cY���]�O}D�����X89f�rFtp����c!��7]Ȕ�L}�}ŠR�D��+������S{Z,
����7��wj�F�*f8��A��_�)������Ht`x�#M�"	�SU��(��}R���n2B��M��e��FE��`��]�_��b"�V�TeΦ�>��n��Gp>����Q0���e�.ɥ�x��W!� !q��{���uĴ�_A�c�c-c��L��$����D�}��mA��P���N\"�kR�O7RPH�����2I��=5먥��g����/	�$ݭ�Ô�Vߴ���4R�����
�������yk�ɟ?�;z��[�����~pFʪ�ǋ�*ԫ���������@��],��V�	�jx����M?C��Q�ԅٱT�¾^�u��=�g�a�M Ň�<�,x��Nw�1�p���2z�5��^c���Jd�h|� @D�\)����(�4?1}�u�TI�^q��io��J�M��Q)�ޏ�����p:�Go����i1c���D�p�^eM���ҿ�$�jiП �ٓ�������I�����oұ"rόYT�4��
	:�@���#cՓ����H0��"!U�~��8_�k+	�ߟ�8$�l�C��yT��#�p}�LZ�E�`���t������ u��v"�"�_=٩����['�OZ�UmSC1�נx� ���+~���ౡg0����"��Q߯�'Q�A�zU..�^d�K�'6G�N�`Ԅ�����.�@E+E��
�p�
=6 ��۶�FФ����<���f]P�A��������,�WW����#��'�ν��l�~ �|	�:qZ����_,���c��I\��j�X�A6�_&�i��؇(u�ƨ�dvٶX��+J��_}D����6,"o��RM���ǡ���;;\>1Lqx�Z���+�6p9O�@׏)���%{��GD�EVj.���F�]e�1@N�d
D����(�6�ڗnq�S����~[��
��b~-bs�(n=
yxP	87�S��2�K&&���O��D1��Zt_�pRF>.����hY�@���}�;ɅY�`m�,�t~h���0�Fڞ��E�R��2R�&DX޽�;|�?�Ќ��0� �NO�}�V�� ���ӊ��u�WL��ף1ViU����J�8�M��]v�bG@M�]	����qO|�"Jl�I|�g��އ��p�˭s�G��:�2��R�����Fk�� �n���Mt��N�+�#�:��� @{��7�o�N�ty���G��w��L�� ������;Vޔᰂ�˱c�ޣF�c�8Wq�:/�D��_�z����Q�#��^����NJ��W�-�񠓦j^w�����JI�Y�IȪC$�������C��u�|Y�$#��:*���p#�Vz����F�!U��*������{�k��J�)�+A+e^�������*RE#�=�.Y�������T�Ѓ����|Trq.��r5�oB0@!D���F�$�5�����G�4JË���4�H;^:8of5��[�o�:���s���1�\����lI��:�v�ƆX&��q}hK�y�/jҖ��CʓZ�ߠ�Q�&'P2��B�P)���y�,G8�Z:5)HT��f-J"�=���ӧ�Cp�ޅ��{Li<;����y�L�ر��(����N1�)�a��^0F2ʖ�q��)�-t�Y��n�3�]�E��\�@/�ǋ�1r[�P�����z���[������cj
Ҡ�Y�E3�K���\�H٠-S\K�ߴ�B����p($4#��&�PA��@��sI�:gl-��u���ǨCwROL����L𐬞�y��_Ao�>`��1��ܭ�rn_Б�R��|�g�$��ݻ��W/�	��3��CT���r�ڵ�������F������vE�Y�U�e�1�I�`��pj2�oX5A�O9�K� ,P%C�#�/8^]X��?T29��nK�KEEJu��+O3�4ٗAc�2 H�:4�t:釋��~�ce�Mne4�	�.���
�>�r���@����F�<�!���P��>]����#�b��"~%���6�Hufu�%tƮ{ۚR{� �3-=����L9Q��3����[!J���/�H!���&�JǍ/z��;m�q}�ǯbI���R��a��� m�̄g6�d+%�xa����N1T�&�N��?�x���8buo|_�Hʀ���\��!1�y�hM@����)F}2(�z��){�ض�S�$	G1;��&MmUẗ�|Z�D��F��g&��fi����U��TM�����AiD�̥��i�q۶�'Z�;Z��Զ�*�#�y�69qp�=�lo|�W����O��m1L��f���U��z�do��m~9�\����!��o��cN�=�"���|�sUﴝ	�s|��g��Y'	\S��#���B��YJ�����e#�4���.'G�V�U�͎�|�<ձ�담Q�O������tf�ewj���sfuXR���w�L�7�a��Zʀ���S�i���~Mt�X�o��v��g��+�z@�")�����
^�E�����dR7�����ӜǙ���i/�4���.!p���O�Ƃ�j�j�ؒ"J��փ��_w:X�+�`�N#�����F��i���"B4��V����H��Y����F)I���d�k�dvFd�V�+�`dd.o]���N{�ڲ�@Gʺl}�����] ?�QJ��p����Y9%�۷�!$���[.H��X�9,�O� ��t7�M�� [��m2@'�C�*=*��ڥ�sb�`����(��v=B�:~�U��kr��Y�W�[ 3.4s�ja����+=�%������T���j�=2�}������2�+pk�D��(�?�h���KC���4��6�vu�Ў��e�Į�`�D}����s��#BD��%=��cZ�#և����\!���bD�*i�c�5��c��!�b�C���<[�FjJ3#��>ޖ�r�]q�ڛb��2���sr��Zx�6����O�+t�>Ar%��!�X/�۴���)oz�k�84��mJ����sNȻ��j{��X�B��6'і�<����*+�]��%�ȸ:�
��`��̪����dl͗SDD���Z�����2,�d¥����b
4O�Qˁc����)^̦���"�ҧch!�m��#���)���tP��`�a"R��Q������>쨺������'FN�^��R�IoY��M�@��;O ��;�\Ъr�bD�=.[��3�;�)��\Pet?NX�g`�	��h����I9�в�8�Y?�i���l͗@�� ������p�����=dS�v� t;��&0̔c5�FƎ��R�66Fs��:O
���$�}�INX<���/���ނ8�&mpB�=��|
��Tܽڤ((�����(3��n�"6hȗ�2�X�}�j���bUN�C�2�G����f�w��p�"L��Ky�|UŶ �|���2�䅘Չ�[wD����-�=:/�m� 5~u��M}7�Cԉ�i��n��������@3�n�4��(3���'�VS�1��Љ�"�>D���>��� �)��:�w@�<�IK�޴@8}A|h��@i٨r ��.q�E>�ZD$����h�Z���	�%0�~�D�Έ����0�[Yzb�j���*BǇ��ŀ1��7;GY^/&�[�in����>7��IG�%?��
�ف#���y�))�d�_��Mq(Ǯ��n���J`��'{T�����*��T��W�k�*1���M��h�N�7���i�~#}�((̓��\��>p��8!�c�ۼ1^�Pz����C��쾍�\]�TM�FD�ԤVO���~�K�3��_`����`�#������Ⱥ^*ͫHN-�=�.J�?)�?�s���������8�X�zhy��A��݈�2m*��z�s!��2h������|�0,z�|m������RJߵׇ��{+��ȵ�(�<v�;��[x]��e����ԕ2A{
�;�
,s�OJ�OH��Tl�����Lm��(�RDP�a��$=���(=�R�r��n��~�2ѩ\�s�PeJnW���.90�w��U��D����C�9�V~��,K�;���]�n�"aW�D�Y�{�ν�)"lj���@}m+,Z ݁���k4�i�K�(SNK��e�ꙍ#�\���(tQ�N
�sO��x� �v��(�u��.a����ز�ʟ��z�y;ޑ�)v��[L�hh\f%�>�~��.��+k�x�h�[ZƝе�/��စu\.�4s��-9|���3l��
M�O+�(������K�:�mG5רn��)UL�"i�cw{}�3:	9�B���K��-0�*$�)�{p&��I3�v)���g� ���:���A7��`�2�W����ZI���V��y���GRM��C���7�����82n���S��i;��`�����kp�B[t�m���)縧|y��C�Jn��"�O�T�RnéI���s95�ʌ#��0�r-?���a���6��������L�ȤVaVQ�O�n�v \ϛ	�X@�a>Q6�ݓ�N�@RP��%sM�vϠ%T�w_]nr��L�{7���uL�e������A���&j�8mcݴK{�wkK�p,��L��5��Q%���J�>=�<�:�B��3vg��V'���� ^��ʾH ��ܣ�g��p�x��q�r��F�� o�aEg��ꃌ��m�|�V�I�D���L����<_��,��>w6����Ox��Z�G��x'�Z9�7�X�ҰWT-�h	�.��DiI3B{{�2=��R��]oɀ�9�\Z������ԅ-"�f�+�M�0d࢒f�<���ES��`F%�l�<��?%.���n��A�c�S
��"�ړ��2�n�'�Տ�N@W}�]�L>�$��`�=��=h7�{���v���*��M�̅�g�r�X�?�J$%ظ�N��Hm�f��3��"�ip@xG�7ѽŸ����t�8�\��s>���E�a���vW�~��@Ɂ�>b;8>���TO�dv7�1�	)8�K�q���!�ΖsB:{^���09W:+rH����ČkD�u�Ѳ��F�9�u���6>_�T��#K�}�;������	�E�wJN����gG��B�XӨ�٠�b6(ttcۏɞŬ:	���#'A�֛q�b(���#����h���;t�eV� �]���be�E+$�4p��Z��6b:6���H���u�t����{<�ax��~�ږD�n=[�kI;��)�w���K����A���5���Y�/��*����kPvd�G����#��@�C�1;;����A �"^��3�c��l��/!��h��;���j?,%�3��oM��]�>����kqq�!�ay,C����	N�I��B￬�� ����@�
�NM7��c;h������NrX��J��� �����xX��54#�m�nѫe��ƃ�˳}�w�$�� ��a�����Tq$���*��R8���nڭ�XȦIe�eF�kvŞ�D�:녅��@��]
M��^E5���m�m�%��9j�0����A��R��C4���b	�/�K'5ht$���!�J;@�$1^��eF�l�-��)l�^��^�i�0:�RS�(�Uw.|y
��WG��x�+�g%����LGǴZ:�U.�y��(�4����\�2)j(��P	� C�(˟����:b��^�fq�d7�.��y��R_��g��K"|f������m|섋�o��҂��o~�{�r���(�6k�-m3�E��4�{�e.�����,�[&�E�NA
��ԩ�F���ĞߗI=�ٳ��I��N�Lֳ����j9u� ��T�q��J@�v#xd��*�rِx�"KC�TH'���f�IE�6(`;佺��S\z�8=u�L�̹�n~��l�Wd�8�5�4�����;�S���?}��v�� x�z`B�@=�T�!k��{k�yڠ}̄/�IWbr~Z���kFK7��<����-�S�Z����i(��_����ږ�w9�����L���N��&�yɘ��IlB�w3U_!��/�������\�4DG4����%��;c,�	�v�-�a=Я,[�8�g�Bq�hf��p=*��O�R����}g��f6����u���Xt~����mm%dr����Q@�Z.��"��K��Eٺ��P@Q!̵T��	��yS�)�C��:"�ix�<�]U8�;�E]�<��,�u#�~�c"��yW�,��/����5�$z3����|�$�t"5�Y�����I��_���{5��4�2��r]�	�=��(+��u��Ζ�}��H�&;=�&^� s0��.���co�s��"~R*gԶw��%G�k^�(>���.��7��3�|�EA���m����^��m��si�n�����Վن}3�������"����Rv����<q@G�����۬{T�h�Q�=��|�o��D�����6/���(��z���꠲G�R:��w�.`G�%�MzG�!;ӎ�+��2̓�i�����gS+��t�����8 ���1��Z�� C�iGE����E<�
Ji�YR6���}�\n|�8�~K{�^ZL�����epPH�iȞr̍4&T�Ц���
��=IR^c��P5^V#�خ��`|�O��;R�e�F����AͬAt���"7�b�z�L^A�{@��o�+Rr���̩�H%�e GM�`�E?��aI��@s��[���3bk�����aZa���A2]�&�6M�wʔ��9���B������n���'�K�����}��]n/��Yk�+��9zX���6���pҸ!Uq0�' Q�!������=�U��_�s��p<��+�����#�r�i����3,`�0m�K*��x����ZN&�Txإ9�����~S��ҭVfB�/�KWi�',Q�M��jI���9��!K���_�U�z�
_�P�J�AJ��o��:7�M*0sĶ�~8#��bL�s�M"�/*����L	��tHHy��M��o���l��hhV��D��AX�H6dG@Q�ͷ��c�������R6c��h��5��H��~>�Z�{s�E�D�W���!6��wU?��8>U�R�B8��vژ����y��~h3�<N�D�v.yz��I�͎����d~�:��{��+.6���F&�����5���7W�H&	�P�N�|Pq���&U<p���f�!#_�l���P��i�c�)�k��!�46|�����޹-+�صi2��V�[z��8z�^�$��VӤvG�������]܇��$5���K$%h��Ċ��~���gҿ3)�[{�B`z�Di��Q�*���z0���_QE�; *��j���P_��̳&��#D�`��p������|�+� ����[Ư3"��Ɉ��G�Whɬf��C��V��`頳~��TN3�Cٓ���`��"A���Z=IG�1:�R[|�T��6^$lZX1Ԉ=����ꅌF~Ff惐�>�z�1 �a�2�.�������T���ōV	�x��R/�g��5�U�3Γ)�>�ks��� ��
�B.��߱��&᳝e��o�������$Jۃ�{!�)�U�ol<,L�6�	~���j�����v6�9��y�������6¹�R:�N���^��f��b[>��#
��Cʁ�~f}(��&�2�X/g�,Ύ�� "�+p��`f�v��m�K��\F���4�"�,o��V�:�^�C��'B=�<��)eLy�c�L����n\���K�2l�. ܉o�W�)�$�b�ţ:ݩj�,��?6EZr�ݑ�HI�s)����^��mޠ1U��"ߤ+1�_���*�-]	��x ߸�>�"�ٔ-@d����K�d��TǕBۍ����*��e�����|����=Y�"����	-̅ų纑s	T�)"�	�I0]��^�w���av��xf�,�9��/D�N��{D|�ή�����(N圭�S�Aj'�ܾ��U�c�v~V>�s��7�fF�e������
�b���t�X�x��d�ץ#���5�]R��jLEd�*�i�3�A(W�[@k��gE�׉��=��ә<J��R�	m�O����K�̂�++f~��L��5|�x��ލ(�2�c
Y��B�O+��V=QB'��$B�����Ӄ;<�W�'{�� ���ى�1cI�螄;�d�;�9j|������^���~N����k4y���k�ox���ͺ�Ԇ�F+�J�%��K3S����Îۭw5�ꁴ,�xH���lvX�|t%��tcռU8���,�J�̠�l����! W�	UYZ���j�=/���[y�`�������Wޱ�87�I���������Y-2��&�9:��
�U�3�`�_�vn���j�:?��S�)a��W>��Z5W�K9̄޴I�%s��5G,��B#l�5}�bsi��d�a��߁(Ԉ������?�e�3E??[��[�,_��C%���t,��zv=�As�D��8����|ûw�Ns&�:'��Q?��W��m/8�1��w�o���
)�b���	��e�D�,K��@�4w�,�c^]ȍ�Y^
���1Ȃ��o���B��t!���/6#���8E�(���������� �Z3.
9I|�r�Z����s�K5ڇռe�ѯk�+/�%� 3�Ӭ�滁����D�j]�����͠A�@�/��d0�kd7�0M#���Ğ:����£��ZLD�r�%���a~��t���k~���rF�k�x����>e��ћoCj5�\�6Neu�Η�I�H�"��W�š�c�)?YgѼ�iD�Y�cd*ֽ�}7,�O��0%�!Q�6��[{�Z�:xZ��){ Z�4Q�{�]Bv+!?a7S!�Z!	7,���&b��6<��e>�������*5�c:% �^Au>u.U���f��:��9~e�i�m�8��_R�jgx6�BP�Z�d�>�b33�U4����S�~�l��0�{��o�o�P��6,�����\GV��Z���(�3���!I�e�ه���;���+�պ\&|ᰎׄs��U�FAۃ���!����N'8_pFx���#�Ѷ?�M�[ټ��?L�V���9�z���{�2��8���$:�G��K9o�=�}�*�a�����Q�F�1r�BR�����c��$�F�kn�8|���/���u������#8ҿ-��
m�C��Ixu�bGjx�:� ���I����i�O �c� ɷ�Jh�G�|��R�Y�{{��XpE$�����w��*2��{V����}%_�M����U�Ѓ�h&	u�K��N��f���6���ڏ"�R�'�,��+7�1,��i�(�9*tp��������Ѻ�*ozeS���5AumPGo*��o��#p�	�Ew;~ې�.�#�5��r4�q9��@zVCq�&Pe\1�k ��ڿ��P6mxm ���r_��X��
��X���g�)���hU�P|��=�_X�}����N��EK��=��L��u��/� ���E{���/b��5*=%�μ!�b���+F&�?%|ؗ5 5�D$|����'X����/OٽO9N�Y��.4�bu�q�K��Ћ(o@F�˦�B�����SĦ�d���@��M��K�K��i\6b��B���F瓼�F[��	����";)��ZV��Zq�N� ��cEw�&!��C��DZ�K2i>�{��.�z�Y�OX%��΄�M�H�R0I��$p��4���`���9�]�� .�F�ңʁm�L��Upʪ�`M�ֽ%xw^��zA�����η��}f��E���_s�G��g-�Cg�, Z�K���<���r/���{��B�H������	�Q��W܊������,�w�go{"Q����ޥDgg7��Ҁ��!���[�ښ�l��:�3B�ݔ3�sY�%�y��x8�vVj�vzBr��`�g�H��J��y��c�c�&�4w9���a�z���_D�o�K��.`鍜\h�GP��V#E��#Ώ����B�64N�rd�l�oNq,�ԉ��T�{���|�f$؞��� �4��$�-�6;����%x��V2	��j6]"S��	jY��ߢ��L&�
���O{%G2<�m_~3_E�i햮IQ�krj�/�i���S�:�9���8�y�C�تN=>��=���(I�0�e}�9U\��w1���o0����P�s꿑M��Ay��4��ϑ+t1í�(��B�J7���g���2�ڇ���f0��㛝�t�w3�� ���A��H�_6&ָ�J\�_����m��(e�GԤ�L����):��lPm&~�P3�X��3����!����B�Z{�}V�!5*�<Oc��!b��ƠF�8�=}!b8��>���1+�K洔�5�5�wx��q���O��R���Ȯ�4.��e%aw[�(��>���5"��\	c�v�Iu���s�y�S�أ�G���?�������K�y_g�ޒ憐odb���ѥ�x�p �.(��㔲���?���vW+���_hV��¦ާ�T���I��^�P���˷+F��w�\j*�Ն����b�Pc�:���a�����VR�4p�4��B��m;��7��$����7����=A�t�ir:�-�!�Mx��
q*R��JU�K� �b�p��YSf����=����q��Pr�j놓�i����� �u�va�UXM%p%���w����ʭ�k��E����V�xt4��!c�u��g�K�$S9�}\*�V�{F���Y�ܑ���Ɗ&�٦����[H#Rq+��z�@���n@����"DJ:Z�ᕪ2T���������v�Am��~+`}�9�k����~O��	�y2� �O~�M���N��L�b)��a\�)Ƨk���:���⭼g���8
n��E\�w�ސ�ҕ���-{�򛮽ә�m�	������%l�CL�y!�=�o���K�ޒ���;�y��O"���A��huS��&J{aχ��HB*U3�����B��L7<�w;��lN���k�ͯ����"�xy���-�F�S��u��&Z;�D܆�
[��SR�{�~驡K�����PV�W*��;��HRmc�q�ާO�0	q�	Ķ&N���SV?v��*+��(���_Zs�{&���.L��5Z��N{�)�7�������|;U��Br.e��f��w;��f��~�?�.wVu �P���C�1�Z��_N�Qkxf�@�U㙳��t������{y�L�5?���oC�y>Ǔ*;;��fr��\��w�
�?��|�)P�]dN�@��y{5Z�8�_sӵ��z��v;���,�L[DB����D[�-V�`��rVO���g�YG8,�L��\�-�����F-�଻���-2OoW��*ԙ���}�� qb�M� Ȓ:~�H2�;6/)x���x�����툀�Y��r �,��%g��k`L5i4!�*�(C��M#�rz�fwC��u�r�>���C�hVT\�ѩ`�������:�׹���b���_�k����u���suz�u��%*�x	`l=C�q�f��n:	L����h���Ň��:�u��|���v�����B.���.������BoC _! ��� �ݸ�[�$3#��%��L���kSI�uD^KaS/{���&�g�Iu�4hkݓHG☦�Y�-!&�F.\�+6��ލ����� ���L�YQ�� �`t�����b�4�[�;��-͕W��[B�|��vc	R.i�C�K�IΦ�fpOY�b�65	� #��b����j�r�33$�#���p*�4`Chb����'���+-~�2"�����n\�`*Rꊼx���渔��6}�����j��+�8d���NV�ӆv�ؔ��jD���@t���m�c��O+�b�#sڈ�RZ�gIr�KZ�n#q�����}�E���8lZ=
׼��=o}[�𭀈�{�'�����Z���x�=���A ���OX��i��w��D1���;�o�o�	����~��%����{��@���prS�^�'>�����g�	�#a�8�u�I9�t�;�j5А_Vn���X��[��9DGtڤ�%#��;�o��d���g�"zQ�Ec3�0���i���Bh\U��k�B�zޤ�#�r皀@���m&�C�,����dz(��椟�u'�Wd>&�K1�����A��w�2�����5
���`�؋$�n���_��?�,�6���T8�Mu�r.&�Z��f��^Ğa�q_.��K_�1�(�A�K)��$�Mw�(�sD��}������3r�h��6m�����/@�T~b7�C}!��i��=.!�c	��ᐝY`+���V�Ե9C��mV�Ɠm��iҫ#�d~sf�ߨ[�I|_�m����;�Wu���ohl;���a^[������3.opu��
@�:����}�]W�|��=�9������c`�G�&G76���(��OD���pJ�ųO���/�L	9+����_�Qҹ'�׃��t�çH䔕gb�y#�f�&���ST�'~$��AY�k�m����[M�����|�cgO�}�@4${_4=�$ ֒�\~}�$:��T����f�'��aC�9�M����Z����Wt;���e�M�B�]f�L�X$b������A�f�e�s�������[��'���������$��VQm��|��C,�~,�*��ŵbOI��˷���᦭�cl)���F:t��
l�#�v�y���c$,��Y���6A�ׇ��[T��.`����%)ӎ�� r���Ի�� ��)/�����l��t>��O�B���ZZ{�1~"u��8�&~�*�}S�c^���Pr�|��!���1�K���-|	��f(�ɇq����a�к�V�7N�}��c�������v
�z��(�_���c��K��d��bS�A�m�cMM#A0[p0��b�3�W����4.�3^ʜ���6Qm�>-�<WM���úk �Ò	%9�T����Sh����=��%ͦ�1uŉ3�����O��"Z��HR&h���p��N�2��ꏢ�q���z0�����*�;�
y�Z>�a�1�1+^���8����\pd�V��b�.�j�@V�L�˧ή��J�ԧ˦g����'?� �Gv�y�;���%8���E�M�T��RpM��L�^j���(^^���`�=��O��&���q�=��nK3�mv�l�&U�	����U	��q^���VrS<:@���B�/��ĳ���	X"搄�"qM��g��ݮ�`-:Yw0x��ulx�x��;�2B�F�f/�J���Znc�e��>��d��QW���ǭ���LЩ��5I
j��)`O�.S�������� �<��ni�&<&�#S.���T[�0t?��QN9�]��D���>�^Z������Y�d���h�Q:l��-�Ԍ'a;K<�,��n��{�yW_Qlq%�d���d�`ߒ 6�ǟ5J�����f�p��P9������w�0$�	�2��{�,C+�	�������K�� F��!�;Gt9�.`A
�r��#�y�{t������,���4�@����B�*��k�Q!� �o��Py��!P�Aި5�V$[k��mίJ>�M�>�n�R�\�t�v*g�dJ#CYq7�܏ʊ�2����v���I9�>^�����P�BzÓX
����{�������ߚ��s�O�aC\ϭ)��e�+���c�w2?���:���s�D�#f������}��0ml?禢��-V����e���G�[���">\H�*���M�U�Y�[��YYzؑ}���ėbo٧^�2$H�+5Ւ+�/�czl�	�e�i
,qL��Y�C7'�G�����_D�0��k�%�n���'�ېV�D-O253mi9-�B���ɿ؁�����EȻ{g�K����,$r�NXH�{��nB���\�-���A�C���c��le5F���ϗn�aB���O6���D�������/*[.��?Ӌ�y��,0��,AcS��+�4=KG?�u�_�up�i꽹�	�̒���ZP����tS�N5{�q��>P�X��t��6��Js�O?��a}2�n4����Z�w��p�e<��Z���zZ�wϧ��̳FG������$8QCZ��M�QA���tf?�n���b��t�
��y��%�%jM46�A�5�oV���3���	]�	>u����>RS�U�����n�|	B�Ghs�gr��g;�QgJ" vX�E�t~�ʵ,�/ukpI�Vv7�p;�/p�����ɥye��4� �?�������3K���������CV '�֛�4�4��(r�w.Y�i���t�02��7\��Eы:,rk�2��L2\���Ȁo�3������EHU�y���3���>�����VƱv��C�R�lW(Ȕ0s�:��+��^��"��T��&E����`���Y3R�7Ɓ������{�E�j
/���:�ƕ|1��T/.�沠��'w�`)`��P/����3��捄׫��eTl�3�gM�9 ��;�Fh7�0Ϡ�d�!GS8���`]s�'KQ�3ޮ��NN���I�>�_��E-h�RN3��l)���j�BLA@������d	��u�(C,�>�ht�*���4�Ufv�Rӡ�|P`7u�SU����f�n�l���2�)8~Y��L�2\w+{��4|� b����ƠI�Q7����Ĩማf��D;��:��Q��ma��HeӲ�g�th�z�z�lԩ̡�W���MD��<�h+:o$ �?�6�{���m
F/GD�Y����j�k��W
Aׅq"bSa{�F���D
f%�ڻݹ�-2���z�ѝV�`�u�O�u??Fg5�4��/e��\ �j���S
�q,v7+ߔr�Y�{
v.P������HM�Ry~>
�)���HSE��U���jw�f�"���Ԭ��h�����!�^	9��O�<l�A�� �0;S�%�v�~>�OժU�;�B?r:[S"%Ќ�`5�$�o��,�"�{�L��4��5��6@�/���m���"�vO�������{�Cd��v��	���H�d�9@���ȋ��G58�B�s���~�E�?�%�5)�\��nXlEYi�~��,���ꦕ<�����P7^�nPo��(Tt��\ׯ�Bzߦg�6�W���'ɦ��OpL� �%TB�c	��
$�V��r� �K{S��%BP]�&��$Ǯ"H��ğ��n{Q�.;���Ճ��y$�BF�Y2��o'ڱ��֠�7�GL��b���Z���&v���]�����ڍ|N�C՘z��*�r��c��N����5ǅ:O�ጃ[�I�<j�mx�C�v��s-�����l�K���)G�=�l-Z�y��I|���~�Df���{?0&:?��co~�`�uX�ೀ_��5]���j�3>�i+ͳ�~�)i��p��F����v���M�8�&��b�h�N%*����Hl[%��c(����>Oc�
�{��T��2�zT��dm��l�ֻ5��4�@�����u�[�A|M �l��\����}k����A�ƅƐ�I�L?,*H��� ��g��z:�N	r-�%μ����n���UZ�~V�~X��o����/^q ]���ڠ[��<߅ ^߅j)T���?�`(<�U��ڡ�m<���%��3����-x5N�{�V�8h�[/6u�����4^�`!�oe.��r�#չ���K�U���.� ZO؃���fQ�0����Cq�'��!
��v�g��&2lrs��\���?I2���[&8N��(�Z�wh�@��!�AD�
�ql5�o���0�g:e �a��Ok��������1�0:p3�{G~_�냨G��j-���V+E̤�A��^��?�awP� 0ն�GkW�����=�叽��8�(|�s����rdc����%��P_��
b����՝��Dzqrp_�Q���g�.�ت,�h�_e5��~�ZssI�tV�����x��l�<QG�v�(�)X:v5P���[�F]���c%�	ѷ��P�eaZ�J)�T�1q�EC�|6�0��{kO&�l���̧܇|�� �7�9�|�. ��ԍU^]�&���dI�ع�=JXS�/�'{��kJN=�)��:��ӣ]�9���9dHF��c�Ci�g���E��,	�I�+�y��j>?;طj�/��^w0�o8��r9vEZ,H�9e���E�f��%vW�{r
��^�W��H��|N0y� ǞG엎�"&].��S����D+%�������9�,"����@h���u���E(�s�� +���I�QsJ�ve(��O��q$�Ɔ�����E��l8���wJ��I%H(�|���� �?���r�
��$�|]��u��R>�ֱ�����GK�宨�m�����Y�2%0��qbƸr�"�����"T��k�՘X�c��*|�����k��32�
Y!���1�2MͯV_���l���>e8���}��&���8�s=ڭiL�h߻u+#ve���g-�U�T����������?.Ya��(O�9�_���3��VH��P��D��|?rhl]�=�Thd�G���9@�-�Fl��-�bw)>�!\��r���7!Ѐ���"~zzBz�6[Ҁ�4�2d�z�8W
#�����&o�_���*�h@""�
��5���"�9����z�8X3���I#D.���ӎL�K&�������Eh*�K'����(�Z��Re$����3K�A�����4�9}X���M�!����Nrr���cxB�z���ħ���_��~(�T��n2>�X�HaxҘ��h�p�<V��a_��.,����fZ=r��~��mʇ%�Pw��Gg
t���}f-i���)�Ҫ����sp���0�.-}Z�_����L��8�][3�G�� w�Qa���.V����tQ�.���ez)��nh�mſy�k��0��Q;W���G�u�ۍ��"����������=΅�+w���"q�{7����~f��6$�\ ���s�#e������/�sG.�6���*�z�FD�-E�f+G"O����͢������c ����rb��XP����Dyp�G����]Bt��U���
o�
")jW�!�͊WO�J_�,�1����H�M4�H|BkG���0@(cZy�1����Bc�&�������S>7�=�Q�o=6���k/֔L&��A���KP0�*Ǐ��n��<OXٜ�>im(7x�Kl����)�C�r��`s��d7܂��5eɲ�.�߅J�卫j��_N�*��Ě����/	������e�08[�0Tyh���׾sͳj���<�炖l������G���ڃ�������R/� oC6�|�^��`��"�rW�#9_c��4��`�l�]�3��1$���M�j�Zl�����r�
&���-�T���u!`_����ة�j0���D��q��iN_��V�K>{م�(��������FΫ�g�WS��ϺX�'�qI�y_���G�;K/����M�?cb�"��ؿ16��O=���y���Y�Ş��@�%��d^ЌB�#�䈹��C���䷋O���SQ<����J����P r��.:ۓ�&�_*�h �i������3���[L��Ժ� �3���8���g ��I �9=#	7{#NI5@�'x���u�ƹ?�I~��CÙ;�������䐐�#K�X��b<��H��MblUE��0�G"%�'���דL%G4�w��;��f_�E�1�$m�&�;��Y����=�G�c6'���3,7h==�C�E�V��q���)��&���q�?n�0���-]	�Eb[���K��O��zW�8�:��j�����n���MP�
HV�7��s"����g�9F�^�L^�CiM��"`���/�$�"��65���b���}T�'����ܷ�.�c^�r��"��̡?Ha_�S�O��</�#w>�YԶs�G������|8sOND�hM�׃cR��J=׉6G��eL �\�������
l:+���`����l��Yr̟���g@�k�&�Q}ҞuF(HO��w����-?O���0�c�܎ 1~17����[�a��!�#�ch� |�k�c�"ݵ-�"S�FN�Qe]�r~�i��x�25*����2�|h�Rz����S��ޭQ'�2���( �7&���nz���$=$N�7~�j�=����o��0zgl೎�įIwO��Mf=�:}��I�@0z��<�Q
�����(#�V\6��_%�(�7�(T�x��$�Wlj�c�GS�F��1��Y$�ȼF�;6�;��b]��H I�\H����4�]�B={�ۦ�2��Sm(»4�l#� (^w4��3*>��hCDK���}O�fDk?��c�ۨ���ݑAG�����^F�ڎ�VӸ�*6��7�f2�#����|qد�����\��|��2�qx��gN�*m�b�	��<0>���;c�t����uˬ�ܚ9�-d���"�uA����@���3��>T�-;Ho�x{'�^b	�u��1����J���A����$��|�����Ț{C�M�F��d�;Z+{t��q�*��7	�@��Ԫ:m!��[✱�X�=!~?8[�8(*ne�	B�;��[�9�|���^^^T�(�jRL�.}�#�M3|�`|�곿���6����9�f�U 
��Ś�6�p%���Z���F�kS<���t�����ѡ�PHr�$�j�.�u��V�e+����C���L)#�?�=8��C���<�Kw%�~��T�PT)뼺��̈́!0����������9�.[��ȍ8�/E=r i���;no|�v�x�3	[x�5�#��_�SF
�k�ZK�.��B"HKbJDM�9��ZN����Y�W�����8���o �l�;:��E���L5�X�Evo���;��%\׷hDm��H�y�	1r�R��[�s���#�$�i"�� �D���Y1�\���n�Y�O4���o򤦙>$�g�9��\I~�4�%9u>k�$\��|���zj�ENN갨^*{�]��s"7w��oP�4|��Y�?�`!.]gٕ2x/�#��L���G_	�z�A�	Vyp"�N�z����-�/?\�dCǈ��3�Q�h ����Ǫ�.���\��ԥ3w+m�;6�r�$0f)�mn��S��f)�MTk����4x'O,��N��S&��@��k�s���|9�L�K��]�m�J���E��7�Χ���f��b)S�s��˪���[�[� �ۼJ�ZR�&�
�}�E��KX�%D��>���Ơ���?Fn�_�Wll�BYg���l�J���W�%��A.?$�-�wm绔�܈����I\Y|�4���xķ>�:3a���m��Ȫ��j��x�5�qb:��l��X��DO!�
�����}f�:QV��b������}��dW@둃��*X����r�`ٖW[���[t���=�(����dS��$`.�C~r��;��,��m�a�@qt�{ՙƋ) �E�N&@F ��:�) qieT+��$���*��i�R^֟��6���[����fg�  #m����������r���,�ٻ������B/��C&���F���=�i*Cq��a�W�s��$�O�I���ۋ	�W򸫃GB�D'�֌)�"X�#��#���>�d��,4�S�R7�x�;Xc)���H.��\�h���(�i�-/x�G����o���BY$j��������9ȓ+�����YȒ�k������y�(+V���)mo��X+�:�e4�̮mR�.¯�V;�Y���X��-�ǵOJN�k��6�TؖK�܈�ΐZty)���s��B��0�R�{�n�Q���sZ3�6��0. �S����vx;�C���a������<~���{�eD�����������Ci���'	H����ͳ�D� ؊o�H�R���A\LǞ5�~�d�xp��2^���}V�_��kDY���nv�)t6��u��c�)����+�R�\�����\���&�1˧�Q֚yǈ4}���6��WON[�YV�B���Ja��a�[>1��~�-ҫ���A�4/���K�����=��Ev�ޤ���n�?3�c�U2�L=r ���ov����������J;d�߄�(*�����t�I��D`6������c�ҳs�~�����xLd�2�O�HX�dnأd'P|��Xj�I]�*tf���ʻN��sK���0]Kt��ԗ�4m�+;J��	�#�	H�J�-�W�Z�I\�b
	c�����GD�7���
D��r;��9���a�	��_�>�N�d�^P�����@-�%���	3�EF8a�s��m��<]����ɨƳ��|�P=L�GM�F+iS!��q5�g�"��-~0ҋ��,K�6nZ���w��ePZ����ۊ�"W�\H��5�g�ћ�y���f���rgJ�<Q0R�Gw��=<hI-,���U���2�q�v ��(_�`3��O��U8.�B�ċ�!;�j\̲�~�8��H[��DG����Cܱ�L�X�K
\�8�-��D�F��(��JX�ƴ��f���I��i\��:�,��eω�~����T�o�f�BP?S�GU!�*�A\��Z�8���׻sn�Wo��\S ���c�<��C�9��n��U'%<13�q�bʺ�$��)�:D4-�&�"�M��}4��8yc{�.���"Rܻ������|���r��Y�K�Π5���p�S[��?��gDr�LC��v:�aAG$��X��8�`6!vu�F$%y�e��8���tp��&�������s��@5�@h��н�\-2Ě����U��-�N�8L��ŝB`��T���jEV9����%��Z��F��w�vQ���r�f��U�e��xߏ��d?�v�oh�)j��J^�EŅz�W;��,��1�Y�	��p+{
N���#��=�z���sr�6&{��T���<$��-千�����+fᘮ��̚���Xo��S��`@?f]���[����&�:?>�l��|�v�r��G,�~�ihzN��vb�7$��s{H��(��3ǭد	�nuO�����b��2#?O_3�.�A��Յ1�h��h/.d^ʞ�p=C�0,�c"�('�T�pv�u�[
��� �
����B�$;K��pq=�3�$Ш	`�.�b�)�6��A"���9��[�}���}qzG��&'�����M���\�7�Lx�/���p�4WG]��X�l��?_�4�+B��r2���mo{�����S�HK�e�H�y�\y�� ���	�>����r����j��^�?_�$kM�߅�Vy5�4�4ᴣ�&f�dB��.�N����ET�2S(H�O�>�Tz.��[���;��5���t�=�+=
Hg�[ӡ\ϰ�ny��F/���nEt�MFBU�k5�p-�� �C���gg3d
�������bʻ�o�?���7��q8r���,��J	K������A�8u \�HӐ$^�&JJ�͊�dOh�䅋��� �/����!*�����t�,�H~�7�H%߅�!b0+���Ů^��o��cp�g].�e�#J �<r���[��.^��(���>
�n��3��A�O���;z�ٺ��?-��8V>��C�A1�t��"*��Y(h��x�<�a��5k�K������\�2'�MJ�\��P�r'5~���8Kx����E�9Hړ��o$��l��cT!9�P�D�4N?Ғh�J0��<r��V��R��iEމ�*���k��D��lә�ʑ�H��1a2E���	�"b�鸄ݡ�/��%{�KȟL,�˪N��KPF�g��l8M��5���2Eyr�w�Y@��J��%3AZt�����p(�?��;"Y?+��t3�Ch��~	��Z ���!Vo�_��բ�S�<�=Q�z8?~IT܍�q�ĠV�H����kd֝�D��Mh]� ?�fx�hV�^h2ɱP.�?'�X
��sD���Z��}�` ��j
ct0���n�ޫ�,ck	K�L0ѱ�n_7����6/��z��.���2t�`J����!�}��ӟ��.���\��b��䧏k?��#���d�l�J#2hFA�I "����C3N8�H���'�a�\G$��p;����z'�߈C��XT��| e�$����z��s+�>���9;tZ��ۡ�`�ؾ�u߀c��vv��e�B�u�fȆX"ܱkf�^�dg�YAO-Y1jg�t�k�M�
��$��vi�g�x>@��si����f,�0������|J���G��t�n{���G�\�fk��'v�N�$�J"V&�\�5&l?���>�p��i�*bҹU���T�9:2>�����q�D�V�� u��&1��;f��e�Ce�`TTղ�-�l��S����須��l��?��"�(x[�,�Z��> ���ֵ$@Ǧ�~�"��9�œM\���2*K�?��n~�.�7�% ���C0Ei����e$��EdS>S؎��ḿzP|d�m�{�m'{B�`)��ͱ���9~�bi��Zo���-C֛]��n� #pO��Mr���v����7��_M���ިZP���'�x�����K���J��~7ڪT�����.#c���Ϫ�4�M1���t��ѨBN��̥@d_��ykq�D4�v͜�(&��E��ϖ=�n�L����<�-�,���䬖��2�3�|y�Ș�W�� :v4�bw�תXtױt�?
s��юb���
Q�\��U2���t���Rg׿=d��x�5y͡���,�@�+*WOfྫE^�vs5�k��mnAb[����vR�q|-��
�!P���V�E[N�� %ʊ����A������h��`�M��H̝�aaw���=e_���:a�{�-5����-��N��ѣ�d,W�6�q�ȩ2\u�]-�X/���rI��d�4��G���ý�N�6����/����'-��;ڡT��:���l����cދ��^1.��#}�u��Vy�=�,� �-����6>��_�����hM�67}�Zb��̏7e����|Č"l���51�^��Z�(��
�=�=
$ir#P��p��Y�{�f꧇b��vd�H�Җ�
�
�|�����f�墛7bӅ7�c���x7w�ˆaD�z�Я�����X��9�R68n!_	����e�%��֎MX���3|���'�5���;="��@"���Qv���#1���M����}Nw#wc�S\|�_+��&��Bt��ł�L��.�������n�?�U����M$T�������G�G�_��G$X�O�$7i'Z>��bU/�'��j{�ǫ�)
+K��O�G���!5ճ8�*,iT���?q�F,_�{��g_���Τ<����z9FD4ig��BH>h6j�5c3v	�HF8�m��]z��\D�fa惌3V�x�m|��m�y}�/䶤����e˵�C��x�}�n�_�Ȝ����Ʀ?7�n�`��gRK��y!6��xN�Nx��5M��T{�
bu�0-Ԯ���á��ނ����"�"�
���
�@�G�b��I(�a�)���v�s�>Q'���5�	��p��h���ɉH�Ḑ��_��:�G��z�����[���0�"�hv��pI�[ɑrP [�=|���b]�h��S(�րt{k�!*k졏78T��t�X	PUy.�Up)�륉�(>࢙
]|�|�H�����O,�Y��rf)�2�%a\dq�-Hv��q[=�n����P��i�b����I�L[�Z��؃ �O�w�������z1��D�j%��Q�-�}	S!v2����7�D"^h��޺�2�ˆJT�7���H���=�5i�9��3r�v$KX�]��#�s�UL�]�8����o8Dk*�[�#BoH�r�|d�PV����!�Y�A�<�B� �Fc63�6�Gq���$E�v�˜�Pd�}��SZl��ug�N��ns�`�<�O6��'�O��N�j����m	A{�.�����"Q����|���&r<^�1өcA�y���5L��?��K�OcM��u�x�y8�KH����ކխYKր1��'�_��>���IC��q�!E�.KT�p�;�'�y}w���E'��'�B�� ��������]����ux�AFP�^܇QeH:I�1	���f�q�yU]�P�Ib�ب� �Bwg�N�V�Ų<le��~������y]�H����X>�g�����^��§�����U��Ӊ��C��~��'K�/���K�y`v�Cy�lg6��`.�I�TK��l�+�+�&�#�
4@P�6����"|�Y�)�ȠO��ZXE���)�Έw�[�	C�]����`�?�I���&���L�_^qϨ>b8��\�)�U�7p�x�R3KO���6�v�uT�)�`�H��M_��c���'C���8춊�aB���:]G�����3�(o��2���cm�"���-�/�S�Ƌ	��1����Jm�����R�c]�h��D����¨ ���KJ������U�ή��XȢM�õ�=���d��L����c�S;z�>"� �fq3�ٚ�A>tb�Mi�5ߘ
����˷�w����`Pԕ5h��nb;9W�#3���`��8/*��f�E�����S$�F�`�FN���Q}�>�|���;;ݩp�n��r�ʋp���V˚ƃ�

��Ą�\d�bI�x�\�x�sL���Y�	�:���3�b�w s<�k�V�����c���� T�]Y�X�	��Rm��� 1~2����@��W&ǖ��yD<�a�kô{����m��c����d��q��g+r~Ǔ/-�I�zK!�vv矪/r~�[��!��.ŋ�����-�(��� �*�
{�w�=P��C[dh)vkƗ6v^&��[��O:�1z(�̳�=��1�'��k����j�9�f�_<&�wKέp��e^�F�����r���c�1c��8h��Y��o~˅GLҶs��ӝt�r��CQMn�6�]��,�[`Z���c&�Ocإ������t���gS�����t~�A}��b�^f���'=� �����t<"���L��O �i �:�(�����ZY�����1	|(������Kg�a�aY`�0IFfA
_��48���X����*W�i/�O��k������.Kx�xO�\��5i��D)�����nTg�5����Z�Zp-EΜN��|Sm��׃��>~���Iɲ�5[X���sp��/�.n�R���J�0�h�4�:�K�eaqL����:��7˫�G���Ǩt� xA��`ڬ�����Cf�����µ��2޷��b:�뵕�Z�i��]n��Sw�aOn�� wIC�Z�9�|��K���BW�3�P�`�VĜ�N���j{��d�rCM�r�������3A?+�h���tyZ.�����A��@Rб�\�ƾ�������ϛ���7B@X�-��E|	�������Qr�t����)G�!�2��1Н)����*�_���=��	���d�y����!f�0J�c��,Jڝ�ЛV�ģ�@s�n)��E'/�oph�*5����Z�~S����dc�G���n�t��q����۳Z�g�8�]v6�w�z�,ڴ�e~̻��qq��r\�=/��,Q��B��f����(��`C%ϛZŴ#;.4��=|aOE�P��5��'��{H�������y�q�yA+�!��s�-����3C�j �ݥNk@2��K��I�2���z8?�� 3p���J��Gz�O�ec�q�c\)���䢿��6(�P�(P�p�`��:�e+ �HM^�?����G�g�K�t����W�ѹ(¹��%���L."Ҹ��1�>K�����5�r>�r5U�S���#d��W
����Z�^�(��_<NciTsg�a��2$��ٍ�.]���>�'�OA������xI�;3|�. n�	���	�謿��h%�Ъ�DRi�wI�ZD�3���e��a$;��t�`�@��t@n9�{ǚ+�`h�e�'��?�}8\�=�?����ьWFOtn��Ȑ��w �W�J�g�Ͷ�{VD��~�K��q��s-%j�(�~�u�H���g��-��6���$�n��Im_�i1g���ͦ�XI �`�W�� ��j��qFU��Z�nGЮ���
��omBU��9��W�s�!M�9�U��*"�+��\��W��c���8��Y��v�%�(ȧEq+�q4��_S��� X
����hɍ��tM��:a���|�[Ŕ,��o�l�p�$�G�e�j�����C��vopG\��R�%M�X�I[ ���