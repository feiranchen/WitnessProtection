��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�ƶ�biA�� ���N���X0�&�2�U�i�zg�����9�n��#��˪>��8��_��^q����O�t�m}�6+�s3b��{��W?[+�dxm�^�T��ס@4o�u�� b�E�$��H�gQI�1�u��{�`���M�3=�Aib�����3q0F������Ѩ,�&=,� ��>KWG1<����S����װ�[�?���[c(t��{8���ȟ)�
b�&��wk�ɢ 6��g'[/ �6�q����o��y;a-�憒�
��;��9�F:�̠c�ɿḱ'����
���L0�8w�)�k�J�M����i��nG�4���J�����Ȳ~|� �'#e3�nO$ǯ;��z�-	|D��/�@�C<�Sc?n!|�1�U�^����(����[Z�^w/�eq�o�7lf:C�����F�����D*�cDf�Y���N�IK���7���%��̥uǝ.~XMy_�dw6�S/�F�g���1#U}���)�r#߳�:ڣ�Ch5�Rҁ�F��)�G���I�c0��OtX=����SK�Шe��b۔c�D��T:���3m�w}� �լ!�� H-��i��s�l4X̿\e�bRt��BK[���gX��TM�A�.�mI��yM��8�|��������L,���@���������ua�Xe�{���;g���7�w,&`��,/q�L7�� �i��xE먛ڊ��d�uR�?Z|(����ۧ�]���`棛u���?9Sw
��^���\u�IpeF��?�x�y�*���R�~������w��2��E�}γE#:��u�B<��)�ep!~x1�Bm�A��뻢�4�c�����U6.�!漜���EуW�M���3 �є�Z��lޯ�g�T��_���zV�zzUE%:A�QU�$o5��1T�9�ð�����-�EӰ|{\���$A�;l�>�4�]�MA��6���T�O�1D8�j"C�V� ��J���Ba����?=�����^ALU�4��fHRB���KYA���������k��b����X�{�V�1�����-�;�/~u���~��{��ԝj�`��J!���o�-����X��~c���� ���R=��ԝ_(R�=�G(e9�F_<���=;��qp�=�R�A��v]?GR)��8�aݪƬ�l؆H8D��<�f,%���B#�MrPx�c2ȿ�x�<��j�&�2:�j�=�͙8��|$�#�\��+Gg�T�r`�!&g�ijDI�2_k��	�n�m�б��;�#c�\q��q~�0�Q��u���N�
3Q66�{'R�L��Ѽ{l�p:J:�q���+�2���:�w��Y��S�����{0�_\��b,	�V��T��|�]tV\���x���|V�����K��šj���&�t�AYNw7Q�o��i�G$�)��t\^�3�F^�{��h�x�	����2)E�̩��E}"�k��SF0~�z�/th�9��Ɯ�Z@=�2�M3
fe��v�&V+i$쬶~]��p�-�5z�j�5	7��B�B��W��h�3�꽡G1���C/��و�Or2�ir����P'��#���S�uBq<s_���� [a��������D������u�BG4����Ӣ��)@.>��6���%��������'v	(�0��^���F��8��t�zN����S�pv��'6:�լ��,P���|��N1]��Gn���$�fs۹�0Q���`��٬4��] lă�J�"�����^�),�$�^S'h|\�j�]~�7xjKѥ�DWU%��~��֥,��bqf�p��?U���#ld��*rjl-KH��w9�60矃�VGz�Y��U~��Ig+�u�[d��>�/��� �y
��N�m����'�k�<��)�P�f����Q���T�gb����/���~�jć�}?;��D��UA�&��Y&2�`k\��.��Y�K05�ҙ�j7Ѱ��q��/)�xi�|F�����?�G8����	��Rm����^�S�F�������|�N/�ݭ�a3�L���$�n���{���b��W�}�n¨�F!T	n�a
��tz��7<��- E�����YC/i��.���N�[F9%<���L��'R;c��1��Qv7(#?�{y2%�tY��]�J�籦�~����Y���jh���B�O)��$�;�ڸ������Dq��=����Z�J�<�z�4?ʆ�7�R����!�
�3K���.��崋d���YX�.�׵��E�r]8��I�9%�~�p��K��-��e�����bG����-� �k���g��o�sJ!:5��[�3��åN��S	�R�Ofc7�����d��E�"��t���c��Os�[:��/�O!>�Ǻm��Z?E���	EE9Ч��	@4��&�޺���.i6A矋D��4$�S0 �}}�yYR*᪌<lY��=4��	
Yh� ����xcǼ�]�$����4�KH�
89�n��_�Ε�X�eRZ�a}�_��h��F��,]E䱩�#U��SW,b%q�#�Qu��d+�kF�k��L�]���peNg�	���CB7d�q�G�Zr��T��]��k���Ϲ)��̈́'&�wC�L��,�n*�0R�p�%�v���Mr}�N|Zo�z�qĜ��߱����,%1L(�&��]����T�;~�v�^��	N�~^�j����Ȗ�v��&��U��pB�j�rt�D��H��G�Q(���8&��`�j�
E6U,�=z��� �!6�RJ�eJ(�7��$�
p2[据�������2� {�L�(���}@�@ I����1�Иݰ���G&�2\���t4 �l����m\�<OOK�<�����ƛ��9�/j}t{XН6��J�uߙA��H�����H����e�:vp7�ec��L "��h�d�bd�v@��9���ne������BZ�[�Ѿ"�vw�TZ<��9��p:��J�	W�5H��k��- L��6I ���O�߮�H�6Y1��	!3X׆	���7V�oځ�F,����<!�8��S7�G���c�a����w�-��
6�����*�W���h���*��C��Hҝ���`��8S���KHH9�?c]F���I��cɍ�{ͯ5t#+3�x����_��W ���²��C�!~���􈄆m���I{�?�M穖e�����M��9�Quָ�a����_s�=��S���#��`������lG�V�_/���3㙱�v΋���eB���D��XiG�����n�x�v�B g:S�?x%*���G���JT���W��pYB��v�*z���$\�����Fڅ�k]MU̀*�U��!r�5���!&ݿ?�ҝ8zg��l�6��&��}���S�[�@ ���.ß���f�􈎘�w��/u��"*��&�t���B p.H����:=�sLj:xq�����SOgЀNF����F�ͳ�����o��F�1��������Tǂ��0ݽX_ڭ�t3�Y�Oy�U���ۿ�ɪ̂/sO�t��A3:�GC��66{>�ϴ��ю�� �.M��2]�5��A=��HR<(���$�R��oqLmv���*4�m���<i�����	[���r8�씧�>���*z���'3�)I�611���>M���^]l����nY::d�^}��{�k�4S����aRL%A��Hx�i_�-ۺ�X�B��Lޯ�(���co���2\��6M�گ?&�����#�?>���J&nb��,O4�%_�N�?�����CB�Oi�V�,K�;��I�p2�[�a5>��$�*��UD�<���m�5�[�;��������u��I/bu`Μ�-8s�K+c���c��{�Z�rk��{�q�e�ȟ�>�Y �������Χ���ŭĘ'4��6��UD�Өɾ��Xw/������d�\��`U�����& �m��K�<;��D�>����s$)+Ĳ_�ʫgD\F��pt�ɒTP�C'%�ȫ��>�P�U吤T�O:�ȶ��q��tY��m��(�\)h	�N,%jw�R�`8���W�g<�5���)",�<��z��`Q��)��m����� �T%2��I��9���Z|'׼N�K�j%����"��D+�� �z����l�����C3����1
��"������(����~8ۢ��*u��D�� w����,�Aʷ���z�-t%�����.V�H�5�}l%o�\�Ŵ����"Q5�~����m�����)&�ދ*�EQ-�#�������1AR�RO��nϴ\���K���F��o�UP��j����&ї���FDw�̵~\�x�&�\�,n�v $8Zg/�|�x�#+~]P�OslIV���g����.o$C�Q��%�?����'�Ԓ��(ʶ�sx�I�@35�>�+M8߱��ȿd*N�iX�A�����e] �u�a��n3�gFUhw��L��CH#w>�R�	^��KCܔ^u�y�9�G�{�7C_��������K��R���,I�2���N�n���0	\��xQFT?p3�ΛI菗v�*KrU����64�롇�������ډ-.��|�I�y^	��O��x��)��X��ẙ�^�ߋ� @���NT�>���B��
����2��;��@P������IK�n�Z�72,(���X�������_�t��^x�i�t�ә��+|��v
��ڜ�s�;{��(صaߏ�Ɔ�)���Fꉆ�Ҕ}����L�+�ʻ��$v�'	�M���;��$I{H�nԊ�:RkPľ���BM�C+���cLC��'�ʅ���r��.�t^ac���J����6H�.9�TnL��o@-1A`��
 �y���P�*��l�1K�+CƊ�8�a���T���`��_u��Y��t~����=�	^���_�Zq:6��q��9�=n%�]+���)�w����c���S���հF���>�T6�K��i:K�D��h�}6K��m��yS��f?��̊���W�ǝQ��Q ��1Pg�o���O�A>�V�^ ғ�]�W\���G�.8��� �s Z_3��ˈ�!{%	Je@(�<���0��ܼ�%�â�ݝ�Zb65E9�ַl��T�b����J+#�]����	��1:ìM��(�C�N���f��=J:��ys��a��s��~f�<w��F�B��	q_�Ng���"���$6f����xD?�ǹ���_+�\%Q���G�����ъ*u�Y��*9� �RW~�0����j7��^ފ�4_��A1扝�ol*�b\b0�	���Ɇ	Қ�m�����g(�9�3z�An���(C�4O���-�����*%��S	�Zq(1>mVW
�+f���~0@�]T6�ߓ{���0P��ǁYR6؍34J�����ol ��Ρ^��uS�J��M-��z���@](idű�ɢ'��\T�C`��V���q��]ĕ��K^�`��^}�P���'��&X��Y�a��8��ҧQm�7�r@љ�'X��y?8���A:�X�t�O��;+1�i����W`%�P)��e��,��&�4�Z5)�r���zRfJڸ���äW����MY��z}��L������>��V��Z�!��i$V��"��_ C6��߲���D�c/c/�N��ﺊ+����$V��_����f�be��p����F|�o��ĵ����T��X+��[4���_���6���6�"p������'ȶ��w$"	b�B兤'��Q�p0R��I��DX��1�r#�2[/6r�>��8PQK��ؐq�x�O wl�.G~S��R�84ڶ3N�W�^j�l����1{�Q{�O� |V{�o�JG�ڊI���O�>�"�	�Ҽ,���w@����	�!�/�R8��DE���@� �r��,'S��X?�����z�f�;A�P���~��fa���jpԪD���3�Ԩ�Q��˛A?2�-�d��qʏ(��
����#�+U\�����EN�nNGpϾ�f]�NM�_V���P]�,`���T�7��+�q�֙�aH�X��w%u���<�W��fa9=}�l�'jȻ�I1EIb}aFx<��v��J"��kT�Ym� vn��.|i{_��1�[T��� ��n��)���,ja��N�(�����r��s��?���/=Ր��Z��։o@=��䃧�%��1��q��������~��H��6V^W�\/�$����vM�ـ��=��b���ԇJ� Lhx��m��xx�_<?BΈ\���x�p ���.j����z;<lU Q*��n�9�$��EG�hH}����"ٿ�[�Z����Z�C:� hf[駏�g��1�e�"�k��?_�5��K�ɝ�\�Y���8��X-Wnj�' Kn<�y\�Jt���5ܬ0�6¨�v	�����We�%����5�j�,i���;���q�ر=K�.a��P�$I���N@���mc�'�Ql�7�")�`-���_��y?���y��͐b���A0�+8�p� �f��7��K��~Ӝ0"E���5%��v�*��W^�	�csq��Er�t:�-r�����d��a�)���S�k���ۆ'���/'�WƂ�_���-�X]z`�;͝�r2��J%R`o_)SHK�I���\wW����6r���������V���wn��K�}"�{�\.nt���j��>�i��X�NB����T��.����O��#�q�������H�/)u>�Sx�d�N1����6���5���)�R�3��XN�y~���xZ���7S�?�K��&�A.�ZYX�3e�P�Z�1n�^�