��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��x���y�{G.z�4�qJ?�8����{4�񂿉����r�^�������5i���c.��9�K�u���z�D��x17��`�ߛ��˰��.kK��ӢGϟ�y*w"�9x*�j��;i��[�d�|r^=+��u���1�����U����@�6Ϋ�*}��<d討�ò�x��q��F����x�E�'t9�ˬ�j�GR�Zf�����4 1y�����?W�;k��jr�=h���ʨ��=;��� �$�����Ǣ�a.F\4����	´sF��D�䃺���0���\u��P��~?�u��j��<��Cw��:S��}�~��� P��i34���F�jjd��&狑��W�D�	ᴌ��.
9{_�@���%b���k�?_��yzߣ_7݁8~Sb�r��D�D��2�aR!�pVAR���^�W�Wtʾ�ݣ���B�j���_�}���F5��1�7��<y��p�$M�%Rב�w�>����vĄ�3�\���.*e�O���O��s�UC����Z�;�=��=��O ϼ�� T�D�6����l���o�;z�E!���D�7מPDx ���r���x4���"��v�h�cc�ח�r�6C��xm"<��/�cIm!� ��t��HҢ�)[@���6~E`dބv�`�+@)H�@�;���g�Yyǲ���^� �	���]D;2P��4F��(6`�w���m�:���^��H���#�X�o�q����"sq_�^Q���z��df�<_b+ߜJ9x�I�:��x$Y!���<���?L�����l}q-�tSp���Vt�Չ>�(t]�F�/ʻDsgŎ"�,&�f7��l��;2�C��>�,|s�;=�F# /���p��R'��'@
J�0�Z��|�p�`���!�^H	����@x� 21�ֹ���@i�>~!������p�s������9*���-{C����ei�s�P����j�5�*m�V�Ä�	��l���`�qV�ZRCˬ�΄n[�q�>0��~[ￄĢ���rK�zW�je��H@�q�P�m
�G8{�#_�7���Uy.p�W0���H���ڶq��2i)ق����j~L+��y�s�^�˼}ѓ�����_���y���~�Vf�O���
_Ic?/� �] ���M�Wʩ �����E�6p�m͋_���:��Q�Zm��zP��I ?5y�5�um�HYJրv��꒪�$J���<���Gg6�:~���I��,Ƈ�U�0Ͽr�nr樟(U��ܠV�@����n~��Ǒ<�plMk*�I,P9-_�ăd�-M�� �x^C<��6tď�w;Y�����rgT�-����wQNQ���u����';�)�A����� =�o�?=�X���M~v��q�[>y�(]�.��q,&���L���V�=��{�-y$lT������R@g�c�b�������Jqn�(�q�̠��I$�Zo�2	����Ds��M���p�۫����n!O����o�j5UC�+W&�܈{{r�@���o�̋���R