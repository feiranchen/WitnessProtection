��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX������`'Ԇ������;��n�:����v�,��Șx6 A�
���։���n��Wo��~�x��R��E�p�Dv�X�W���߳�V�����9�H�~�U�T�`�T��iw�c}��_���Z$�����_�7���\��t��7W�c� W/G���hF�V_J1!&AG���t���yu��~3^%�f�;��ƖG��G�-:�aW��ͧ��ȩ`�P��T���y�s�.�o�w+9�ʹ�������Oq*���q�����&��DIČh��"�ѡ�C���O�N��e�.��B+�r4E+��0�ʀVJ�:��P>�&���7��k��g�H�3�U{�C��X��� &�����`;�7��&���.s�G��C��&��}T��Yk��map0�çN��&�e+_{�j=K� �Yy���q�����+1�E�����Q+�v��-&���O	�bI
`IZ3�.�I�F@�O�ˆ���ܓ�A�j��]�W�ck���[�(���U�Rq·�4�召�����4�3%��e�)�2� Ot�ԩ�ס\����S
�U��
�
��L���\�br��{���@+k���kɛO�3�/��WN�����h豚
b!��z`o�+?	�hEq/T�:�|�k}�3�Gb|�:[Q��v���3[	�B��������<��I� �4��e���=�Ά���F�J�}�U�gH��&y�O,,�d\�g?�� <)���3��}?���q�c�`V�oG {5��`Y�Zׅ� Ho����,�����N�-Y���l����5V���;:�B~����x�%`��͞���� ��=i"�wn�E��se����S-��q~/,身��w�DJ�z�obv�ơܙjVM=�y��>$9O|��6��hT
��Q�t�6����T�rz�~�����!��`A���C5�M&T�ՓE} Hz�N��,Q��T���]0G	�eU��k�>SN�����M��}i���pl�x4��*��FF�5��c�6ݱsW�*�����d�}I���z�Z�p^�XS���*#4w��r��~�l����/����-���vwF�Tި��!!?�{+�Q�F-.a�'X��%K;t�Cw�m�u��Պ7ES�xK�B�#���'J��ʖ�~s>������cY�Hӆ[X�yNر#)�1�!V�6*P�ڀ06�%��o����ރ�=���{8n��Ap�+�ֽ��d�9��\m\C��~{g�<y�U;g�p�9h#���B�V��M*���Pb:��2��٦ƃ:`D�#Y�O�Զ�r̪ݸ�ᒥ��^)��?h�а;.y��3��� h���+�1G���Wa)�+���QI��ل����]P�GN�~7Y�����N�g�H��Z���H�}�9����@:T�N᜸����f�h�?�R���I;X��T�D�9�3�
Ga�fr0���PBH5��	�lI�`z�c���:& Iw	�qٶ]U{|�3�6� ��lo�� ��W�^�MU�[�9i��\C ���%z0m�� �`��wn�7�I����6�	M����x	�����X-��@�7�������`+l����zS�ݕ1�F2J_�>#�TQv��h����l|3N}޳	Q�ܟ�?_��wڮ�E|B)yf�Q�+>��:'�|���j�����s�{ף��V�$޹���@��W�������͇R���jfN,s���k ��{{��=**�a�����>e�P�rd�	�b�m4eT�EE��h�w���h%������0�1<5�� �D䘸�@sJ�x�`$m#��������ݪ
Qn�Q���A�!(��h�9��zg3����P��b$�d�v�(���i�Q��	_ّ���K��P��)��h�_`�EUuen���E	�1�m��0��K�����~95�M��ЦJ�)ʯ�=����Ӗ�V��/�w5��t�zׅgk=s^��.E�o��]Wm����T���[i��[�!��9�]Ι6���uσ�.$�R�� �A��:����:=���F{hF$�QP U���KP�MlKR�bM�yeO4�^b{��i�Z��%��F؛��ڶ���i,2����Q%��*�9�-T��@1��k2�lwHW��h�ż�2���ۛ�׵4/�j@B|��M�b�`��S����o*��-�`� 
���b��>�ѩ�����N��/�c#�!�6�y�}���?����0�~;��v�,Q{�<�y�n'����H��:`{�>=k78���~�vK���4)�v7�*�v6_�F9D�Y_�t�BU�vҢ3��d���Ln�
;��$l��0�������cU)"E������\��.�@��������Kc>��	d��[��������C�M�b*�`�RG�۔���)c�A����հpsU����[� |�����_������6���r�S ��4T�a	;�q&�]��0(c�� f٢PK�v8�!�� �� Ǆ��\z�u�:v��a�O�)��[F����ǖ�^ =Ȋ#0{`\P��0kIj�,�{�Uu+��c�N5������tY�6�A�#L.�	忚4���D�i�����$�^�N�^$SZ�ۆ�$j��/�#�_#�.��x�3A����$,,�A��H��?�h -�&�x>��O�y�g�)�[w��9m7\��t��*}�B8��~蝞%�a
ˉ�Na�����Fc<�V	�~[w�49B�ARD=���90,Dޘ�`3��o�v��A<��硷L��>��^	*M��2L��{�WB' ��_cu�鏛~�gߺ�\Dy�=����cr�5 PT�WJGոP�0Gd�0�lT�����,���A?��������P�hH�d3�!�1�����w��>�J�ƕ���Sʠ����і��FtM��2=�@!���#�Z�Qۋ�%h�y�����ݛ�2�a�����|"B�o ����L_�=�J')ՍOI ԨT�����Uj"�T����jYO[9��#u���A�o�C`��{`%��mx�Dg�/D�G{JAf!��AGY�P�zKy�E��i(�	�EK=��K��5˓���aF�s��=^�U�.��J�Ow��;�o}i��Ĥ�$�Î��Ļ�O�Z���F$�ԌĨ��vZ�3��B����\nTb|fP�����"���W-�Rx��墫�ٜ��� Q�$��M~�u���$�jQ�>�;�%}K��ń%,e��9��#"v��)v?O#肙��7pw����;����K�x;Aq��3�F��+��=�݂>� 8�����B�nh�*i�}��eM�B�`��ZMo�U&o��q9�°����?k�5��3ae5��Ջ١�Tz�054�Nu�.��������u"Qs�c�r�Qg��h�����7d�����hk���Hw�C��T��}A��k	���8tFV�ȴF�-k�$�l>�˒��d��X6�����9�x4ۯ��o��R��^sb9����k�D墸�C���bi!�����hy���D�X�����A�
��&ݣ�g���!q��qČ�ܕz��1�I<#��7�X�>��Y�F�������)�Z��!~����J��?n��[�|%Ȳާ�rڊ�q�ABfz��-���VK
(KV��:/ܛ)=�M�+�N�q��O�Zvd�S��4Wr�"a�}�����I��;��R���ke5B�J��f8�����:Br��A��IN�ZI
"����V*UMqSr�^����~.p�O%�nd:Xۛ����?S\	N�J��D��w��h)�Jf��B�q�*���t.Y� ���Z���AA"�l�v`�n�%ə&�(�ZjZ��Hu4�rW>�~���{�d�����=�3`���V�h����@�U��2kSS�-K�>�.m�Ἡ��F��'�$�k���0)Lg�VV�><���O�)g�X�A��ݬ#K?���8F;��{���5�vH|z���
�?�����ǒ�@ϴ�JQnn:���2q/g;�\f�F�I����!��U"�`@�N�p���i�V
}O���6�Cp�������ׯĭ�+7��|PͰ���w[�8�t�X=��J�eԿ���Yg<�
׋ţ �/�8d4dM���D���M��\P��zb7�~FߕL���9�N��� ��q���4�橇Ƒm�jhA���C��S�H�u|(g�4�gvZ#
ݞ�~�t�qN� Ә������[禢�8���J����(6�:�^v�fU�N��B>���d!�O�y�{aI3�X��8j����4��,���u#��8��ġaT�[hl?���L�hs����7��EŁX��~j�
�*kcLK� )����򞆗�S{2ͼ��<���.0�/�����́j�����0��]1���L�r�o��֏-|�e|��h����eH:r��
�r~�j�"BG���M��1���ߌ��J��]�����V)��~����f/\c�:j�t��S�9�s�Aͽ��-�5���f8ۃ^7lm:Oc�\��/�9��e�$���:�H�C����SNL 7��������a��`~�(�ij4R� 	��G5��`|�z�/~}M�F�kd��O���*jLP\mi���[y��E�B�� ��F��;��F�A��Nl��5�Zn?<�yl#�.�\*lXvǆ�`d.��^`�d�K�|�e��,���ٞ|\���3�fv��־X��Tg�ܚ1�	�W��z��Tٺb�z�e���~�=?��:u!T�#Q�BgM����5�����\�1���Є�����-	0�n���%>,������oE!!d��ȱ�}Ih��:��0a;�m���q�,��d1��拴ފʜ ��DO�j�A1�5��D��ͧ5��g�H�l�_^;���7!��0����HI��"p;始Ba"�M��������zH��a4L���TS/��'���R��-�����1E��7��V�UR�lS ��쨵�'!�ю��&t�Gv>��<�i���B�[%"N$�=��P���Ƭ<zSY���C�A�C�y�ز�X���};!A���G��p��JuU��5�o0�_֟���H?~�O;�����hM����>�BL��N�;pŌ9,�<&�����w���.�S��[_���H.����PF�C���B���w[��Rkj�CA"
K��d��r.�-�����&�`y�Xs���,��p>{ful~R���J�Ax��Hd����O�^F"�줓��37��|r�w��لHO�� ̐n|�d���G�U)o�Idr0*�,�-�`�!��[)�g_`�������@�����|p�}vʩCjzp"��_E]�f�2zvz�Կ�`���V{��d7��*/|�txVw��/�K'�3�it�=��&���;9H�{��� k==����Z�+*��w"��uf��ۖ�{.��>9��VQ\ذ�8a�u*S�����T.�Z��}1�����ђ��~׼��k��kD�,��׿B��EW7���;�*����>�o��3n^,�NM�D��и��EY�9m�t�A a5$Ya�wX�P�x��������~#?n�m�d2���4��I�e@���n����N&�)R�z�'�5C&ø�"i�E�hvy��� X��X�s����G��0J`�;XdZ8±}�ޒ�\����%��'˧Ϲ�?4�#�L���j!e�K�u�Xm��Ƥ~�F�\�T��_�����ЃW��ۃ؂m�
�,�4J��'(�jsO�3�vJb�kx/{�e�V?�i:LW�h�\W�%sc����� !׳
"ެ����.�1`d9��;� n��5�`��$r����ܷ�1�j���oY����D�B�#`�$|��X=V�)�ޘ܂t���O��)����}�V��.��뢸q�4�A������(��ly�>�e�P��ɠ"�|���ջfT|�&�&�s�,ݿ�$*��Qq���0����BJ�[R\ưn7�̃���Kx����oOt�k�Z�X׷�4��ˡ<���F�E]8�0����"�6�k��`h������V�sl��,	�t�2�ߖ��t2C}Q��0�X�Kv�\Û�Rn����q�g�i�|`���X�&����I��k4����O�Kd��B��1��˿R�aǴh��.>sB�.سt1˫N_������ɟ��⃅�d�����^N�R�M�f�2��>{|u	��ª���;P>B�L��uje���a����
���\z�,�'C)w2VĊ�:�NsKV@�꽖�����W��L����B<f�u5O*B�]5�A%L	�h>9kGH��lԠ�LCk��bbo�K9�ŒÝ�B=����Ǫ&�r"mXy�X@]	l�M�!��� �#l����O��{�Ċ��z�����c��`A��x�y\�x]_��/ZdB�+�:X�UxӇ�[ɏ���i3$Tm�Fm�=K�@[��KH�V�{M"~�;�k��.�~�ח�nD�2 �ĸZ.� #/�H��3���5�����Y���������rv���T+�/t.4���?F1�5vw�o���d�C]O�̆:;��q�'�N"d����Fڅ�qNy-VL}6+�k���w��:ۈ��UPɆ	/�
��������M�y��Ȉ�DW���H����)������B�\��^2�� $.ŕ����n���K���7���l�uVB�/�IP<�0�� j��Xd?l�Y85$� ��
F�iq�I�2dV�+�j��km�����I�\/���}rn�䴽�����%���� &QeO����#Fk�b��ʹzJ����||4k���}F��8<Cu$�
�2�c�C0j�벴��[�smW�Cp#�[��f8G�V8�`N����d4DwW[��$����r/e��33�u��o��΍�A�}�T��������#��[y��ֈi��ah�l���g���Q��8�[�����]���>���J�A��ܔ���M�:N����f�8w�dK)'�|�?��Z�r��BW�ӡ>E[�~0K^�	\JF��.�6	,f����ȗ2�D�O�Ȏ�Q�ϟ�/�c_݆y�1���C����Գ����{n2�y�� p�J�$Sxܗ��h�F��ssl9�v����9����,�sx n����ನr��niN�%S7���m��g�Tj�o���]���R�4=�(]����I|��E����vH��7s�%�:��A�]�]Ѽ?<�f��1I�ϋ�3��Lw���E&?�{]ΐ7�W_��pޏ�̎1[���O�����gѧ$i�1�<%����: �����)=`�c2:c���yٓ_|0�ׇ-����-��'�,�ȄUP�D���'��~����!���e��KD�@./�W�q,�CZ��"6��y0�|I�Q1�i�X��1A0I�pWٷ���7�C��?��������o�fT��([�ɂ�.�r��fr5��jJ���yҢw���~+}B��i�g<���,���P:8����=ߞ��a���ܼ̚��ř ��5��X8�k�t��X0ƭ�g. gF����u�~� �G��z�o[D]�9�+�G�ͼf�04az��O�W/�A�t�'�E;%��ϼP}~��)u�&����w��3clI�g�i-`#=n�̣^��"�$�a�a�%�͗�*!\;P�����R�r���j�-v�<.)���Y{��K@�	.���F%\>�h�X@�Ь��,�ܷ(��악i�{/g��@�Ę�?��ğA��#�&�P*4ↆԼ�����SӃ�����E���uVY�|oʔY�}��`[��!�v&6��G��[P|%�~"�<�	�P���!f�[�c/�ry�/m������(HJicz�]]�B��,aJo�Տ[��J��Vx�^�<�	���h?Ŭ2�Z�8�W׿)�ʃf�퍫�Z�[k,I0To}y����XL�^�������m:��}�[�mα���f�F&�^�j�����+�:S;�.��	�����SM��N���8�ḷՠ.𼫲^��\���"�{@�6ɼR���o����9L��%�*�v���S޺+�ی̾�zxyKM7��h�T��*ր�aڷ�-�Z,$�͙��n$v[Bf�=�n�ԏ2�1���v��o[�����J��:�u�����w�96�3��ŉ��3H�x!=�-�󰷸/�(�i��5����9~, F��i���h+n�A���!|���n�mP&��Q��y7˾�_D�f���zp�D��ۀ��Z���,1/p:��ᤊ�������o�@�J���3�8�.d��(�z9H��+��'�(SO��/,�g-�����h��]Ii�!��#K�8���ױ4�Ti��g^���"���j�Iާ ���= ����U��k~�6���q5��/f�80��P��(+�ҿ��@����zg�2،82֠Q�BɉqI���y
v��W���H�ȭX76~��Q�A����|n7C�k�؞mb�b$9�4)�=R�K���� }�=�Mu��_oK���ܾ�0�tF�ӣb����9�Ȣ�"�D�	�JOB-쎰}��	~r��N� ���W����?���������f�eԂ���k����8C�|����Q�]/�!6�Dq���m/��)��y�!`�_��{��,H.C�m�FÐ�"�����4���)�������{�S�b�G �G��H�xt~��i���[l�H�6�]I��m	�%�B�x�Ifv����|�����������9�=	N�����흷�-��0��ְ^��f������W�r|�˂	N���<��R^$�Ff�*����Wѓ�rC �:��N;�h���z�3�@*��Z��<	���><H���:9׷so/#���)��v��A%es���~���ހ��~��3P�2tR�6@<mg��|^|�o��h�b���e���5x�v�oo���'�x��!n�.i�2���,���H��z�"�i�_� $b� �meӯ�cx��Ic!�-נr�3���
����`s�+����_EO�����D�G����<�)��T�:]��Щ>�8Ndˎ�󅁣|�D�L_
J¾�ӵ�{�e9�tY$�{�͘��(���Σ>'���q8y��\�ɝ�\c���Gۊ�N� ��������zR{N8�ﯦ�����>7^�\��V��Mb��f�2���IvH�����v�(�+��*#��~uC�5�q���XH��p2�/�>d��rq ����%�U��W�j�5�C5m�\s>S�!��Q���.!BSs��Z��T��^��^�',Eagf�A��Y�-�LѣB�U�0�Ph4�ep��A�A��Y\�������u)֒.s��Ի�e�r �Ykfn���>�� �ﳦ�?�ȧ�+������T��[�h�O ����+JR�h��R��[k=���O0��~5{�Y�� J��C�F��5C{\�=#�Nybqв����u-˚���N�[y:k�eT�/��y�;�A���o-��1C�:�bkj�-��Ü"gsY�8��=&7�����{߄��)� S�o3��y�F�ޝ͗%hZ3�o� �M{��!Q�S���M�+�d���ؒ�&͜B|�F@��!T��Xj�	��T{��_�6�A\��� ��{��Ӷ×:~��d��%�ҵ��;��F�j��!�����l��->��߯��_#0rZ&�{�������.�����Y�i{���I%3����%����^��1v�X��V�K:_�ws��}/�C~L�]��e\9��,�@��F�>��kL����}09K������;�m�X����i��a��Zt��f���\��j��;��T��5��b�;��P��i�Ḡ	�	=��4:��NlYB��t�Ir]�wt-�뀼�}��Iuh5[i�u!8��P�q�PF�sq}���?b��%7�Zm^�Q�;��Q��͂� �1�y��$=
��I�] Z�( ��/y��,ؓ5�����W�q�k�������q�#K>�z�]�`{�6��K��qH�H��*�<h�,	�*���̵�>i�SK����^^r���/���ϫ*�	��[mۘK��h�G��g��uE��p"L~"j�&z�Y�����"�C������������]_7�t́x�0�a�K�ȃ�!�"��K���jFQ���Y���T^̭n:k�7	��ѠF\�W�s�bl	���m���D�MB76]����v����4�F�6�������m�>��|�w��05&����AlTg{K;��a"���V���Ie�T��骠�bf3nJV�YZy��a��Ƽw?�$�#������Žr�2\"9/[����w�!�XSEhԣ���o|���bM�!����'����^��Z�OoH?�@��Ɔ��ȃ��^�a\H�VQ�%��]���E	�Ūm�9ƅ��q���G�j|�%1����:�==����U�M��sD5n`���`Z�T=����$S��£tHh�+	���b�Z�MP��4=(�xe�w$%��s|p~MQ��K[Eb��8�&�'m�+V�)�6��3�N׺)6��� �L����rx��q�+k!Y���������j�O`9�}��-�n�I�\�2jP,pToW�Puo�V=
��w�Ր��`24_�Y	V�5t���l����T�f���;��VY�ߜ;���Һ"Q���{�6E)�T��
�8o�����g:���"S�[V2�ك�)�r��y���1��\�NF��Tx�b�
�b�H�@O{p[,k�<�۶�p ����NP�]�]?,>��Ć�y����-0�SUƀ�O�%v&��Z���d�4�'n< �����_>]��֨�k��݃�E���+�),X6Y�
 x�S6�E��,4M�*��_�j�x#�]!�)�s��p��:`�N��y�Q�-���/;N��չ,�MQ�7���]�}د�9�����㪒BH���-#�N.Ґg��ȿ�\s�X�Y}���<���ަ}=v\�� -Z��'���l̤ؒ�r�v������.�����kP�\`��|lDAa�W[�	�ēz��!D�ո���EZ"���`�D��x�����@��i�����68�38�aHc9�����г#���Xcv�gY�%NX�L�T�}����:⾵��S�H��_��}���}����"U$��V��P7���Gp����w �Ϗ������K]�ű�|1��we��#g~��}iJ�SunI�v�n���[Y�@TS�/���Ք�3a�K�=��ng�[ID*Oa
��̨ۇ?�����n��H��Ҁ�z���>J�~L���N���cJ^W��r�9��!��У6������f���o��#w��R#"c�4���?�3 x���~]|Ii�՟��dַ�p���+?x��aYm�D��}h0� ���6]V�0{)OK,4���,�vϵ����Il���{ w䏏�#h��/� ����m�%�Dv��&�t�'���QzЦ�"����������Ed�@�|e��G��R1��Vg.�V�7L|]�	���S���&Bd}P�K^��,�+��TL3 f��lL�����J�zb$?��B?��rڌ�V �B�"��|7/Di���w�s��'���������_�27�:��T�����zZ�;��i%�dn�j�y���b:�ɧg����	ӗ�MP��̅��J�Sv)<��Q09�e��?3V�/��s4��O�Ig0Բ¿�yA�ӣwk�Z�P���2��>o�~{�v���R�����HzSR��Mn�%����?� ��<��T�/o�+4 �J�*X�?y��^����g+�w㎵�=��}P�00����	dl.Aҫ���tZ��x�r|ա�6��:�k��仠q
U�N��Pz������V�c�LR@����v�E�2���i�U#Gxc�jӿfBM�����+�!��׊T��|�]G[������nY@xK�y�W�^%�@��
�D��T��DtM3Nd�o�����$/����:��;ڮ�sQ���F0�i���4-z��=����1�@R�]Th�AɌ�%�&��AH
�.O('��i(�$Q�mq�p_�X�6v��[�}�C�1k��\�k�K�A�5�.�|��+�t��#b|G$�H�ͱ�lvjJwы�Y��]Q7g|A��B�n2�+��ib�P�&��ʉ�t����^k��
�!��6/([=��7]~��"����:r֥]�/d !��sw����[��w����ژ F����� ��k��*���u�¯�v$!���e��Λ�7���uyF0�	ɴ��Ak�\��:�z�տ5��.��3N��hw ���"Zg'��t�e@L�C��SD��o�	�a��m�q}�w6���*��k�0-z)�HI���shG�5+���
4������m�=+=�O�Oefae��<���Kd(��6�<�;|��n�H	H�d?�Q�ݦT�e�a��(���j��+���dt������K��$\GTT��'��%\��P?�`%ONg�ÔM�x�Qϱ�<U)��'qR_��g��~x���#w�Xk+% ��FX�T�"_u0��(����R��cU=5�>���w-ڕ�?��K�6�<K�8R�L~ٲ-��x�*̴��:ldUԉ2�����%���K��Bs�4B鍅6}0!�>�#�V���\�����uZ��m�,�
������"���E����D�>X�6�`��2�ܦ����3�i����TP�Q/1�md�8��TH���Ǿ ��#�K�T�/�9�l���W;23Ez�h���Z5.M�mG��L�xS��:��s�!��b!��ha�ݪA<'R�R'ӄ���J��Zcƃ)= ;�״����Ikw��W�Vc��4�|�x�_i&�HP�I�a/ƶ��l�-��W��}g�W|_���VB@}~�_�_S/Vtd��H�e�{	���kD{�^�z�Z�&� r�z4�9�b�-:��hD���i�}�"(�M��۞�פgg��>��nv��� ��}���$9�|����?��,:m ����']��B��,.N{��D4({Df�/�{��$�f�pZ�C�cG�r�`4!�&F�f!5�ҳ��,Mvd�b-�F��C��b����_�P��V+E^��W��&�i>���`:��)�o3�Ç2��D�P�@�9��%������u@�p~=uf��֫���͒���"ӖW��MtS	7�BR�@��W��@�[(�-ű�8D��N��vr&�6��pMU��'$u&���b-�.�X�nfB����bw>����at��Y7�����Kz��Q4���r�Vi4J��4d^�v�PAQ��z|l���=����O���A� E� Ln��~�s�V�I8��ڳ�҆�����r����}�Pȸx�#�oZ�wJYj��1�ͳ�y���q���u�) ߑ7�H�tim$�p���K�)v�ST�25e�)�?XM��וC^W[�,��(�5��e:�,s'�M_Du��o)�M*h���buޜn]�؟��u���{���8S��+.�J&�u�3��!N���<)rX1���I���Z��5�X9mZ�܋?S��ٜEs�Ď���&Td�Th���%��',�H�:�}	1$_<Ms�i�{�:u�u�#���}�g&|%lC�_ȹ����!>��mgi�a��34��G�!C�{$�`C��f���A�M�D=�+�p��Gj�Y��a��O"H#��;�yh�4�`u�3�`��V��Ff'��Ղn�6�y��O#�u@֖6w�v�(��������H��	�@bR�">���Ո�d^�P��������Ւǽ�����R��q�]J�g�b9(�15n^~������C;,�~íU`=���	N�����7ez��SeqghG�0��r���b��9���	�g���5���f�F"�u	����F
�6$�J�V!�n�fk�dF�Ԃ9t��<����+���䛫xXJ��>��v��3 �?U�T�HW� :�럤�l��@?Ƹ��m�r^l���[�Y���$��vA�Ύ�Ҙ�KE���7'��
�<v�lh9���Y�2t�X5���n�51���`��@�������pMX�h�
ϥ����&��@�����~C|;��)��u�DdP+-<y�Lf�,ax���G�P#�����A�W���,���㫓 �	�ɠ�%��T�RbQ�����
4��
�����И�6�1u7=kS>وp�#���?�Q��آ�Qs˳���`_���=�/���'\���{�m$��a^�5����Q���Ssjo }��j�����12N2ḙM�^��kE�gč�}a������.�.��Ы����X<�/ŧ��	(��Ri޿�u2|簫)Α��&��<O*F����ˑ�ܚ��;�ӣl���o} *��Ze��VtAq[��+=�~#����R�ô�|q������\���8�X�>uZ˪���rP��q����j���s��Z.��<�? b1.��E����,x}|4�*��2�n����w?Mw�bkj!!�$�����ˀ>c�K�����q��ۃ�3��8M�B�U�^�칧"���E��uQۗ�N��h*���v����&M��a I%��ɶ#G�D32��3$N��e+����xG�������e%�;z�*�WKħ�� �+4tR�Jwx��&����C�=%�D�'AD��L4�9�b�scAF����L--(�f��CQf�D�1�+` �m�B�%O�~�t���O@w����{>��n[@�&��#X����,b����nC3u{B)��(�n�Mc���+�B��M��@��ŷs�h����~}�y�+��9oKC�r\)��5���0�f&x_��?�(�G:�;��B��uI����ȧ�9L�.��ŏ��y��S���~�^��QS��A�5�g�G�2!�IQ2pe��d6!���0�&�[���|�yc~����.�'SEZh\�#X�X%����*�=-E� :Q?|?w���-���ǖ5�s��v��?T)b�ȮSVt#�C (����˾��*�5�T�/S	>�����Y�Q��]�*ۚ��n:��[j×4)�lj/�'��kuG~��̲�4m��$hD��%��C�6.!��l��h�p`�7�;�-P'	�}���A2F��n���h׹M�z|n�ܥ9�n�7E��a�F�O��C�ٛ� �슈��%�9��\]Z#F�G&1����fE��^J�*�[+hC�i?2|����J����1�}�nV���X��*B?�[t��	{��:��.��,���OV�;O�����
��N�ؘ��%�'��|1\�+|���+T]�=�}�=�+��|.ѽ3߿Q�} �^Z�'&g|F�����FDq@Nt�'�ݾu�<�1$��6�Д�/���sI;� ����D^�GM�Xܿ.���� x?����x?L�[�.��=�SE���|�wP6b@�X+u��U\���ʕ`���קB82��JWyW�[L��A��W c���L�k�ݷޯ��I�ռ�7�1��m���C�'T���0�P���[c��q6��N�v������-�<��JU�%5Gg���,ܗ;��-M%v>�y�/�h1}��x��t1 �e��Qqv	>Xi�Ų���tI�t{�ճ@β��8�L�Fpks`A�jk��܃��	�j��� X	�c���Ęƌ˃ů��
F��^>�%u��a��S���E��^a�7Iq*���E�]cB���}�~�������J�nzB�z���zS�u���t��fS�XaU�]J`&'
�1�z�&�
��z�	��.�fUC�5��ƹ�p�Ǘú}����|}y��[h|����K�yh?�V�n�����>��0��Rf#�Y�r%���z�\�����j<]n���A�V )xH��.�Ӛ�gr��M�1q��)��d��PQ
�$�ϔ�D/akb�����rX&72��Zps\ju��5�z���~a^6��Η!���֎J,?5�G��'�� YV��*Gg=�4�p�S =�$������h"̃@t�\j;kJf��ݎx4z���+�(}�Ĵ	��ù*���e�ً�Ug��H��u�����M����{QA���G��Pd�h9�g�gv�~���$g���k4�z��O���E�h����c�$�f��.���8����ؑ���ʑ�
�K�+�n*FG�/���)yq�1�}n��tE���4蹵�0&�����c����E�@	F˪�y��\�dp�=A�x��u	�����>ƕ���5#`�D��V-ɻ���������R�w�4�X$�62@����NKGJjv���3�/	�P����#\�ꬑ4g�j4� 0�R6k:c<^7h9<n��l�(��� "�b�;g^i+�6���:�*s,��y�p?������R���&���pm�Ӏ�GbN���юV6Ӥ"�����FF�VI$T9�X*���w�0��������b��G��%{��x����~/>�k�9�8�%�i�E�$~4@���y!�/�,��'2 �`9<�A[��Le�jĚ�p�0� ��R~�;ɝ@���j��Ua*4�@Hw�#
��G�MC�	�IK<X<��7�#^�&^&w9l@ld]��R��R���f�vk���2�q��x�nB���ZhJ#ź�oj��mUaM��6|O�~
!�f�f�M���ϣ[�֮���?2iUȈ��r�D�aW��7p
�Mm%���� ��
�Q�_�n���J��#-�Q]Y(�\������ ���H[�@u���@������v�'q�U����7����L��f��^�k.U��Dd��D	 "\޹��XL5B�o깎"��"ۥ��F��Z��}��;�W;�B|[�i�w�R�TU�S�?��n�����J:�7�������d�_�)93��Pu㸫����p�����U��9P����ҟ����I�gp��ഐх��|+5�a�����Qe_�^{�����|�Վ�2�r$,@Ce];�JbCs3C�����m�|��D���x�## ��B��i@��?�j�w1�7�����ÿh����t̕i>�Ov�� �簓}iq���v�k�dӾ�e�&��PR+�ną$��V��NBdŝA�S���1.ۛ�gD-8���s���355��]�دF���nL�v�:�`�����b�5)�Y��y���C
�є'q���$=)�ҧ޺�#~�/��a�i�b 8�bA�@�?$����{R�x�I/;ۼ﮼��;V�2. �s����z��_�]��^���Ĺ�(���<H��,2��a	��R� ��N��S��=�[�%�~�u1�g���Bug�x����D��Gn,�P��d��g�,�fA֤�zM�I���d�&�=q����Ud�].p�T�$���v�в>ݪ?4��n�����O���ݓ�ޟ	��S�0��$�7_��٤m!���`�-�=�:���pSy�"j��lTrA�od�#�(I��ML�&�TL�=pP�U�"8u4g���y��yN'�W7tD5�k���/xQ×G:X�$�Oj�c��s����!f*9�S(ʉ��"�X��ߵώ���'Βbk������N3Z��l��!�Y1�Z[�V�2G�Ry�Y��b�UC<��&.+�ػ���Ix�Y}�1�[�JAA)ܣ�t��RW���{-�b{",��y��zE+�:��� I�S8��ED���)S�Ñ���jɐ�md����;�
ʨ�^&٪%!qWn�ui� �~�q��4-7TIa얶��"=�)��X��~�9�U{�tF����e�E0��?�'Q&ҽ�Ǖ�yE�U�!k�x�v��s.#A�����'�1m�%p��r�A��ˌ��j��=}׹֣���j7��k3Hyt�.��b6��T��vE�$�|�O��bOo6�}�U1g��<}�'���!����5��,BI<#�X��wi%�����T	�q$�kֽ�>����,�G�����&x_˥M��ȣ�׍�㡂����\CKb�+3r��Յ|�ao>� z���g�o���>��lG�a���2�pu����,^�gg�.8j��ӆ��h��r��^�7��_l��=�*�^����� ��DSZ�13lC�,����f�?�3��*��Q���"VN -zL�8�a����
�C�]Hx.'s&"uQi���-�f�Uo�Oـg�����+��փ8��Z*x�;14
���c]����Mj�0��=;°���y�U˯,�RnmP�|n*X��,e	������oF���w��A䗈ھ��µ���Wv�j����8^X���S�v���kۼL�+g��m��QY;.XЛ�)�rU�;��G�����WvP�t �)��-O"�$�&�^>J���~NF�`]"]���7)��#�'���,8�Cw�D��{�BE��ݯe?�S����M�1��"pB9ͭ@���㶅�`')@�̤W����pJ�B��e@�=��5bH�M�ڑ{�s^(@�_��%�Ʊ�;��$-)��|9(�}�FV���O����ݗ����{n�Z/m�w�5A^ v�|	���z����Bo�D�qn2I�ʓ�y>,K��葱"�d��6�<��%���Y�E��x�m�b��r����rs~�"�Ӗ#Ⱥ�������x��4�4�տ]<�����5/矨��AZ\�r����P���MP��j�̑�)֟	�-r����%�pO�b�ĩ�ۦR�v���r؞�J�RJ�o�N�v�MmT�b���6"���ù���Y� 1W���#%@Շ��Qg��)g�b?o�IT��k��� ���*qM҅8fpEy)  �<6��璁�]" ��1+���okb/i�$�mg�O���$5��w�������6��A���{��T�w;���C�5'2̩t 󛴜�]��(f�.��!�'��N�AmSgy+^)h�]i��rqRԻhAo�B����o���
��[�7N�5����*%se��(/��ƐΓ�$�r>�s����D�V��Jш�8���M^[hJBb�n��~sp!���=�Y���M�Ԭ�v7��zNh,$6!�d4�^�b͍�@`i������;��/8s�"mI�I��k{�:��l�i���|�J
��
\���l �
&�g�
�򃼹AZ�K�8p����3�Û�:�VQc���l��`���z}k��u.�!� 0t?=�M��
�Ʉ������Jc��R3�<u~v����ۨ�9y����q==n�D�f?�bͽ [�x`�sk�/4�^11| Ӯ	K1N�R�[q+��L�����qH�����J�.:�:�n��q��	�iF�A��K1�g+E�V�<�^$������
��h�D7k=r�d�Ĉ��R(�=���W>����vm@��U���s�.�[J3��?�Ԅ�ݗb*��y!��9|��;�#�j��,dV�g��s ��M�BC��m��EX��-���I�J�i/���{�1vƎZg��R�1�I ��+����,��D���� ��ڔ ���"��10�p���]��a'�T6C�Ӭ�v��Ѫ58[8����`/�Щ\����1�_;5D��x��Ӕ��Ű�C�cH��eC?��}�y&����%lq���#ʤ15AwS�p������a�Q�&���|(֖ʁ(eY���z��8*ˋ#Cl����򩍞C��p��뇑��Y4 1kƜr.���~��YN�r��vet�yh|%��Qc"띅5���m��R#�O��<]�x�'��h?�P'UH��i�5b8�۝�>JA�ѫ`�OLw��U5��c�o�(lC�K�&�.�D���_�G�7Ɐ��c�a����������o�]����ƛ����hf1AY���s2��-��,��!g�D,����,�^������� X��kf�6��M�VTȹ�S��r����=4\�		;9�w"���Rq-�12�n�u�ӽ��.�5�m��
�y�}B����J6�Ҟ��T�V�u;����c��E�%vx ���W@n����yr����k(�T>���!�x�b�wY렀��`U�w5������C9bǊ
�%��?��5�-�\P�vJ�dL,�E�HX�%����v��qb�{��Q*���{�+i���sa���� ��x2��W1�D%
����BH��@�v��h�C��]�*$cp$���v�ꙑ&�Ӑ�oڞX�1������Gj��$��������&�Qe�P����$O<�g:Apq{q�������&������AO�"�n~6�u��\��(g���C�D��@���v��J��Á1�C�~�`[�]�V�_L�hf3�z�e�>��
��2jb�s������������Sx�GcK�'PO�� �
��/7$m;Q� �A�sdC��eQ�=�WTk�7e�n���4ɸd\�ANs�JE�M��Ժ��T"�G�!_��ºx�@6�g�lъ@>���h��-:��PT|
<.����>�&���4,�S��=�N��?�a��0�c����2�����%�b��EM���ݐi9�1�\�RatN�d/�cu_�#@�\Ά�*Ͻ�ff'�z$�/��{��ŏ���SaF�����Ŭa�.�3�[v.�c�Q�n/R�2��-c�7P���g�l�AV2�qv;��:�����{��)q�f�`�{�m6N�{�o�~e%��{;ڦ���y�o��upm�i��5{���Q��I���3D �.����yٿ��O8���T`G��g?c�!>�w���;�%ȗo��4g�)��H�Ѡ�H1�`G�����.��\�H=��[.8���!Hd�/�9,n)�F��}ݏݭ�w��X��9/8CY�]<'� �>.�T��+19#U!���N*Xj�A����]٥�f.r�)u�17�Ñ����dg$��n�M��!���o�N���Mlr��1ߗz!��� 5�hY�>G����hC�sID;3&#k">4"�*8�q�>������*�a�֘Gs�L
o_u�UI�u
$
�<����)9��5_�c��0��P!l�U?��c�w�iZ��.��]���O!l���A�L6u`W��s�t3�ǷV	��$t|�[m�S{������OIL��-"��Yٹ,$t=>	�C>�y��Ɋ�N	�=F�Ǝ��<8}��6�@���Q�#�sw�!���oA��S%,|~|�������������a���
�+�=n%�7�ԏ����p���8�`���E��]-tʚn#�j�}�9ZZ�>����K��`�Y7"���&&�@?-WU��רA�jG�o�0�|w5N���h�+��7���|�S�7��X��>r�>����z��,%�B����?
�/����"��4^�%J���TX�'�������V!�ς� �;Y�uaM�5p&�B �*�n�L��H-`&��i�osO}�D�oQ�E62����J��t��~#1Xr�t�a�n����u��{��Ac.;W�X�������c!��jX�z]���X-�-\%����*������9��c��5(׻��B�`��/?M�p�N�U�+��>��ß�:�\F;��UNSCOkC�� �S]hy(���J ��ۃ&������"���txF���.�I2e�����μ��@OK0_��<��n�dIx���x�;�Rs'������ �Q�>Ϡ�k�L�̂5�x��>����,TG-�ܝ��R�����/���.O��&�v�F�w	Ι[8f�~x�K5���$W?��o?���7ct��H�#}��}��9�h9�_W�;gN2)f��"�	Ѕ�,+|�Ԑ��0˪&��qb�Eomi���J�0T�W�s���zK����٬�o6�RM�P��F���ς�z#S@�ZT��!�&�$�����+�+����)��X�Ơ"�4�����(�Q�1�0�u�
B� �/ ���e��m���?���r eЇb�~5{�%�~�L������xGܯ���]��8�*���̗ �hIv�r�����>程��#��P0[�����9 E(Q�N޳���bT��Ȱ��R��e�m�B��e�&x4�";?7��-�8X��9v��E(X
;�:_Ƒ�\�T#HA^L��~˖�n���Py��f�?�םjW+$�Alԛ�E"�z���Cd���đ��
h.ϓ��K�i)�.�Ʃ	'�6�r`�7/�����6+�d���I���?m0iN(|�ܖE_+��xU2��7Ri�(M(��;�7t&��b��U˄6�i��
r��?ة`�����e&����+�g�GX
���C�D++�U��B+�頎яA�mo�HBYk�`�kܡ�*�H�D�CT�������v?�F#�v�����-�m��������ɳ��~H+�U�F�%�in���z=�_A�6}�O�5Q� ��0<�]}��Ǡ��>9v����5�	�y�^���1}F�����w��v���83ߝ��� `8�hKa�O9E_�*9W��?"!e�m��D:E�(
7����ܽMכ��v���~�L��X��$B>l0夕4L���$ݘ^��7�����[Á6����*x�\)���j�t���7�_@�`�e����~q<��Q�k�-m�>����:�l�+��zr�*����$]��%C�DT�fFz
 �`!,����:L��b�Tx�6�9���M()�
�P�X���?_���J�"�I�sr	���ZC��oFr=̫�f_f�h��Y�4���qC?�6��#{�_��"��T�l*q�XC�D�ا���@ZÄ9OE���4Y���b�,zP�<y��U��ܣ�:+� ����u��Ͼ��Gc�9�Q�ݰ����'gG�.�q��]�8C&���6�5�l��*��v;��m[K:�u;�������^4^勁�t�8��翚b��#�v���FT`@���>��O�"Ři�4?�VSFAOr��F��_��b�M*�ƶу!��%��o�^
�[+���^�JѮ��C@w��ٜ7�#�ܶ�N7ޤM� �cr�H`�"�H	=��oG�M[�$�8��<
bO(
q�F�V�P�|tAu��*�GI�#lz���А��l����ҫ��Y�'m�+7E��J�gc.�\
�(�&t)���Zg�43��U�!�4w�F�ޡG��L��Z*��S@���r�D"lTjw�h����2L�K���K7 b�7m`��ݐ3ު���}w��H�)/�@�^i�`\���L�v2�?/�{Ը6wP�g�ĳ�c��H�w�v����7]F�L����Oƞ�/��ؓ����N����/��h��B��-��]�%	�8�!o��Mv�&�d����L��2�~Q������&�e�ma{�;ϛ.@��O�|��;�	½ᖞ�ť
,󨥝�W�+�����R",�n\�_�rc\�G����N�����o��HMr���W+A�����W��b߂� k��
��{�_}Ϙz��H(6L~�z�1�]d̝�[О�y��f���y��������G���tĉ�^j�?��o�1)e&���Pԩ����%��ν�&���\ *OvTf��{x�90�jєJ�����[$)��{\za���aa4kn$ק��ٱ��+�>���Pv[��O�47����f��(��E�z|����o��_>�@)pS�(�-#��K	�,n��p�)Zق���|�k���"5�V�G�f2F�|o[���`�	�T����LYV>p+[r��iBa���!n�Mb�]tff *��B{�q�^��}Pa��S8��t����ZI����_�j�4��kY������h��t�zi������ұRr1��5�/��}�`��&�ѻWL2Z�8�o���
���B�i���P���&��W��}ϩ��u�8�"�so�1'�g�J
χ&�ۍ���8��=g�ʤ��O�4>�����4���j+��[\cV4'k����!`����O«��b�Ӊ����RnT��ѩ,�/�����-4ܲ&��G�
xk.3�mk�9?�Ś�\D��d��L���߆�ݱ
�0��9Ŕ��=e�@[<��!C�;}�Q�8�v��/���: �P���Q׵��=F�5D$���?�Ǽ��~��EV���{�CN�$ѽo�5�B2�j<����#�����*Y��^�F��gSB�BI�)D@��^��7�\% ����f������Aq/c͉'��o��B�-!��58c}j�y��gw�}��j
��cf꥔µ�����o+c�s�v,P�}��cg�]#ɚ�T!9y�VN6�5iaq<ca�iY�C Rh-��k��=k6`��X�֜�*9��֬T9�2d��'T�A�ﯸG��I�x�uj�Um�h�f��\�a�bK���Y�.�D
�}�R&�Z��'��9�S�����>��-}�s�Je��/�Jh�4���Q�#T-{�~�Y�Ŕ�%}Vd���:����"{���2�X��UW�⵩P_�����
�ڋft��C�
a�}P�&K�1���w�b���A(Pm�-�m��3N	�Ri0ߩ�X�ʴ�j����}��KT�d��Z*(�7}��h�����[�}`҉�w�HVv��O'm$��U���]o��q���6�/�3s��J���v0�2~��ٝ��~��eg��볕�P�A�.�k(���A�,U�81BH����TR����aL2�e_��t�{�-��8��u����X�K�L���`�ӄt������9R�ٿR2mq�(+�^ʐ�j�ZW�l?Y�Ȇp��fa2�n'˔X�L��'x
D(ss�|]�#�W���擪�a��~oy7������gh����G®�LW�N�0�E)��S��|B�h�E��##�RZ�m�y��-W(�M���X�Z�*����.w�K�4B3��>��ez�S4�~HD�ӱ���8j�+ )���w�&�$L�j<1Clq��_�Wh����M� )WjN�:�R흊���l(��Ʉ0�-�)�F�,Q(�p0���v@�$l�sS��i��U�������Zr��3(�G��۩��v'aBM�+����zn?�K^,Z(d�F�&�>oBl
�B�u>0N��G�'k�ؿ���>�@%Vk�3TzX^������܀�����;�p����m�j�u4�c
E	8g��<����LQv���@z��?/���͡�4�aW%��I��߼]���yx����鴚 6��XW���<�e�>��vw�wO��w��J5ʺ�B���W*��ۦ��l�_R�ų��+Yf�c ��-��
��͛�C��N�ĸ&��iiH�2V����C3Rd�6
��];z�K�O 0���)EkD!�'E%��d%����ȣ�(��/GԚL���@���#M�����R�V[D���j��γ'��w���N�0�'O�n<¯^�I6���a���&ˡ������<�niT��[�����%!<a�0�1k2YKtF�t^bh�[c�h�EGũ*o&֢H����$�]�JH{���/���l�ӗY�������zfGLYןk�{�Sڀ���t��)�L,�`��uz�uw6��?�������@�����~%��@�8 �� �ܪ�~��g���huE��1���8���*��)�&>�m�9�nÛ�h���~�Q�(�����ߨ�k(\����q )n%dNNgcL���i���1�X�5�h���ى7�v�X�53�
b'?�\�.C���`7$&�)!���	] ��K�3�b�$�U��!4���n���7�C����qu�Ӆ�E͗�.y�H����'��O�_(� �D��U��⃆��A�� Xޮ�0Ǆ�HTj=.ygM��l�7��1��	3�ǝv��H��
��ïCT<�K��F����M����T����O'6xsu��s�1ҏݓZ�C���rkؠ�{�F��m#�nC5W��5�(���@����(n�=W���z8�V���	ë��:��/����M��@�vr�4�!�t�d����P�^�^����A��IJ^���*�����ԧ����'����U?q���$*�+G�m��؀�6cw�q*�ܛ��K,�B�xH�{�?��I���MT(�=��c��(AO �<g�}\�Wd]&~���m>�W7i�'>��|�~f��^�,�21y�w�����6�>=�@� R�Ax���:�~��{&wy����fR��F��1�p�	
��\K��LtcU��u�a�	s�	a�j�o�m�zB#�s��"�Ν�|�jr�z���4�'59�����=/#V�U"urA!�6����[J�I^t�F^M?�Si_������Գ=o��E|���%�h��
�H�����;��?��1�.�x�IceCݨ��^%���p��
�9���Wy�a�/)R�Ǩ��t6��9�Q��m�׻�� �q��^�M'1��"67�oT�$aJɽ ?��O4AO����%�QZ6HP%@Ec�����:b��J��������q�y5�=3�_r��fUxf����@���i���<�c��M����?�Af+p�j����-`��'c5V�T� ���`^=���6>B�0�#�[�iյ��wl)��z~m
��MA!����ˏ��3�Jd�h�.�A�1'�j4�8�BSa,l�wǌ���@�i���ۖ1^��c���E�E[�c��������qC ��ĸ�k��ղ8��l��4'*�#'������I���W��θ�EV�%�:!�kD5!̉u��d��e�g|(\Lۜ��7�4!S6����o�����00��m���$�Ļ�5Ai��A��$6���Ҧ2a�R����D�Ҙ�9������yٰ��2u����{z.�T��a�dD`�������~����$�4�|p��t�p�6����Q�<P�&-�Ú��489�C�F#��|y&����Z����pZ"z3�ʗa��f[���$j1'�f�ע����x�q�U̐N�<1E�r�=�����q���
�U��~�dW�
8O����r�síV,�ș)+k*M�S2  �C��fa�����$��5~����[�Q)ۺ���[6��^_|�hf���8�B�ܪiT�$��T��	�6�V�ǒ����k�+�u�QAx@[c��XA�V��8��*�z8�P�!6�����/p�k��ڍ�O]a|�'p�_�M��EE��Ea4U|����̄ �����ÆI&q)[ߚ��mV�	z�Q��E��;����[,���M����~`�v����l~�5�P����+oD�>O[���nO� C@(Wj�r؏ >V\�8�?����J��M��q�9���"t��:�ܙ�^�?6=q=N�g
D����G��sz1�����I����:U`F�*_0U5����,��::"���1�9��r��a"�����Oz���E�2~F�
\�K����"x��خ��a

	C!<����!:x�P����»�Nn�+����O��Ĭؗ�q��ګ6���B��Q@g-)�t�%}�~��G2+�;�c9f��x5��ly�$���]�B�.�E�Ct��p�c����p-\*΍�oz	����7.i�+����&�H}_���[M3�^�<�@�r:~廟���Dퟛ�Ѫ�5]ɪym��6hz~"z��a[��>�qlG�����=x�w3�-�]��`ҭ�����P�V琭>��I��M�];j��������ݮ�q�ӯ��5�h�1��\��9�i�8݆;��(9T�Y��wE��[ꥯI����X/����Z�����x���
��r��W�UJ�O�#˚���1lW}�Bl���򠸊BL�B1��t���
V%K��.�ݺG�ű1�� |��	t�&��'ݧ����EɎ)��J<itj;[�"	E�ۇ_��cc�f���}��mO�PZ���t2���;�����vd7��¬/l[O���)j]�3,����e�m��޻��\��� ��-�q?ɹ��'>���b�Ec�	/Ǥ��a�j���`$|F��L�B�_[�����fFV����lXn�%�|��:8�&MlE[��Z#^��*4�c�=��.e��L�9�Ӧ�0ݮ.���pb��̐����	GٱH2�>�^zY<��v� RЪ
��;�#X�pz�}\}����g�p	�6�9[�,մ��$�\o\�������«�~jy�5\�tʈ[S�������r�G�\���9B����X �dջ"��� v|�3�^/��V�`x�C_�;M=E�34Ri=�)��/`����r���=�`%�#$��2��v}�!$%Q������*FH@�9e�a�Ab<�?6yz!be|�:�g�����LǸd�p1�M����X�לKRVܿz��˫&u�7�3e�G���H5���� ��(�,S��(��V�]�dk{b$�6'}�����wpm9�.[�Ax��uW�"l�lD�R%�z��^��P9��2z�V��X�M���A�L���uZ: ���	QJ�C�{*����V��d~x3t�G�~]6��;ߦJ������5��*zi!�V��\b#g�!OK)"�-����Z̝f�v̵���29�X�'@�M+�	�k�=4�^��Hy��1�����編c�	QB�w�#���L�z\��n��ёc&i�0OԊ���Bd�G{,�ſ���	����lx����.R-ZJ]���+�񶵝3�P6��}�̜]fLGP��~��-�#�R��>�'~y(��+A�'�51�RbÑ���˰�2��{�J��1$+���V�U:U�}��R��w��k��`�9a���sA��`��H��QV��e�i���P�^q�<���޶_�]2�����
c`�a��(���e}�+�h���d�J������>����6��e����~�L/8 ٜ����A��Y��@��7�6��x:S|�/��?T�KFH�v����=I��~$�^�'2n��y���_1t�*ÚR�����a�C������a �����|���H��/�˺i[-��>[��:���1j�ޝ��7�Y�t$���M�Hii!�xdk�A���h����Z.Aө�-_�Y��d�0��������'��� �pH�R|f��M�T]��B���X���O�"���|&v��V۟�p�l��d4��	�u��5z��<ô&Jp�Vc0Aͷ���s����xp�H���{��c��[�H�pU!��A_����!���eI�Z��Ϋ�#�b�/Y�K;rʝ�Z?iW��yKc�LQ�%-\%魞�6~{�g�G���/��X�a������|Q���Zx��:%�]��()'���Y������F*\�~�F�{���l,e,+�ݣ�G��'���o.@����d/Q���zТw'���w�ʱ��-�2��v�kj����Hc�}�^W�Pjd���Z����]���f��;��Z�-��bhy�i�/8�h��
I�r�A#�D��L�!m��.�>�5�{�<uE�˓j�
ؽ{Q�Bq���[��J��,���@X���s�M8��X�C=Q�AV6`&	�x�n��
�����*H�@^ƗPgl��Ǜ*�Z�����1O�-u�Q��i���Eo�����0����o�H��V�%�78�!Q����,�<+�GM��S��U2s�=z��e��PF�(1wN0�X�5Q�&e�\:�M|��n<����?%B>2B#[O�j���8��w��Yz�.��)���]#��A���"�̅;}���n\���Bs�!S�5� @2+t[n/����c�I=�O�_����J�-�|h��%�7�4�&�H���p'@ �Y+���=�h��W��T���d�ȯnpA}�jp?]�\l�g>���$eʝ5�M;�$3�s$���lg��m >r�d���͎W|=ދ�+�u�?^=��7O�:��J,99�#�<��}�Y���f!fK�/���롂��B1�}J�ҸT�ԍbՕ��nKC�e��i:��G#�
���֦��ٟ�R���?���R�B�Jf&�,��r+a�u�׸j�ƿ���\�֮��{Mk��~N���_E�O,4g��5��n��!I[�:�Կ��B5p}u�WrX�pT�F�M�_�h/M�Z�i����K��u4\8m}����aF��1�@�[�U������ktY�H��5ħtG�{���	���K���.x�x���V(V�{{Y-,IQ !�}�^ܑ�`/�5���l�4��2z�\-/�>��a�
A�z�m�ɮs$*�E�M�,G6-���0�����Q������QqiRCCiGQ~���lw��r���y0m���2<;�I���q�f'����[���l�0!Ժ�&M�����0���*��m��,�ٙ�٥x�Ŭ��H����w7O��]ҹ���#;�J�ύSܯ�`�ǡ�c�'����&���ǜ� Bl�ƲC@���7�<�g[����H@�֢$��W ���K8S�"�Z�����Fb��o�L{�ʴ�F6B�C�
�Ǩ�^�ǎ��8��l��[js(��'2����yW�jq���e��Kg�u��z��V\	S`����cL)�؆�>M��,5Y��o?<e�6ݍk��bpx�Ƌ=3�c���q��'�W��(GRг>��c5O$q���ɬ�R8�h�r���Ӟ�E,��rt�;<آV.�4KA����������#�0�˿�x�+׵ U�����\�`؜��''�8+�;\�Z����oyO�
[�⎉�i����/J�Q��ԁ%����$z(7����͉���LQ���޵8+����M�����3�!�&=�bJ���&t�M���
�uշ��AT��p�ON��,y�LP�2���N����I�@�P��yX���kH$�5� t'X��B�H�.F`��L�\�C�����W�#�����ڬo�N3�@-�{�!���?��!��[>�Q��x�ٕ1��(W�{�z���>�JV�9W�̇�z��z���Ѷ��-����cglP�� ��ea������VF�{ѷ�,�D>暯K\�RekL�ң�fv��,Yi)B9�ܙ��J����Oȉ���~�3��ſ���u��sl��h
�^$���!g�눵}���i L6�����C�&���uop��iW���,���S���y['��p����9���+i2pL�t��k\��v�x�����Ȇ<P%��x�S7�l�m7XĘn��94ݏB���l��Yh�u�/M���K�Pm��!ԗ���s�[t��tu84A�zÃ�P8�N!�W̾w(/,T������Qc��#�I���5�VyF9|�p��^I�^���hL�۾�]�'�A���ʖ��NUW����W�x�V���wҠ������nA#�m�g|����ݨ�rV�ZG�&R�X��}�j8�5�33ੲ����G��_k�2޷�����:�k�������o.6�(z�>�-cf-� �7~���B���yX�^�*+�o�p��L����R�Z�
 �����A�S?J|fu 5���Z��춊A������Xx���
��xۓR�x��pFAݯ�Q���z2�O�c6���XU��//=a�%�wj~Ɗ��\'���#�'�^,}8/���"3�%F�Fb��u���$&g�t�����b�je;��Gb���O?L�2��'i�]lG2�_�,O�r�U���V�TM����$JDJ ��T_VAĢ����U��բp�WhHy-�vtI��n��rp�T=��ի@��ʻ
�}*��ްL|�e�3�y'I�>	�������[k�D��D�Ru)�Ɲ��\&u�GEÕ���~H��1��]&0fX���'��P�6�]y>���C�Z�i��	'�������g�m��^�=�[��M�9q�e,��݈��w�gg��\��<�=�?I��e@e��*�¾>������%�,2�0�hj�bTz�fk����7
�YK��y 0��0N\��~mʎ�?P��8nt�!�|���6X�-l���W��u���Q�;�Ԍ��=��o��f���ڟ�hX���sC�LXM�K۞0�#-�<U(<�k½҆��`}G�i�k���'t�����X�����¢o[Y��V��+��ơ)W����<�y� \�J<�9��j��@ʟ�g�^�Ug���&����G��r]�(�`W��B�~��<7P������M���Q��(k�@�$��2OJ.X�O��F�G���*_ �K����k�w:�
�R����|�W\��QI������j��3UW���|�j\��GG����M�	��
WD����:ob�=m=J�����.k>+Ȁ���IU?��@h����C����s|,e��I[�9���G6���Vs���]ǣ�Ft}\O>k��AR�n���3n���GZ�M�3ו} R�ͩ��v�/����s��v�7䉝>$�����@��P��x�)�$Li����+���N�'��	��ۃ����/��զc*>������H#|���g]6)P�f���5���yJ|�4c��QC���<cv�K�{,��\V��E�]�v6%����5�������=+}��f���Ҩ��oG�yo�9f��l���/�P�(����IT�㞶�G��͑E��ﳲ�4�ؔl��a�ֲk\Uc� �foCN��	�q�u�E-ey��<(���On˭8�>�<��F=�p+�i�\s������u��������C�4.	[ǯS�����l�U���2$^>?��԰�ZM�/�ҲLi�ݐ������( _�� J��{�ȗ�ux�Z�=(��s�2������0n��	���O�*;I���\�ZR�/L��Nk��^�l���ɠ��M�E�\̈́�ğ=:��+s[�fŨL.`+�I��:�+�Ke���h����=uS^OKYȏ��V���Q62^��.of\������V�������Lyx���/q%�B���Ǒ�AÀF�B���~<��XwDس�]z�Y�4�PWwV���5�6C�L%'_/��N?.�w����Jş��%e�B�;=���L����~�P
�����%:8�2����9�+!�'7�bӛ�/x+3^j�B�V��Ӭ�&��I{�C���{���]rL�d�)�T�RC��Yl���R���T�7A�>G��-�S�� ���,О�k[d�l��̄4CWK�����b���bI�pP��ꌪxI��|����צ����,�:��i~��P}��ٙ����,����@,��@Lg�3ɕj(Zd����[Rv�h�w�r#����ɕ�i���C[͌t({c��AP 9��	@\0�� :���X�)s�c�殗�GC���#;�Q���H&����N;`�'^9�4��>CKH��3L̙��xf��P��]f�����L@4S,�Y߇� Q*�3�W��՟��R�������ƚ��{B��l�X'F �<X�.�(9��X@��}�$Ы,Y
V�����a$��V��VzҌǁ>)o�Q��x�h�p�T��2C	��%h�'ӎF�b���:E��eP�V���>���x��ǰ��{.�A��).\KBs�d׷��;ԌK��C�ݘ�e��w�Y��{L[7ɚj^�1�{�ل��Z�($�ퟞ���<=�u����-,e��o�&z��T`��1�t�t�h���Rэ��ڷ[z�kH3�r�6���g�����������uv�Ё��q�fs�3��L6����e�1�ռ�f��
;T����<��;Ur�9�د�6lʐdjފ�����W�n�yW��[�Qѣ�St�V�C7�]��Ov�(s*�=c�uJ���	�=��O�FI�٢m�q��X��*-�uAe�"V�fȆ��4F�3�&������S�a��4<X�~���A3ҿ�H�8���w��ud���k���"�[��� �3u�G(
!L�i�w6�V>��l p�O��4��W���|�|@h��>�kM{M(���]�5;�?���հ�2eQ|Ӓ� �Pؗ��O->���<=���Rc{�F�.k�ٴ+ܠcTfAÝ
�z�����I��賖����6���	.�ul��
[<T�e|Ę�#L9dmU���b�h �m�\�������T���#�)3[b�.�s���q�$�T�����,sB�(d��bG�����հ4��3a	M��6�.���QծAbomİ��uP��$a7�r%�0�,04n7����(�V��pFJ�⺷�O<������c���Ȳ�X]�*=dNƲ�CU��9"I<�wUm��M�glWW� �Z�,���de���փ��w�]���!.����0���;�8<��lU��h$P�>�S��bד�6LԲ��]"��I@�[�umC>kA\�q���1��`���*^���p�"����5ܼ0B=����C����:����8�RkE�ߦ��%��at�=vD:vͬ�t�͕��h��J�a�s9��<\3��N�06}Я0#T �g��^7���gG>��.�Q~�ւ�OM�Z-v�4b^�l�b��y����d�c�'FC� ��&���VQ=BFFR�Ӑ0@��=~q)}�f�0Z^}sO$6��W$�t	M��C@�v�D��E�V�:d�b/�6����T������1��2DPvHa�qK+ؗ%,��� hg�b��h;$��0r˩�騝0�����pf�]�Z������4�r ������ # �H~��(����� G�� �+NM��E�J&>nf�lI�Pl>�h���E4��8��ǐ\��g��q!�_P���U ���w�f$fz����e��p�)�1�,N�G��>y��=^\?[wU�m��7�\	�]��	����"L:ea��)d��ƛ��!��WA,=G�bU�M��XH7[�*��KJ��Z�uF�5G�����E�n;��jx�(L�,,��|�%]�,� ����ٲ3�7�^{��II��-�vWeH.>\��9��]9̀�f���)����'���)�E��`���7 �ቕPfI�[G* �1+o�S�� �s�д����F�y;�%?iD�✌A����U���GWu	��UE���;	�p6ͪK_kyR�".�|J?~���s��B�0��J�-J.t�9\�)͸�����!����<���9;@t����mx�H�$�:�=ր�y�Eb�>�]���e<��Ȃ{Az�P[�P  u��*Td��Kr^��K��� 0l�����"�Q��|OH����e7�֘!����7���� ��iZ��<��s z.�*37ZW��@�EͶ�:�֌�p[��E�L~L���D���WAi]�R��Va��>�s>�&��G<ҥq���˱!Ҷ���e��̰bRlZ������X����iӸ�[��D��0�����������Ά���¾�7��O �)>ƪ�׫o�D�I�v5T��ctT��Xn�-�)����U�1�ǔ+���7�&&���0j��ܩQ�Ô�g��_q���|I��� !�b8�o	�&|�t�15��4������CJ��Y�������Q�o���p������*F !�]-��2�e��T�4�/��o]pU��M�S��Os2i�F����*���ppQ��w`4�'��W�-���P����$R��շ�G d@��nj�IÔ�2�ҟ�0%���e`�%cU4�6N�%�J�W$;ˬٸYNmמ��l9��祍����C$��IX���]���!$n�'kF[�Of�?v���E��\F�Ǜ�}�M���D�S1����
iѼ��]D�\}ȃs���w/|��D�=V�hE�����o��y�@��P7���mqkŽ��I��;DĞ�>�ɟ#�����$s=�?I#����}M�6[���T/B��)���.?��&�T����L�����LV�v���y��Yؔ��OcԬ�j�k��ز����W#�L)�.�X��ax��Y���+��n�9�O� ��Ϊ���v�����w�{|�ΡLj<$���R}���O�e�<Ќ�[Z���mf���UL����sA�(><�3��;�e�6�`N�4+���/Q��/�|��j��$�n��#��?\�(l�Q��$�ӪH��bS��h<Z^6�OYq6�t��
{�6j�a6��#+����߰ѵ�����F2�t\��ʵT���<�Q9��6Y3'Ǩy���29�������� �7�q�U;�J�`� w�čB�_���0c���$p>`�_ѐY`����a�1f��� ;Qq:~ƫE|z&ɍ��K\��#�U�j���D����YF�x��H��C��H�{.���N��X-D�A^g���D񚧆#�$�r:�;K��D	wH��D��
6����E����N��D��yx;��]^��f�``ĶW�yרG��������I'=ł�fS����.�˶��(&)$; ��4�p�C���S�*���.9\ڰ��dC��a��z����df�j����}�5���3� âRu�����-rZtr����G��@f��̦vԸ]��[[i����}�!��x:���}ׯ(��[ܧS��|�&z�ģվ�[D�*ih��N�A�!A�Cj���Q���]i6�j� d��X�<��o?a�*��.�w���c�؏p��u��s	�z�R��Y�1�����4�6�!0�a>�ŚXu;��.U���r��4�0�s":eۖ�GOwc��vX�K>}^cL�.����i���A�vC�*��ͽ�����95���!��1G����f~��XXw��9���m�I;S�P�X����):j6�]b��M��W��r��W�H�P�̢
o���`��z"$`�ߨp%X�'����2A+�~����mǒ_�&�y,�������Á��23�>�T5m�N����Oؿ��H�?��������avO��n(���`gk��Wa'��:�_In�4wp�.]�?�����D���OUEBBmݓ��t���b��E�	ӽJ4��Q2�8%;�  �^R�Ls3��c��MQ=>����v;���؝1�i���m)�_7�'���PW��0���FP��ΰh'�����N}�'zF�����5��F-���7�Ǫb�Gă�4���M5�a���M6]Ǔ����+�sa}���"p����(���0?��
~r�`�lѽ��〗�P�,��'YU���Cu��U����޶[D�V��Y��#�O���pc��b�EeB�r��sb����hP�.U�3[� z��n-���?������]�ht�������k���'�@m=���s�1��4=<���HO=�!I��_!Y���Y���Yfe��8�[t̈"��G�~�����M�0��s�l�񊲴��׍[+�Åa�jD�� U����2'�w�	Tw$���kC<_O� �N�]����}/�6qT�y��)�m�~zt���j
�m����:�h�r0,s'��I:C�&�	P��b?*�🋹͇$k"���J3�/���05�(�gӄ�/�t�vg�<~��5��;�,�δj$��z�"����b>&	�_�^f�𠹞?��H�,?�f\���,�Eb���o�Q3e���|�8�3�o�dP0(�`&���.�xw������w�IY~�8�Y=�����Q�|��~���"�@�*�X\������	S��j�QRJ�Έ>m��f�I�x�й��QL[�%|�f����}���`�O}�����B�um6��)��U�!����Rh�f��9��}��MH�/�υգ �o*6]�#&�D;-<]23ծ>P�ň�x,&]1'IP��h��U١��!�or>��xk�#if�mm��Qrj04.�s�����)	��7��x��)z�)�S�6��M`����j�H�v�eT�Ұ"9ptلA���i��<]Ũ�h�G��1f��qw�m=���'c�m&�X���-(�fT�@���w��s�\�Y���l������\;�E�T1*exd"�
e���	�<(�')+���gW�3l{gj��`��	���`��=J� W{��4Xf���>c`�j�G���8+���?��u9J5j/��x��Z��,�)Z��2G6���,�H!>\[�}?8��U
�}gS�V�ޓEt��_ �cס��5;�gň����ƛ�?��ә����I�RT�c@��"��~�/���"&��jd���U؆��|�4�/>�5��٤���5K�c˽O���	BU��(8B��L�V��\�c/��W��sH"iRd^�I�@ѭ��/��?�2;��3��7%�ֱF� ��<�-�ODíC�'Ek3�&����a�t�Xnb5��Ŗ�^��C�T])qhn�+"�M�a@��'��`*n�U�K"^;NJ.6���7�f�(<=r=���ɢǌƹ����K�g!�h��p�t`�sk��ƌקS�?�S��#�Rov���Wc����*�uNww<�����'�u��I��	��n��9#� �C~��d�%���M�[��˃6��M�r���n����4$șY�%�y�$%wK��y��v»�x҅�FyO�{��)��h�Hi�����/҇O��%���~�����l�+Ọ̑����GkXV�ۅ��f��~B��x�b�Y�����	��W'YHY�DUSs��A8�x��Ms&��� 9�Ɖn��d��Ӗ���f���+�ulK�#q�LY��4���-��w��P|����U��547K9����L(ݼً�3ɿ���Or�p���34�G64>��?�����|���<f�5ʭ�e�W%��I�!@l격O!O59��_֋T�]]?��%aR���&�U�P�c�i�%�2��R(�ޯ�}�|'A3 @��f�aIs9ƀ�ȱ�v?8
�7�WJ��:���'0"�-�e�����p��D=�*��<�?P8msj`��b"�!9*�>P�8Q�z�{6��&�Z�H��:���I�Ƭee�<��~��h�?ej�IM�"!p�������4cg$^$�ȅ��<칬0||^���@���k��י�/Zig��R�b$�s��^l�m�X���#ˊ�xS��V'jh���&+|:�~� ���a�Q,|q��Mr�<��pq�:ς/:�[��9���:d���v�<�����7(hs�k�Z!���Z]�W@[�Wۛ�z?�f���3�a�� � ��]�+�:�my��wmIR�.yƮ�s�t���
�á��|�PR�}6,UD͐]��{�t����S3��ɚL�
�ƍ44Q}��Sf�;�fvvLɫt=�����o�w�;.���T��y$(ye�(h��4��b��G{�!��)IlA��w=�s� v�zA�b�	5�:ב�hclt����1 �1e�3F~���N��&C��s���U�+�6��~��`��<g�RFs>���Y��/��&K L^����}��9�#_���Á�Vƍ;�0�O��>�'��!4��6�q7�'�3ZZ�J�ԔzT	x���Y*�ZҺׯ �T:՞}g-g=�]�7��uAr!UC�W놤
�l�ε$�:G�5�t��c
"���ې|��Π���Z6�����
{R�@k���������۷�ĸdC^c9/�7��px��q�:0$�-{m�£�=hs��L*`�G��7�Й���lF��o\ά_�N�`�ڤ��|�^A���s�^�5|6E����ډ[-
�:���8W��Eg��mM���蜭� �8&�{Ct�w�n��/��%6���1����\]Clu�a��m������
<�=_ys<)<��Bm;U˒٣�]ƅ� :���Q��4�^�:�a0���~�B�lN�&�v�wP����P�Ei}@��|� �+K���]r����8���b��vޘ�*��2-;$�hK�z��(=�����S�oi�����=�o����e���079��=o<�E_F�0_UVܾ�yd�M�����|�J-�Q��z��(��B�^z}�\��-�,X��ݫ
�ZJ�rE���6\Cf�ŭ|17�US}"�V��Q�u�eɫ�Yakތu��J 6�U��'$3��H}��vl�������GJ-ɜDp�17�.�ģ[����d{��H(�����-���$Rs0b˦ki[�����B�7vy��LL���X�}�F2�K0i,I�\썎�~��Cv��99�Ut�ڇ��0hH��[�p	�'O׆�ؑ<M{��0�`�k�M�E5t�^<��̖�(Bʥ�6�
��D
�K�hv�=�7����eJ�b!ZM>��f�W{#���NC(3 ��^�^:���(��؄R�|O��q�5 j�M�2 ����h	�t��e$ٹߴ�P�'� ؐ��	�y�߂�s�WLa,g��5��()r��{���1s��P�����(n�17պo0U?sh� �$:S��}Kx<�#�����c�����(k��c��rZt ϛ�P5*f|��O� }�⾿��}"W�K�ߒ�j?w$��� ?�tx�JO���)�<����g��1�'��I6S������O��-t���P�9�`�����&��<	��]�`�������N�Fex�Nu�eO7��|"��]�iM�2pJ0�`�q��ӰY��T�~��)� �L�ӱ c��!��7�oQ�e�=d���@�+��?:1���Qp�{xh0���AP�,}�P<$�I)Rp|-�X�O9>�cy��&�	���Gt��~ZPgIҰ9�+�62�.���b����|-ƈ��Tba��r�R�3qUzvA��U�E�9�,��g�-FD{��.����%���] ����A�Sՠ"�y������ï#���ږ`�@c_������O�����p��|�6ӯ��P<�tp!����?�^�un;� ��M�/��a⫸S���eI�<a�ʷU� ��̕�F	yh�M��5���`$@sDM�7Jǖ-��G�Kt0���H��ֆU�[������7��N_;٨-�pM��!�Y�1^���Jhb��k(��U�mlEN�%0�_k���E�%\�sH��։7�3�/x� ,Rw"e�v��6�Sk�1'�Ӕ���!�Cv�m|x2�t'����|���sJ��ʚ~�G�X<�'Hp�k�P����{��6&LB�R�,9��?�ݚ����n�$(�Q{��,~,rW���4���������A�L��گ�D�j�_��Pٱ �7����{7xl�gA��9zcW���SeB![YK�nW���=`(2�K��sr��_��܇b}�1����xY�dj�U���:��R��փ�'1�X!��t���v/D��5�����,��ǿX^�IZ}�Pr�N|��F`W��Ng�%<�d�UṎFٍ�s��o|��>,/둛�h�%1[�����zb�Z#$RF`���}�X�yR�?PR��,�U�X~M
�/Ą(Q��dlA�nh��K���(B ��(�Y��p1��B.�_�o�*dL�;�M
G�ڱ�'>�-?�F��p�g]�Ro�rMj��V�]ڃG�͛w`��ga��/XS�p�x�O^4��QR����r��jF`���*_������ˊ�tb�8��&	ǥ&�n+Rk�%R(�s�f����M�G[��X���,d�)y��E�knN��J���&]�"���!�0�;Ģ�.���n	i���$������t<����7�!N��=/�Z��2Ҝ!"���~�Zfs55���4�*�N�1<��ȣ��גZF~ �Qz_��9$/SY-j?ȱ�I��9l>ow��0�U
��5��-'SQ>��{��V"�����g������ 0}���ҧ���[D����:���&�,�^P���-=K�8�Ֆ�w����pp���)�U(�S^����|藤�N��s�֔`%
螷K�{�P��B��z.�B?��챳~��7jQ{eRiޢm���:�ղnܛ!cNەT>!���|�ެ�zl@����X�D��h/�}�x�Wp���&�{8��_�I��cpę�ڹ�P�^���|�C�k��v���PP,���]��Rr%�UAp�$�S:I��
t��(-�a@2k()T��uwF䵸L��݌�/��a�������W��%�s��+x{�G
���+�r��ic�ˮ�U�M��g���@��G޸�%` �_&\Ȉ�*�\9N|�k���H������v���$3��ٌ_�a뻶��D�����/"��Vd�%E�r���^�Swן��w͏35`w{!�Y8���-~?J�O�T��HȆ�γf>��<ȱ�AѶ0'��aJ����e�v�M��e��B!�Xۥ�k�g]���޵3Ep��-��ޅ]��*��*����2���p_�)>t<�]J�Y '�[���1�����޿/��"F�$��#�թ؁�r���.`H�#�c���@���~��g?���,����nd-E 5"�F�C�x9���o��j����إǛ��K�h�y%�6�>A�%7+���*�O��ÆO��8:��l Р�,��W��~#��eZ�_7X�UC�8��V��l5R9@n�4��';%�פ�O.�zA���'K�-���~|��-R��Q�R*�UKdv8?p��΁�o}^̾�%d��K���6\���ڦWӼ�2Ol��%��#�p�����r�h��y��mcIԏt>/AC��a�)ώ��E�Ψ�i4�]������
Y���+��o���b��c/�ߢ/D����㬧 �B
���S��/k�ǝ}q``F�#4h��a���vp~��r���T�
���x␹G����Ӕb�խ�T����*x[����3SEUV�W07!����pT�����b��y�S��S��4bI��M-�js_�� 
�#d�,V���C���g� Fnt�=*� ��͹�t>���$6#,���(ۤvH�3UYL�9�~����M�����`��}��.al��(G�}�#	d��Ĉ\�hC��b|(%��6R��~!�J����^���o�����z�=�Si>c��J݃4D؂45s$C
�v�̍�Ng����P1�V���L�d��T�ɴ�`@��r�?%m��'������<\� N y\��ω0!Ǡ��0��њ�i:�Ȕ�,@m��y�1����wP��3���-��Q񽣓������mWY	�@,v<W����5�*�������Edӹ���
k��8�5�uO�)�Z����0�I�R�2����4ȶ�ȓ�5ȁX-L9(S�2�lE�7��a�.)�و��9��|}ܵ�Qk�Y��6Nc���fX�i+��^-�3W��+�{�X�.}�M���g�L=�^�I����U��S��f!�=6�U~�Edp�;U��F�&W��`*b����P�O���鯲��pI�'cz{��c�Yq@�5>���y��H����0y��y\�A �$���p;C�4��yY֘ɖv�rC�<f�q�g<�������O�W��HB�HJ�i��H�N�ܥ��VơGF����k�_�ճd�0��������UG�js��,�*N�����2�w2������!櫖
���D�TA��r����W�C�۟���t`R�o~D�:
f���W���?*-߇�	[�gF����6A�r=&r���[�p�^��w�.ך��ޞ\ep�i�7���"A��-�3�5An����{<�GP�2;DwZ�d���g����w��n~����+2]D�S���B�J�sOkr��*h1/���R��!�1O0Qd��}�D{�=N�|;� �\�<�(O�8X�[�~X�Q�c��g���P��0Sg��ڕ��<(�IZj>:e��qɕe�e�����N|�N���}Ɓ|���@NH�o� �h�[0�^�<*)�-��f]��I�r�x��t#Qr�5��τ�"
��זu���yҬ/j�p�[�����h(J��^��ٱ׼��A);kh)�pc�˥~�_wМ+�*Dt2��u$PW[#��a��b蜐��K�]�^B�S`�s����_� �Uc̧���0��K�6��ؿ�����K���;F��r��JX��E��K[�T{U���S �x��Z�����}�W�i���}�-$���|r� �0LQ��� �5�_K\��������x�iD�K�A�|�4���aT�z �	�˥��	��~Qh秳5-���I)(����|yYQ���G�O����;���q�b5ȼ̨��V��Mц��ۮK9��i-�G�G�],	�t���9FZrxل5���3���V쳎�zᬮ�[p�hy�a[�����T��7:�^�(�ә��v<aZ����pޅ�M�ѽDp.�MđX��=6��[�㰔�I�1�B;��
�Ѽ�ꌨV{����1�0[ ��I�i��c���K䍡�̝�	�Q�?~�������+����� �~�p��h��W���yݿ�������/N k�I�+��<�mU���t�����n�V��n:�N�+�/`ƶ��3�Y>MH	������&V�cTN>O�K%�&W�0�i!��,����t �� 9л,��k��8�p?q���E���0��[S��gn�
���ђ�K�󯚡 ��I}��c�ȼ_y�����Y��l�Zw+"��4��~j��2�R��<�q���e{��=!�rsy<��9���<�a�"�a����O�X����R��}�Z��"���hl��[��$��������?�LS� K�|ҵ;�>x����G��F����S���<g]�TZ�zD'�z%I��Z[��i��5��ezܪ�@i,8�q9{�*k��$�`�StlG���/�z��g���"8�:�.�k:2й)��g*N4(aא�� ���:\��?�g�U�*�n��_$8�"7�׋��Mܗi��Cw ��@���yK~����V��VeY��8o��v<�Њe"�Ũ]?����G-h�|2�h��8�>�H����ޕMl9��ve����]�����CQy$������0A��T$�r|�P�L�	R	o?8�� E��VU�W1.��x�{�Wɇ�=2�����ktP����c%���NC=�<m�.�q���B8���j�.8��]f	�^	/��jML1�HH��M�ոJ�U���:��l3JhĂ�[_��y@��DTwHJ�.��������G����|\���4.+�+��Vq)>�H��C]�,�15�n��5�W}�� �$��gF�h�4��/	��gd؝���ڔ��\����Q���g�s���t8�F��ڱg!�=dADR�ߔ[r�D#v���U�Uc�*�|r�	�Q¾z�l�0ZX�|l�<�&c	T�^�3���J-<��4ܗ��v]N�y5��T ���@��.���r��O(@����\��3��4y�c`���ݞ�#�
eU�7T���!�ڊ���d�I���[�Hw��i�����=k��"�����
^�L?<�V.+�Vtfǅ=O�8aASR��H��[�sI�¢3#]Ӎ��%uꊶ|M	��)��O�P��K�/��'Y���R����X��A�̽N�jٌ;�9ѓDo/f
¢��{зl�3�G\S5��;3Q�X
biX��&	�C��0��?�6k;A�m�T�iJ@}]L2q����|�����O�@�Ƞ��Rb�� �#*��	_���3PsȀ������y@���Y�}����j�G��ch��N	Hfs�[�kʨ��' �>G��"�����z�>��M�߹v�Z������:�/A Oé1�7�t-��*�����03��r���1�*tw���;hB�Z]+�#ft���-�G��k9a�������rW2�ٰ0Ϧ��ȉW��Ʉa�?�]u?*��)hg.I{�sבV }l��3�����)~�pL��]��	1���+v�ōz|_U�j
�����=k�I�#�[k���AcNڰ�������fB8-�S]��Q��x|�U5gڠ�i݀���X��0_|_-4�������<�Mm�~eE��p�9}�A�htu����ߚQ/�r!MN�i������6���3�����	ۜ�g-l��V,a�"�JV���+eY��
t��|�"�"�􀞌Ec�=�K~�e,S#��2���_��2z�|=�S�ű;{>Py��]��t��*�$��g Ҵ��beO실��hj� N�y v/���&4���Ԙ!��	�lU˯3U�tK�-�Q^�j�#�8��<�~qbbW�I.�"�rU�Քd�����;�*z��@�E:�|*��07,�j]idg`��y*�ߏꬹ=�W쪠c�8 ���[T_A��?����[����,�VO��|Wl"�����ú��%���W#g`Q�u��f�!u���͛�ֹP����-R�]/Hy\̞&>�t��>k&��D��癀"�G���4E��	F ħ�Q7SB�=\�&�(e�Q� �����A��O!X�!��w#|� 8��::ź㢂G,aF��}paG�}h)Ȧ&Kj%�����ޤ%Ճ�GSZ�W6b�L��4H{�#�Qr���߅,2�(��Ч�K��⍢Z>Lr�d� ��XM`)�L[wн�JV�%�X����CZ����3ٜ4�m+<����JGH����AW��S��7H-VzNE��F3yL�C���/x)���נ�U.e���t�%2���gz��=&M���T+%J��L0��@L�0����˙	B�|�Z��Q�)�
�k7_�s��y.a\���Y��-ӁH�M�����8VOײ3�XÈr��o�.��]Ff#b@Ve�F�Ci˗����J?�ܣ$�GdTT�q�yQ�����1Ղ��0�qd0�<�B�<>b��C��J!Q�*`߅al��Q�2�8v���}���m�`J��W���b�ɣ��,oe-�G�����QJ��$�`��y!����ПL3�a.I�g��e�sl����/L�S}!��C6G�����6&�ߊ�]�ի�W�����)��=��L��8t ��:J�*N0ľ_�;/7���E�-����Q�036�҇rHW^��������g�5�ŉėe��x�մ�<�����~o�ϝG{�G�Ĳ���#�`���y�<M����d8ޘC�r��aH`���n�g|Z�\Ċ���x%u�Y�V�,�Ey܋;a-�"��g,ܾIiAY�7"�B.��穰 i.��$z��e篡�7*�|��OXg!���30��n�*��5G��񖞝�M�Ʒ)-b�o�z9�S��A�b�w��zD��C}�f�MP����Y���ޮYzYy7U9'܏������N�wJ��g=3P)x+́X��ڶ�~�o&��:8F�����wyf�
�6ڏaNSst�R��9��9�Ұ-D�>���م��$%q�Z��t�sC���a�z���\�ƪ{Ӵl���膱p��O�)\�����UL��
���^�o�ljN`��fD2�:�A	`�p��Eu�v�2�n����ӏ���%']j�1�� i�3�O�'	�&u���pr����"��(RL�m�0.b����G�i�"��A�OKꌖ���Q�C:�I��F2"k��������>�`��0e�,��EG%;L�Tb�<����u�Z���O�ah3]� `�>E� �;B����֐�Lx�H��H�qF�G��O:�򏩢�f�Y���oOG�����hG
[�x}����6�O0����t�|��7w6 7if�~�2һ6 n�qhj$_�5�L�wp�`f�a� �u>�W���I�-�'J�dN㪶J �����G���h��s���7��uk�M�?�jv�ٓi��O���ו����rJ�s�7u��Lc�:�uX�|�i#�<1����z@�	��G&b^���^�s̒H�0߁%��cO;���Z�1�, D}���x38�A���B�xS�Q���!=���m��r��*b��w>���i���ǉ@�^ÃĹlB�/�����2a��"�ـ����%Βyޏk���L$�b�Z��6�������q✔8�e4�a'�R��"�="�=��3��ڣ�f�Q�=և���G��Gb ��GFj�XQ=)��OR-؆��k�O�%=�_�nxK�q�T)�3�|#u�7������ln�c��y��x ߏ�&��2� �K�d��lO1��vZgv��]�u@1�k��=�Z�!Lo��ǥ�'7�Jg��\�b�S�/�@�:Y���N~v�9��Ĝ���8>2���2��p���\^>�M�O�N_� �Q��j�ۂh�À!F�]����$�w-��vx�v7�a��&���.PiуD�Y |�"�0��wE��c��
����\?�{�F!s���t���FQ�#�)���;G����"ԗ쟓� <��R|^Z�=`��hcw�g&׈b'n�p5-�$���@g�b 	���T�����g�]�K@��ͣ��Ш�:p��
Yh�HZ(=cO@v�1�g�ث0KJC5���j�k�}T`�]�!+��z~�E�`Z��q"��$�q�$������c��3���*Ku_��1^[�Vf�԰3.3J4��>�m�
��C�K�����
�$)�����+�}��0�x�d7�O#��!�I�C��j�/��б(J��)9����[�2��04x��FT3W��r�P>��ܑO�/��C�ƛ��	����#P���Q�����=�ƣ��WO����J�7B�	���jDiƣ�L�Ly�p�`���f� �me���?}�#���ʔ�U�Xkb%j#�ڐ��F�����1a�~dO5�dS`�5�s��%��7�dv��ɶ��YQu�NX�iU���� �&�cQ����e)�,�|�$���_Һ�k�=|<�L���C���pj{W]����/$�i��,������������[�l��)A�� ��>�b4]�]�o),I���5�+��U_^���ȸ��I��V_���ߴ���3w�i�2��2�����}����ա��ϥ��-���k�Hf
G�T�w�P\�w&Fj�Iؼ�6�6�/jl��G�p�cE��V��wPM�Xf�VXY���hzJե�-Fg��i���ylA���� ��;*�QS�ĒY��a+1��F[�n��9헙AaW��Rx�!�W7og��^���WE���)'�"��!�W0���:$��)]ކ���x��n�ݺ�k;��tE��ٸ���Z��~P�/�C¸���/�>��̄R1�1>���g�;�y��z�s�ô�SG�����b�ԯy@�
�X_��o� =�>Ȃą!�h�ٱ����rQ�����uNa2I#l�m�v;}5��lTi��VlZ7FB��?��	S���8!D�s������$ٿm�����8��(�]�Qg9�`���{��Y�ϋ}�,N���^J��n$�v�O/ʕ�K@��N%����}��M�$r���͚�{|����˿�CRO3Oh @�7th8m�ky����A� c�5N���,>������~��;��P����"���N�`cU��������m3�N�<wwmY+�j�%r��#K�-~x,���gZ����ec���"�$�0����*��ؖ�#�1`�%�.�N��80�����(�lj��_m�g3O84;���.�F��F�"yĵU�Ƥ��^{}�+�s�t**7��?�I��eYw�5�-B_��E�3��Ԩ�OH�R��[s����f���dvT[��S�l�S�=)p|sH���r���-M�I��H�t���!!�5�F��I��%:v'��s2 ��7i'|�g��w9����Lߚ_Z��K'~ߙ�6Ľ��P�&4@�D<���i͐A��"��L���M��r��wdX�k4�	�P⁻��RDG�߭������/V��X�N�8��b�N9�\5!$L�swG=6�D�O��:�λ�����C���J���R���WE�?{�n�Իt�z�q%�z��?$�����W'3�^��h��oۉ�Y&���8��ǐ��FS�d����k�$�L��<a��Y[h*z5K&�P���;�D�E�[�,r?(�'�KfKY=��t��72P/;�Jgy�M^gC\�H�����NU�¥�8��@��#�)��<�u�u����چ+?W��U�K�?������ӹ�
������w�O�O�&���Rtr�.��訴zL�E�i٬��Q���|�!B7*��Q9�D}C�l�jq1ImZ������Y�^K3�u<Q��'Hef}�p8iuKiڏ�A��:߉���"@�4�d���ᎇ��^"�9I����d/����~�� 1hW��#%#҄OP��t\Ʃ�k�T��H~�	�7����3Tt2��j�qL����5�Eӛ[�/����W���:�ܬ��z�>���;'P�mE���	/��)B�Kp��-�`'�(	�Q�e<"bRU�#��6tJ��J�T�Ԏ*� �aN_�U�(v%�,ђ �Na���O����d��'��pҁc����"��k�py�1|������BD�
���ue�X�#S�b�{L�?�Ik%Z���-������ $«��r(��Ime�?GA�X۹�H �"Z/6��=Sڳ��`fd�̐n�h�=9yg'��WϪj�:U�q0��]q��V�mRPl�tWj�
����N��+n�Z;w���o�p �5q](�zq���6�@�֍�f.����;���M|_Haw���l:� �mƢ�3���-��U������v���zy�@��"�{��-�x9�N�*��B�r�8�h�0�Cֈ��<5S�7�@3kM�,Y���r��.��Ǩ��a�U�hޣZN�=�i�8��/ݑ'��.	AыzNյ�B7��9�Fl�u�Si�D s�0��]޹�mB�����AH	��o���s���X*V��+�.��"�!���?�L#�=]�x�w�^e�
�cv����L��$������������:j�9B�8��4PI�6�f��F��l/e�?�|�inW,�y��7��G_c��>�Uިm*�*�i�}"�X���ȼ"�x����q������q�i����k��:uLR�	�k?�
<�@g�3�3F� %z!�v�+�8�.��vuZ-��582c,Z�[�D�����]�Sy�HZЊ(�#���9+0
�����O`��9�����i!^&Ռ��	7�E,��+��t��w�`~�"���]pONk����a �jM��vD� :YI�<�o���TrDV�� �/ħ���c�y�}�$(2��H�S�S$x�ɰ�8#}ǎ��|#c�
��4��Lw�3tb�2�S���S�DTD�j�Z'�� kw2fb���$�AJ-���ϛ���*��l۴����ɖ�E�}ћw�J9"Ra3OE=��/;�1���7F����`<:Kg:�)��O�����ˑDԺ֥P��*{A��Dg�M�p� 3�M%Fe#ge @�@�&�6�t�7LA�-r��@�<�'E�*9��.�w>*����J�`����Ć�����cr����G�%�l1�eS�I0�W˅�z��5��p�H	Tc={ "�W%�d/n����R�~�o�[Q�/�jFe~t��"C��Zc�����Ln��k���u-O�����
�Ze�+'q\�}��\����%$�؞c�|�jbJ�`xg}�JP[Ŀ���d��1Ȝ? ��ʁ��Mp���X�,����1�����^Y$9��B��@�4�rӁc;�sýɲN�]�&)���:5�i�1�&�|�)�&fn隗����ОE�C�ۆc�p�fbƨ��f��P�/ф`1��&�q�þO9�®��s+���4�`� &��g�� z0�`
:�3$��pF�	ņ �q�߱�����&伛��Y/��5���u������g���_�,�,t�c�ӕ0^9z���{+d���FN���WոӺ�C�[�-�cŜ��s�1C�ȧ�j��D��=c1I�_��d�د�g�&��5�sU�=_�[�c?^����.,���d�:�$y��/��j�Yv��W�nu�7q��Z_��x2�5�Ĩk�,�(�6fFę/R�d��������CO��b�[�P�'���7`�]o�5�E��)���R��lc'�G���ifqPE�	4B�a��]���A���;�iS~�v�C���6��=	���U���t�����m�q�Z�BO�60����2�W�aһԋ��+z����Y�)�]�j;2&��0�3�gq$*Dҥ��;�X_&RV�S�*��n�%>/o;�Q��9 ��?iT����E��vcQI���>Qs٠F�N�8AZQE���[E�/�1ق�Xx���Zà ���t��SA�
�D�PP̬}�{6cf�V���%��E�孥d��|�q'�����VS�g`�Y/>G������:��Ί�z[�2u{�2O�Z��d��u�J����
H�	r�ާ.�����'����Y4��z��:�{��|a߻�[���\�b|�B4L��縸��0�[R�G������j^�Y[���/'-���8,z��*kG�,2������l<�me3�L�ϜE�t]�������7ʹ�@T�2v���\��y°��#!+��;�i\ΟR4S
�V3������9�T����B��� �%���6�R-��Ȣ��6bE麺�"�+D@�� s��Ű�H
�a�p����qB�sg��N}��N�� �L�v�!��%�@���48���
��hc�;���x��������[�yO��t�Xd� Oɍ��G8��O�#���:�D�-�Y��A�+|�+�B/ �.����#�BvI{q�Gt��V��f�ӌ{դ��L'��㚽�f��QW�;�v�I�[f�6�'1����*���+e45o�Ae�M(��1�f(����D󛪎���^*.��t~J)O�b^~�6���-@p3�7ȑ~�{@����6S��m{gY�T�.�X���N
��)�R
�'�����)�Z���F�H�:@�ݬ�������U�tң�p-���BqKUX_E�h;��3��wp�͑��K��y���~�۝s��mA�p�h8)�(A*��i�f`)īyv��=��	�;�'�7�WF��l
/&S_0��A���F�u"���C7�-��u��L�i���'��B�����&�Ea�{�"���õ7f��]R^�P�7b�7�J^4�c���H�g|���8gM� W�s���v#F3eڶ��}���,�� ^�ˇ�B,f`	8DͺŜ",��*��bTa���[E������a�'��Wh)t��X"��Bg�X�H��&�A�fݍ��,,��.m�m!���XԔ�,�_���T�Ff��F{�jl��9���gIȅ��/q\�����H?���p,m�˭���,�T>��[�T�T�e���k�T�-f��+�֛��Wdy�rq�-C�0��/���a��%#�.G�I&��y֏`���DV^�S�Ek#~�wG>����$ݟޅ�i^K���;�j-ҫ)Lf�ꧪ�=��or�����!9��]h啚��$]P���� <�I�/��j$#ܠ�P,\o�@�'P�+�7�f8^r�E�+a#σy���/h���L���7���Y�sʽQ�F:�-+�(#סC��j���z$��d�IQ�5CW���i���4E�ɒ���J$�χ���RW���Y�nQW�'ܘ���w�w�� 1�ߏ�]�Q�@$��8�j�k�A�W��;3�B5��c�6���w�]�� Nj�#$��F��vޢ�]��O�{�F���ގ�^�Ӗ����P��?������Gw�<���	Am�įh�!�=HJ,Qvg��3�L����V#'{!��C��'�I��_��>M���2��	�ʏTx���WZ�,��6�⍉
*��������Y��=t��.S�F�b��I$�s{>������X]F�Q2�jk� &��-%}�<e�h��9f��-�Kq�����t�FH"�ة�;ь����80��i��Ą�O��7��Gح�Rx������7�a�C�Y9Z}4�>�1V��zY,.5��Sg JVg����6X�U|Jk6V�7��(B�ZtpS��X{uQ�H9	AH1 .F��Y�����C��\W��w����9�`���C�ȁ`�o8��,�0�c��U�wޯt�-|\�N�HP>��!��C(�5�*��3�CY���yPi�_e��$�Eo!���<!xv�/�0O�`"��O L=%�!�`��XI�;ҟ�-�1���	��g:io@�J�����%*��\��Y�tRre�H��G�e�,(bvE��9P8��ۨ=�
�X�k��վ+c7I�����Z=�z�g��:�R`XwU���[�ߴs>E#3k��ƶJg�kRqQ=��{m3�#z�cOM�/#X�M�'D��c���МѲo<Ĭ��UD�a�~�ѽ+]�)����L�{�|s��~����9��Ƅp���&Ǌ���ݛ��}��v�gp�Hk���O�����C�$��7��X ��:�O��K�5�=i�%�W�~T��2�>�[�z��c�,��ndoՎm�w�i=�T���B�-�@#�h�]����D��Û�|\�� c�Y]�v�9�mݭ�|:vsK�^� ��Z��B�2�k�`������k�$vw��{�^m�
�"X�=����h��˕����+"��$6�vP�����i��%�� v\ ���AZgǂɘ]St\�`A-��f�qu�����-{��Jy�ry?��!O$���ا��&y�w�桝�E'O)toh����w����_�4V���V�aHz��:�T&��s���2�O];ʝ8 �'ǳW_�q��H�n2�qڶ��R>'E4
��g�m��n�W���`TI�F�֟m��,'#c�L��AC��M�ʟ�r����T�TNr�! �p���K�/Jl���u{�ae������yi0?��	�A�:�A�;�D�Q���]8�����r�nr�-�V5�}j���=ѾwXt�����Mߚ��I���c�-<���	wn1s6Hc��!\#G��2��ҖQ탒�S�\�sf�����m1�Z���sr5��b�c��K�N���.���'ܟ���f��V�ܬXrb����w���r�{G�b!�4u^ēo���h� �ҏk�VӰ.qW��蠆�Y\�wW��v1�$���U	��zIt��\7�%�,�2! V���P4�>��zᱎx�$�|�,-0�\. w��"#�,A8���\�J{�d��a�Zeޤ���~��ow��Å��AvΑ]D��m��W��@m!�����^��՛�O9Q���:�+,�I�ͅv�!̓�QK�6�Z�h���<������{D��y)<��`�#�o�9�|7o��H��5`��K6�L�d��of�c��|���xm'{]�,���z9ayއ��ԭ�b�c$�N�H|RNL�8��k�~#+��F�YM�3�!�z�i������U[T�$4�Z�`��9�����e���HWc���� ��xk�X�M��<݃��s��:��1S�`_r�ˍ��P~��DuΔ_�5x"ai&�2L>��`'��C.��gAxt�q�/�i%t��j9���ݼ'��劙
��߶D�C)��;݊�4h e�ʬ�VD$����X<����3���慿��W41�("��m�TU�T�-�׉��0�I�SbIӶ��Vv���<t�����Yƥ�19�(4�4z���ʇr�Q�%�_G��M�_����(���U��|�f��ұmuw�Z�S��aZ��e���sy[Zδ*e��ao��	k6�WH�<*�W��f���hAP�}��I6|J^��l�-䚬j��W��ؑ*nO�q�[P���,�po�i8���x��49� Xzs�v�dB:���ɕ1|vؿFc ^�~a+>��M�)�H���Y�bLvA�`9��;G07�<Bg�J��c�#|%�L��^�wL�U"�sܠ�ۿ�i�,��E������:tO�e���"Ȇa;����K���3�X�0�<%�	D���7�Z8�"�$�Z�2�ܵF��[�t�ǈ�׼�W�.�)��z���<}N�.5��usB,-jۮ�P��Og��������y�n��N,�f��0��`L���lm�	_G��ݠ ���+H�{J0����h0c@��J
��	�tL_��H��Q��D%^^�VCQ3Q�Q�"���ݛ'Qt�j��<�K��m���^�#,��z��Cw�����Ѿ�!T�A�.���Q�muy�_�����E��a�&�C��w��SĖ����RǨ��*ϳ$+��B>�׫"#Ա�K�\;}G��@T�o�W�loп
�2ѯ�Bv'���J��֦Fvz]>���'Ⱁm�Ò��2W�x�M�N���w�^T��M��|u������L�~Á���x�=�ZY�k�8b�]��Ⱥ���M]��?�t����*c��խt8c��w�HCgY\���S��U��0Қ���)��fk�qы��j?;c֣/���̳��oҖ_�1���;����fi�����4 ��� R;�ta�G_?gJ�>r������̆�j���{��+U��?�V���7��Q�����"��`�-����u9���n��ɾL��/��w>>�VpOI�~�m�����[�z���IU*�w+�r�xQ���%�%�l��:�v����Z���-��K�E$uﭤ��B��8��a���-��ǭ��,/X�>U(B�޸�dTf�L_�r�‗-�Ʊ�
�b�c:��5����*���f��`@nʝ*�vF
�v�(����;�Z5S#�.�[1}r���A����"�D%}'%O�����L�Щ�i��f��-q��Ў�D`]Q7"̧[���j��8�����\"Me"��ܿF�6xI$� �`N��z��Ou�;~\���쓋l)��`G��5X���XMd>\ߴ�-�m&X����P������gY��]P������i���|�D9��� �/����GQs9}�ih4D���_�s�K��b&�s�x���+a�e��HŔ���g����N��:_�2b��שs*�z����q���~,5�R'=MNU3t�>�U�c 0��r��l+���0r�bċr@Vwz��I>ga-�/��Uf��=�cH�"̌pg�5R4���
�U3��%ʎ��I�Tw�j���΃?H[�]�������-��wy8��>ȏf�%�z��<�M�_,�
s�3A��8њ���&���v�W�h��o�Xel�Ҟ�G%����5
%���l6��/�1�E!���7��EU���T����^�~���1$��q�@�V��]���i��5r�-��-�6';-rA��3�+[�^j���/u�7�b�k��1�0?]R%��>�����Bo�{�u,�eNX��hNR�Q����ĺ�@B�hۏN���,t,Us�m���?��$� �ذ�������1N���'9c�'��^Hx�{�n�|^xLx��������8g��z;���N����M�maS�(�	��*����?�??J�~���# B�_���4@��o.{�:�C�l��ct��5;���A	"��n$2{������n�|/��9�?i~���d��eM�k~��ڮ�tSQJLҡ���2tW˓�K8�W,���0,n϶fώ��:6齃���KTZ4�{�]���ƱZB�1�S��;�$y��O���f�ė3�ha��HĽ�����ʍ�+[��1����<����y��a����t����L��#f�yZ��;�y��q��vA����Y�%n�� �W6ޕ���B�SԆH���O7��$)X=�?�7�{�i�8_!Щfp�R�hy�~>�ӆ�����e���]66�8�6����������R� K(Y_
[ܓ�MO^%Ҥ��h�����xI�w�Zm����g�$�&v��2?Ts���񻏸7`�'��d�W�\��g��h2��|Y���)0U��\�aHq�YIW@���}��-d��>�M��x���������?����B�@�<t����N���df�/w�b��QLI_q�-#���Փ^�C�{x������
�Z۶M%g�<)�8 ܞ�Ԭ�������X~�Tn0�VL�3tBZu�B{��EX3FU��y>�*)�KpSHWvr�ڈB���^��G�S���cX��㹞)di���=�h�R)k�;g4OG6���gbf�*��F�O�CT�.�4�+)�:����m�$��Ģ���P�L|�IH^��2���̫�;��QG��n����bB�e;���.��t�����'�{�����%�����H�I9�kF��ܢ�
�|i�9�8\JQ��&�T�J���@K����@��A������z|_oP��>�?���l!w�(?&�<�67D{��WX׽А�x!r��'�9���XY��i����L�P�PN�,G;<6����|����ŮW�g��p<l����ǆ���p� ٚ��/�&T7�ᜱ\US��������(m�i���k�`����.��'���6ս{��|�M��:�$�m�|_�SR��ZqNs|S��"P�%)ol��J�i4O_�hf���4�F^�.��+9��O�&x��6bۇ!��L�+�ۓ�/��1�B�����>�<�8������J��42JT�Ҵ*�������Qj�/--)!�*�����+F
�;�09Y���j�����\vPb;2Ȅ�S�a��w�k�Lm�p��`S�VH��-1(1���0�a����^��IȦ`����c=�v��Kw�9��4��T�!���B<�#L��`�*�j_ک(*7������nU�
;p�!��v���t�(ԟvZq\�ޅ�$��4!���3���/���G��X�#����[�5���t���6~��ԿN�W$�����y�@�&H8�k�h)xH�2e�9/���5|���JJ���ʾ�n ��`ΘlçR���+O�(���V�D�����Ξ��9"xR[�����0�W��Bs*�!����x�y� b{�!DF�x 0	�ME�=�_{�AX��Ʌ�V̉.K<$S����H�@--�������nqv!vM��B�=�{}��~t�j;,���A��}g�'Vg8t+ahPO�wh�6����͈��"�����`�2Ǘ��a�7��-*��T��H���z��ÑJTi+��h܂�0`��)�Q܄���Q��)x�q���KN���6pS����6��F�d3B(T�!+��n�$��c���K{�Xj�5$A�y������D�\t�`�M�;�^����,�6�ȍp9�W]5�m	ʔ�]�*Լ���[�0�) h�p�	�q�l֛��I���թ�C�$��H�B +&�#�.�Nz#n����9�k���y��r^-$����D��)k˖7��Y�N������|����f��T�G��t���9��M;�=̫O�aQ4iy>Eg�GMm��^E�+&��]>��D`�8<�������7x7 �������ݲ��%k��VvN8�ǁY���0�&K@��i���я�!6�~��+��o�X��:B� �֩loV]:�rU�2b��m
���F�H-1���6M"�6/��m�3�8��5�	�^�ێ���D�֓���N���9؉6,1;���-�^
p����4= �7��^�e��%�GUo��:_G0z��*�&��M����IB2�R&��㰯���9�Po'�q.J�c�TU�MA0!���v���y�n������:�L�6b��ִҥ �����n�w�%�28��ΌX;���K4���P��Ql҉�ў�͒��]L`,4+e�3�__g��k.�W����ѽ���<�� ��ՂvxoA���x����Z�B�b�w=�'���b��e5k�m!Uo�Գ����4�
����q����ړ
�*��&�A��,+�0�~� 5W���`���emDM��b� �ƻ	T���0����$[���L� �ι�#0�D6��[��KEk
�x�v�9yT�5.��O^�4;�Ҩ�3���`��X|o�j���;��k駯����*z�es����YAޒ��]� ��ޞk�9��[�s�ّ�L���]Ǎ�Z�gۿɅƛN�����t�����պ|37�yS �o��e�����X�<4��3�H�;j���B����A*F���{�L�1���?sc��2�Ư?<�#�#tAs�c's
�T��O~%螓J-2l�94=�su��`/�g��h�1p�kx��\n�����9JdҝQ��L�/~_��Mei�7~o�3�%�tMzp��<@rrfZ{�e���������Xzg�[?�Ų�XeRc�̄�DĿ�[���ٖ���Z3�H*R�h��}�B%�����Ra���rj��9�F�S�\�W�ŏW��
-��/�B�vӏ�;)�S�w�
{���7)�l��v�X��>X�}���A�C�E~U�e9.=���|�5�������ߔ�㇩�߸��A�&;{��L��(v�8[��1����/Op�j�`鸾�/X�c�ڞry�O@s��!��7-P�A-L��ױ���3h\@k���|�eAv�ߑb=����P9����)9�A��";��Pwd�t=tT��@�0���:���4m���A�l��]�C�v�.^q�!�X� ^-ϧd<�o���v�����:ߚ����Z%Cx9�`eUw���K�V�l2�+_e �	�����y�'�P0 �μr�Z��ϻ��Ҁv�\4�Wn/�k*�a����Ɩ�6��˫�=�h�r���p�<))Z?1�Z?C�lO��{3��2Q5R-i�tYѦ� ����h?�Ҙ�7	�̰��0���v9�jȾ�SP��f<����d�90�r�>�v�����@yM+�h��F�7c�^ΛU�����i��G��aL0>N��F ���]�=,�h��4�+��׿��kzj�����V��0p+��7<~��z"�����}a�h��4\έm���{��%7�D˜��i���G8��eo(�t�@@�>6E]~cd��j�k~�1w`-!x��܍����m���@�eg=�4ac4Jش!�M�e2��Ҷ���To�FT�%�}K���Ua2b�X}]4T�Hn����p�"�q���jF���+���A�d����.��q�5s�;d��h}��g=+��ѩL�+ �T8���?��9�a��N&[���ֲ!�g!��ϓ�s�h�O(�����UD�s}�ɳ���.�+����O�R���h�R�>�� �FQ���nUq1����9\f��Xb�&D2�.��'  ����9�����j��5�\}!\�J���h�܄�t�u�M�~;iguc�.�����QN���)�z�v�0�ތ����tp!Q���sZ\�ZOq��o a�)O�؆��5ui�)��Ei9��4�����0���'�����/p�~幚�+tgo��Z�*�D���L��B�������r��p���G�"9\~È����ˊҤP�K��E��;f�_�w���3�2�B����edO]z�9����H���*�<o����$�n��O�!rw+2���;�� ��ڔe���»����a%L���7�t��'��F9�5T�yK�'0��"�"�n/�t&{bZ�bLN!�C@��o)��DC�{pF�ST��o�`�g��,Lٿ�JA5/� �?p1����*7de�^�Ɩ�یeΨeO�u�ϳ:�cb����E�I�,*Ih'h[\i�����Z���n��:�O��-%�| ��_�hr3LE���3\��N�J-2)��o߬I�;�^��(���q�S�� d�E���)3�CAbH�ϲ	ж�R�\���/U���ǶJ�E"؁ �ҁ
WvF6ܙ�#zR�p������n?��|l�	����j�XHQ)@�:se�¨k��Ik4���y�4�ڄ�k��Ц�-�.R��f�fY�,�Kmd�$ce���t�<��ɤP3����	�"�#D����篣��%s܆/W�\�F��X��vWi�G����ִ�`� �*��~!������4>μ�Tӑ��(k��d�9���v���ڸ��1��X���'��m���[�!��Fd�
�˶����ìNǀqs°{Q�Ip:�T�J�����Qn�%Rj�w�f�)��3�R+���(pOR�����B<U�9a����q��O�u.8[��o�G�է��>�W ��syس���T���Is��I�	� Yj�%�cE��Ϲ�QȫDb����∌,ZN�5� �.���,�{��wM�C��~�q��n�ne�@F�)8�fL�ju(��ŴG0�>�&�?-�g[��Ģ��,0f�����DL��hR���03 *_k"���_쓯�X"k���S�H���Ĳ馋S�i�C�
n3@y��ǚi������4bDz�#��6(��}-ܗDH�9}���C�($�(F*0�^��}�]���u��i<M���IY&�Mtǹ�Ѱ1��j��vKs8K�±Z�� 	*�$^!3�Xh��HXr�O�(	�Ɓ�5�d��9s���"��T��Ƚ=5 ���rB%��ԗ�'gN�`U�B�-t$b��q��~k�'� ��/�";���E�~�\�/j� _��{�	O��(���s[�;C�2�Qwʂ�$5�	v�W�˔������W!)JB�}�Qưzv�ӿC[-�J@�Χ�Ƀ��m���n����dS�ݵ��)Y�M/�[��7���~4�N��Z��%c��&���z���te�o�#�
���	rW�2��ۈƸ̜&脜!�S���4W��f�g}�x�ϒq@����"�E<��W2Բr\8���� �,|j/'ị �Zdm�n�x3���MNf�a/N�0�)D�8j�v}^�k�'zq� �_�3{�-?L)n�_Ď�+�s����8�[�?_�p?m��Cڠ��Pn�m��ca�3�J9������i�1h�ʨ�5��'����+�����O!�Q���Q���Xː8˹;�B���y�0_��/�}D��,���m���m���GN�ֶ ��`˔�����9�����hH)=|�B��ѽ���kJ1���e5�`����|�m�&~�Ʋ��^� ?}i;Q��[>��9�����"G���_��F51��fF����w3���C�&�T�$듧�7��
�zɈ=���ֹ�w�Sr���3V���<h��g%'8�'�i,# ��k�;�v#R�q	DOn0�G�%?B��1�e.ȕ��o~~F��?1��f�ۑ���x����������<ív�}"�H;KX�SC�1�����:sw����=��E���O�H�r�(7��!�9�sE��1�C�y��H�O���q����`�a0�A��8����1�6 	5 ��}�J8�%r��2��K��7�bGG4����<(���P��^�']��7�sj�vF[���4�.𘟿6���e����'?OLX��%dm�_��"U�JR"THؖ�$�"��7��3�Ԟ��қ�8�x��A�t�;G�Vl�m���=F��tE:�|�HH.+��آ-�����q@䠺<�6��s�D�Enј�-���z��G_m���r��M���c[L?B������3&.r��P���?g�/Z"f/T�qp������N(pg��.Rm�O��8����T�:�J�#z���IlI�ml�b4s2.j_�ˌ_Q��}�B��j$PU0�o��E ��vr}�.z�>�6aҨA������Rq�W�(�*�%{|{�؟���9�w#g�q�gI����
�~ �b�D���TA��E!䕞���C��:�v���j� O�x��o���!��O��Q�`0��n ޵N!�b(3��hǪ�_n�Z�g�~��%RU�'�j�o��̉�d�:�^{S���z�s|1���+��z� �>����>y~wp����.Yz�	iE�������6$��d�	�%[lt���� W-��opr<��5��5��S��n&55ڥo�e+|��u�/,K��LV��<s�����!�GAulu���B���
�hp���.{�_�d_�=5(0SeB���g����B�A�"m�-M���t�ޖvK�IlX �
Q��t.1[��5���	�]��f���%�1��	�~���5��(|�j59�=_:(4(�0kx�1We0w����.�e����z&zc���E�z���p�>)� ��<M���y���M����#�ui1 ���u�辍���PS��W� ����X�h��eޯ�Rw8<��j�u�w-Z*�m:������T�.`��j_���씊�W����e�l��}-��nt�!?��1����{j;�+˱���yBF�U�3Z���mo�CG0�;��e��YT��6`�`���)8�κ�S��֍�>j^V=q���P�޷A�ߩ��ND?Ձ-.�`d"^aTW��8Ծ3D
�,�tzQ�[�m=�����I���+�2GHR�ߧ�T�Kp����4ӳ�r9��x�|.��缥� d�3�R�$�ɦ
��B	��o��/���"D�U#U�������҅fe�'�f�P��l1�� I��������Ƙ�}9�<=������̘�CJ�I�ܶ�-�'*g�	7Z�W�KƄ��^�����jd��*px�Qz�bR3QCAP��ߎᾹI|rX�/\�B�E&	�.�vC�u1aB�{Oy�_?]d�׽0K�䲆	kL��w}����g�+����5"��85�H�Ʒ�ȳ4p��x��0�n�<ݾ�ݍ�2$ a�>�ۨXS�|��nߤz@b�m5�8$��i��3NpU�[�总Ƈ��1~��OG�.�����,2�cs��Y��b|��mpq�G.�e����/٪^���iyK��Ĕ�������i6�k�qa%|̡Rʦ���ͷ�f>Oq�y
w��_�%?'�c���ݚ#���]���k��ȾO�*Q����E�XP��ajΩf59���w���yF��*��v)�G�t������h��u²>u�:�.�G�;Q,X�����m��1U��JO}��Q���掸�v��Q�R�Z+�H*����W�g]W=��,q��*��z�?dh��Pc�
���^쎴��������~ʏ-~՚ ��a����=���, 2�ܰ��԰W�z��d�נ�+���W����U��,�TA}]/@���(H(' $U�E8��<�Y��dEo��S���M3
,��i�(:�1^ꔞ�4��u�4�*Y�٥��D9v��{��0���Xn�^_l��e)�3P��
L�8~�~_�'� ��Q���S˽8q5���hſń�lG����8�A8Q�{CpH}��\����_ω�x����Y�EDf�d,����R���^��wwX	T�����X���/M��^\�,,��,��"�e�U%^�E�,;6�E4jC=�,d$2�I�8�,���4���n b�׏�!o���;Ʃ#|��W��%cg(�ڿ��x�r�Nz��:���#EfV�y�v*�+~���ߠ6
�e��.F]�6�)���\J�R��G����rJ�; ���8��h�z�Ž�:G�Gٍ�,B����R��nT/�m%(p���n�˺�c���E�d�a�D������� X�j���_JB`��5��[����i����t^��Op��gp�{���w��=�\dOJ�A��޿Ѝ˘���,Fx�p�P1#�Z=z���/�����l!��+�~bO ���u m�$@�`�-jm���u���ꋥ�ᢏ3���L�9A��yŕ�;�˒��`���x��\��Wr�<���1���ɇ$ �A�f�zć|�9�J��
,Z+O=K%7��C��Mp�m��fB��E�M�÷<�}cOȉ^���ţ0��w*�Q\�P�y��.�h+e�gP�I��wb��w?F��T@b#!��$0��W4EP��R�����������cc˩���;�)��3�聻��h��&�!}p�8t����dP]�sb��B��B�d)u.�M��Wt_��f�F��[
����k�s;cUXL������S���뎞��0��+jS	r��!gz���P�k'̶4ޓ4�	�=��(����'���U �&�O�Æ�J���[��/^!ƙ��.���C��~��%V�i~@߆#��Xg�5��� ʌ�����M�.] :a��1�S���β�K?gO��_J�&i�p-;��5���s.}�o���� ��#(JV³�ͯE�dߜ�Q�ՃAI<������Rnq&_Վ�믕`�ht¢� 3�MJ=��� �)���l8l�X(��5M;�sNpn���q3�gF���r�o�7�QȔ%q#�!�lʑ�����/�kU��'�m;(�.`]D����:�I˿͘����*��ߕk�`^���@�c�,I�V(j�j/�:/�*���'��yYYh���%�#��㦽����x�7rN��x�����Bo�����D�v�u����K���ťZ$&H����Б��d��œ�.Mmw���@|��=���i��H~��b,�1�83��śj<�x��=�̅��
�3l�z"����H��8�%'�����b�e�{��^�9㩀Zݶ*+�iA�����+}�ZU):S`a��I���L֌�þůc�KUx�O���K�A����I|���X'C�⃦����Q��ϛd��f����a�v��6�K�$�.Z/^C����<v�~MM�[!ݽN��Ϣ�So�|�,�(�'�Q1
͐���b�31�I�a��l��S���_g~Y��'��a[�	t`o�<��bi��#|��9�$q@���5�W���1�R3@�=v76�囌EA=i!!�X
�JE�T:���0��p�:xM��m���a4\���߽�l��M��l^.��� x���rxE �=4��58m�٤P��%�!���#���Ž�o���~�M�x�G�XN���gGܲ$��9]�x�&'܆��O���H+�g���7��L�_JaT���T�LyUi���Z�D�s���K��^Y���t1@Q��궙��ύtVjwG+���m�_�	k��])d�k���i>G���i9(@��!9��=&%�!���� �s�*�!��u�u43M�qBJ$�Ɖ�h�\b���l�Y���-���Ȏ�dq:��ɣ��Y�7�ý������P完���Y���8���&�@�5�%?��k����n�s��F@��T藃�לf:�"�>�<9@ E�0g����4-��˷��c��L\D�H~`�/+t�[�r/���,�/����[\��g�4���<v=����1!�chQ`S��Lz�
7`<��Z(�\�/F���"�$�$�X� G�B�#*��;��%���:a,�W��j�7Ц��K�ӬF��:�&!���ަA�����H_��ܘ-�Hp�?f ������k�V����xi8�d��g���#����t<�$z˺m�����������~ b��H�N�@Cfϻ����m16(cFA��p/r�vro�'����}���K -k$6����Y��4f�GƸ��)����k� ν��2�S� &R����r�];n����*țG��3�J�k4�o�0/�llR�@��M������@v�v���Rg9�)<e��K����\.B�J�eA�]	�Z}�A��|Լ�e�̈MI7�VFx��O$���H{�����m?��SDԐV\�c�(���#�y�
����z\ �?JN ��_1���a�h���UZl�-*�a�
�#��z���0���~h�F���j.B2�ȗM��`}al���q#����M�.н�:�"Ɏ�a"	��a��V]�+�C�3Z�E+|�=�.�C=QN�~"ٺ������[s����u�	P�-\Q�s���iE{y�m���h5�S���D��Z
b��H��>'+F�����R��J쫐�>־"K�8t�w{w-�0њ�O�z���>��̺S��
��j�0k;�\�y�!k�L���{�*`���Tr�p�!�J�v ;��	:�����5i�M�J\�˶�":
l��^X"�6^6,�O��z���x�M�;k-�%.�8�@�.�_rD����X"�?���e���ů���9z���z!(Jp^�gJOO��ۢ���>�E��l���@�r�bLKZn̪2h�]��[9�ҥ6a@N�Μ�RL��\�֥�HY�3��S�`܀���,%��5/��s�"���?��_ukS7{�uޖQ
�1��'��l�Au?�N�c���Xfb��^R���k9�{r�����P$�\��,��Ӏlj�<��s��ױ�rTƲj�b6�����f<������W���j6"h�Qn���^Ӕ,wQ|�l� f�x��EbD��Z��z؃���,t?�kX��q����������x͙�S��'�������F�M��6�)�~�@��.N4m��08�?�1��9u#}�a���")�(W�>"��
��s�5��6#���	7]Z�n1��g�oVHu�p
A�;]#�OJ��`�[G��w������!T���D��-e�l:��U��1�vE�|����I��p�u���]�m�����J�
�^ �H�Ԑ�J3`r����kOq�:J� 
:����e��J"=���|G�W}U������2�o��+����E�����9�j���<C�Ÿ۝�7c�Z6��U�y}��|�5����Rm��'�}�9�j�W�,DD�%_Ys��KQ�T�z��~����;�Hl��ch"ݚU��? ��}�"�����x�y.
�)hG�[� �ضy������B��H�u�OrP�g���^O���k�L�V9�v��K�؀G5B�ܹ3��%M�nUU��I3�S��5¤�j'wɬJ�O	|��>���}3�M/4_�%��Z�t�g.��y7J����*�@���_{��;��5�j�`�)�~lxhۜ��;WT-� j!�]�ó������&���nf ����F�{��||��#�wE�Ut�רΔ�D�9��X��"�:g<
.���`*�H��MuiE,��@�����ߥG��ոs��ٕ�A���&�4�z����� �e!*&~*���^J�&=a����3g����(�t��y�E+y
�^̩mS)��י�:$^�`uK��R�$Da�[���8{DO��&�Ҭ���ݢ�`�w��N���X��r{F�~Y�A]��ͬ��WB�Y��w��<]T��p�j-W��eH�e�ƨe�7����%
���l�m"� n-`<��>�:aa�/�����ʭ�Kt��S�f2�`j��݈���62�`+}�YңR�;�(��vSi�|7��J~^���d4]6�������^�9�@��$�}H�c�Q�M \��u�q���������H��;%`�T�MAr�{�6A���e���G4b���Gz~��.�tq�Ĥ䡊�C�ʾ1G�L�ϟ�&N�f7�xj�h�ϵz�����2�౻�_�	y�Q�HrY�� �#���u�T�K�\�c~=��o��n_����;k[7���(����;X]黑�Ƥ:����ƈ���gےx`��c���f���8.�*�3*�����2���E�'K�H
tC���8M\@b�
�c|� ��{��d���	n�8`��	j����,�����'���1�X���k0�f��_��R�d��U`�z�;�;�Б�Z|>N��������ū��L̇����.��^n�8b�(]�0����O��=)��zPv�}���(���� L��M_�C��+�^9L���M�bgUk�}���3�:?��7b��7�b;`B���{�)B�i%��G�@�QN�#���
e��ߡ�r�(1�2523�na�N�O�@�^Ҍ̸̔&�_��{�A�RQ]g���,����1����;e!�S���?���5�y'i#NH���Ȗ�oX�;j�y�j `���q+�c0��8��T+�T�3��F�
��w��<�Qi�?�q$M(fAٳ�[��_U�]�Q�����!𝗲���m+���"�}��*V�[�n��fXfL<
%�L��F�c��#���B��=�^w�4����B�Lw�Ɨ�t��C�g
���a�Iq8u��w7�l߯���wv�H��+\�z!f^�"��˒$2ՋeKr|���c5b�����(��uv��b���.bL�IsZg͘��|^9
���z�<Ӑ1�>�Q��PJ�42'"���:�O�����S�WC�^�-�X~�:R3,�^��f\��ON2%��1I4Ĥ�5��@�7��m��V�@
H�i�W?U��xu}��S����qoa>�����$748S�ի{����z�1�s�����g�cզ��s@
����ȿ���m�c&� N)��}+p��0��UFĀ6�*Wo����+���, �{g|�2qSp]�6���������Nj���z�w7j�|���>��Q �kE��7�[�<L~��|4��i�){E'
�ҥ��:{y��2O���<,"*h'*���G�h�1вT�D+/^��J9�C���UlW8D�Pq�P_b���$�Ox5��7Wm��$Q�LZq�~A�{OgHU,���4*]���I�c� N��4��.8!���YpVE9���I.Û��lM��4P�[@�T�q���MQ�ˣ�rb(O*��cOØ#]�I�gi�8l�����j�����-"�ӍBB��6Fd?�z��8���	SQ���s�,��;�9x3?�p��c		:E�}�2�1K���~ѥ����i㡻��ޢi�WjS�נ��)���>$%�KL�);���?�e�K�7+�=���t��$����	X�ӿ��~��l���r;QNu8�5����ev Kŭ.*!�8k�J32;Kh:T�7�%Vܑ� e���f'N���7��� ��l1��A4>Qػ�_�d�u�!�Q��Q�&W���#�����m��0�/S"��k,�����4�CSJ�O	5�x������d6i�� c��4�4��K�3J=���4��\���ؽ5�Af9&d��Ż���"+����J���?�8��K�6���h37�T;���P1W ���]��L��j�u�6�<�Ls����=�eN`TN�4��C?� F�m,��Т� G:���eV8���^�e�Eqqe��B^׈�!4a,�Leۊ�P1�=�����%2������%G͖'�f��������`Ϭ��a=�o�-y�b ��� ��[GF�^�8%��M�&@�\`��\#�|� ����]i)�NI3�v2J΋�A�:��ILu�1�K��B h���>�"4u}@Se�m�I��[4���8�3������bZ,�L>mL�ll�@�K�8�~V�0�G��k��*��j��ř2b<��ś`�X)G��Aյ�c��l��X��&�(�u> �Ne�q�������1�*�l �̯�6.�~�ݣ��5t�E{7��%��"�|�57QE���3��?[T����Ҳ���Sh�w�["��z1z�C�-]ޗ��Xl�LoKF蟛B�0�����L��K�)�<����80ٽ��p�^98��R�R;4������Z��͓�f����2#�s�����^&mV��	����.�1OY=v�>�څ��Y��^F8"��o[�<���4�B�[�ƚ��<v
=J��7�,����T�.�]Y'fSu���� l�>t�V�A����������4$��� ?�p�Ҩ�.��!	�ڊ�=�e���%.��]�����+|����~���SU��)C�?�3�d�/?�Ą��j���O��Ie�ɱ�b�S3C�y�uwo'�\7�xCOGI�����ѧ.���V�\�^
#A	��I�5�f�XF31�#�Ǝ�%P��mh�3l��R�`�����b��ta�6��.�-���I��zVPɋ��#;{��k!)1��m�ھ# �����,Ĉ0��p3k)��=��L3!Nv�1r5)�x���ww�����gA�ZKE�u��O!�GQ��^vMd�dYN���W-�ٮ�I�;y��+Gz2��Z�?���M@�>U���x��GGAq���A�t�A�a%N�����9w*UP�x�cQ)7��2.�S}UA}t������EK�C��v�z�@=�C�I��o���{����p�J�v�q�w�����&=��\�]�-�����m�}goy�%Q�Wlj�����m\b)��|�X���&�I`��2�dJ}�D�̖�L�4�-�_f@��F��fj<��Wi;�l�>����fP��%����ܽw�5�F��)l�I�Y�0�j�#w�$�W����[��a����V�n���X���8^p�-��^�>�T��N�?)�=o��RWC� �Z�f�_�$$?L��@X�.p$�a���� ܛ�0̮�:�/��q
c�u��3��}b�j(9JL2�S��[�R��͖����Ba��?7ߔ�����E�2��3nM��=�ϸ��!6��<ܢ(�i �O��9�)��
�+��x����h�Nѐ�α��#xJwoÃ�U�K ��m��k3Ǟ�4�Z���,B�Al�B<Z�'��6 �p�+~
C�I79����b�=k��k���/��H�@�d�����:�8&�n֢��s��Udm�7��N�t{���0F��;�#�ӌ�Ǿ�sG��z!N>i\���c���)6$$%;;/.���/{�渇�M��w�2�_@���ښ[�7�N�sU���P�dl����"����ܱ��c�A ę��3Bˤ�|�HH�w_�d˴�K�շ��zK�0 seoJ��u�dhB�UT��I�: E�lYe#�S(����V��8|6P�����s�^F�E$�3�,�"��_e�;ٚ�h��2N4�Tx�w<i�����4nR���p5�I����"ki-hzî��L\R8~Xp�<���0�ƚ8pBƎ���;��}UZxU���O��ݢ�x��Nf#"2=#�/qGLiZ�~ �T��p�<���-V2�Ӧj�h��a6ر���d���Ȋ<u󢓉Fi���rо	�I��UB<+⁏�����ĩ����2C�D#zCZ��S�x��sȕ��u]��D~���k�f��rJ��$|�h�y�Lyü{b6�g��e3�5-|�֭�Q���j$g���;��,	w��Mjd�M'���|6X��s
>F�8˗�K�ڰD^Q��
�CXV��m�m��߻G��&�m���z�h1>��� ������{����1Y���-��^��{(�p�K�����ƣ���ʘ!��,>P�Vh��*���Sǲwn�>7����7y�p(9*v���q�z�A>����ge�U��+f�K�m�A�l�LX��Y�3���H&Xl�����x��q>C�Nu�e'�����F�[�e5�y(tl�� I��4�o�s�L��v���	ɻR��\DꟉn��.�Ce��{m�+=��B5��=��V����|يwV}�e��A�1x�*X�?�� �2�'���/VO��5�� ��^h=&"�|��	�/v�h���0a ����*����Z�m�ޒL�N��U��� F����m%���>d�Ɖ�)�e恵�2�%��}��/�%+\���ʮ(k[W��C]xQU�8�^�3ʬ,��؝��$���n�
.��o�RIhI�}���<��ݑ�5�d��)9Z1��G�(#�55�&���ޯ�,��4��O���_d����k^�]����'�0�6�{7�|i	2M�/ʽ���0/zg�QL��m�q�"a�]p���$I�Βu����<�kO��6��⺳�Mouf�{�Ԝu��V�� ��*l��f��\Y��x�_���U4��E��X4��еpH��2Ӯ��D+�3n��&,&沂!��B��;om�_�VpuW\�_t)J�W�U4�l� �ĪY�:yB8;!sD��zp����A��?����e�� �X6{�'X���I��J���������ybS6��G�~@�ğH���@��iSf���Kt��o�&V0�>���_P
M�0\9���5���.a �Z��?��yN�}վ�&��}��K+ҜT�;2_�߫��vB�S�;!K������1XnV F��T��[�4[R�� OV^�9���7�r)̳l�m;���<�g�� �&���N�$}F��V���Қ�>w���EN՜]����0zuX'M���[�*��fG���=2
ٝT5$�MT:E.EwV��G�n��uM�8��k[�6%���|p
ś�6Æ�28�ʽ��f=Qd���p�"��m���Ԯ�!\lpaZqE ��'eq��fT[ ����#�*\R"a��?V�����2��6w3�īg������Y~PP���X6�c[O뼨�;�����"bI}��ܹFH�-�5^;�Ά�84�q��,윾��٢탂Xd�tL~��+�2��(4(A��B0ʨ���L����G�]�Ϛ�F�w���������
�3*y��F�Դ��i��u�L�A]&J��"�L&Џ<u���	: I��Fy�b,����s���l�5��C]��źk�IU��S��ҼTϝӝ��V�.�L��N4���sЍ�g���}���Ypsd������Ӽ��
���"ST���$3k�}Cn��l�:��6�F '�K(��`^_
�q�.,Yx��6AM����w'z�qpw��@�v�ѹ��I��*�7�	恁�:uVҏq.�"���\c%0��hL:L�"���[�V�q#r��J5��.�np��9P^�$��/w�.�75��uM$b�o��)AL}�e���:��@q������Jr�>�w���8.�nt�4��/8%qV�Y�^[��3ج��0��,2��!F�^�$�MX�p�:�DM�8}>��Gb��-v�T�j��N�ַC��CР ��bA��6I�g�C ����M�1zH��f�c���9���D7�$��a{Eʙ����I�Fն�d�ڽ�c3�@0H��0R��}<��܂	m�l	��Y�юHʶ�$��?�<���N�LfNñ��5�t����'N��#�@��%�ƱD���4����`��k�*�� �Ά��R�ːl�Έ=��y
!M�R�_�F�m�4���zz��eI)9u�Q�&�Tz�L�������/m�Ro��?����,M�S	�GY6���i�S�1&�,H{���i	Ē�����L��iQ�K[)��7[n�Y�`4���W� Q��eԡs�M�2zǜ�fs�[ނ89�s���
5��m�D�%V��.7��G��@��ZzqeV��'�!��}˰�L�H�ɤ�4��x���t)J[*Rp��u��4OY��Hϭ�~.�Lb���=�l�_�L����/������D��6,�#*,K�!��v���pO�Ȳ�+C�� �f��h���6�%�?=uH	���b�Б��G����z�ђ��	�6��Eη/���s����s��K�CuoEc�F���袐*�HQ0��r����4�'~e� H�`n&5�T��nz+*�2�A���5<ȴ)��w�/�J�>�A0��D3�{�CU��J,�p����#
�s�6���M�6@h�u�(���;{Fi�����t�Z;��T+:ۅd���o�	�N� �*5��a"�~[��m8<���4�A��z��9I-ƪn �S��V;!�!��t�ә��>����9Yt��~�Fv�K�j����=�cݧ���X��F:Z'0�_�������m�s�e�a��Y��b���k��gݖF�z�bD�;h����	�g�r�aIz&y��C�o��qD�6��2%GN96o��D9]��,{#�d�^F�^�7�G��3����N�	4^�}�D�: =�f��1{�kUU��I���|���[�W<ѵ4�O�"7�2(�� �ZY����t�:DV�cn���)�G�D"[@��Z��䞽m`+l]M	F���v��1XЦÿ�,�k�}��A�,=S���m8Ϧ��'�=3��zJ+�C����,�	���8�OV��ٺ�jh����)>�+��p��!��x������}��.oW]�_S�&�AwC���$n�Q����t$�y �Gmz�7A��6�aH2�&��%��0��m(ϋ��2eϗ�'v�e��p�MQ�����支���1�y������iL4�RG��-	��$m*����)�f����\��3����i�B��m
w� �1�?O��QZ�:�'̫~��):���ǡt�~m�"=��X�/=�pm/�:�M������ii����\���"����/�ژj�zOg8���4h����̕��?��� (dˍ�DF�h�