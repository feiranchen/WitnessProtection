��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX������`�k(f�MT����|����E�do���j�i_G�G;E7|`�3D����"A� F��=�z/� ���o��	�
*��	~�1�=��F �:.`��q�2^���X��,a�2*M�	U9%2a?��Q���|6f�]m�},̚��Ȇ�,~%9��ꄼ�S�:x�=��>�Vʂ��BtS��w��q�J�M�7�JW�i��\�y7�m�NM1;"�U��HKll�b%� �p!��G�)9���R�,)bR�Y�d�C�!�(&�2���fH�3�Q)I}�4f���M�ԋ�"���]��2@ŭ8 ��CH�ќ��� ����}����Ҍ
{�
}r�r8$P?�W����K-Q> !�| ���J��~��:]Aβ����� ��K�� �[�[' _j&8<������g)% �s����O���vݲ�����>x�74=���`�����b�s�<[!�]�������;h��le0-l��	)۲��-����ߛ!0`P��O)|ތBR�Άs+�_
fB�6GTm劾��1F�ݝ)��+��Z�w�v��� t=��aFv��-׋aƼ�s��\Q;����T��{~��wEc��>$�j4�s,
�W�\E�p�OX
���_��K!^sx���cK��xb�Fx7^u֝�E@ ֳM�\@�GA�$z��y=��@ٔ\�)���\��9=�4T��@�N�C� �p�9�eRZL�ڍ��a,Jb�_���\4���\�{{��(ldp**�`'�[�
2?R=�-g\;��^��*/ ���Y��ށ��>�?I����|a`�N���vS��;�|͟O+��#�W��46R���h�{�;�B���,��u��iKд�>�6�<�g5}7M{�����-���'�S����9X=Ȣ��(�mp�X`x�7��-S<Hr��m��s�"P�6�����׃���_*�#;n����T����1 p�y[���yB����䛆ܜ��N{���y�>�sA����̙�r�оy����\���gnd�~��S���_���ű��Er������X�8	��,����Ki��A�[M%u��AN�霥L�5�e��?�"AN��5Q�Q�\�PD<c1���Z1��3u�rR'7��24�!T(���Yi�z��.XR��1�A$��!庥���/(L�X-Ք�����8�k����*K����U �,8����U׿��+�@�� o&�̍��^;aW�I�c@�w��V��&WgJ�E󁼨�K�W%�*�"]FH�*��~���+�[�y̨�0S?�9,7E~���_�\q��� 3Ӿ.\P��<e�dՉ��*h:&�O�W턢{�[�Ȩ��2�
Q��:&Xſ|�o��&nɢ���%���/S&d�DI4��rE����!J;rd����=��ٕ�{Z�����! ��Ân��l���|���	�޵�����7��B
����Pq;��U�籟w22ywp�o�D㸺�s՞"�\�����?��[k����,�?����f�[ݮu^S��+QI���1�A���1�3��Pv��'��ѹh�PP�*����'�<�	�|���BA��6���L<s��"�3��g�ɦEe�s�>,d�q�=-�����˲��-�,����2jA�M!��0�m��ҡ��8rqi6�L;��H(�6 F�i�{�d������ �E�b��\����ǒ�;����d��T��s�45b���G<D=u�w\Qg��svgz	��3N7�n�k����nA�����Hd7�pdƅ��	���D��)1�+"���J�(���W�d�tצ��$#4]%(��������%#_�_�0�Q{�-�֟}��_�����	xҞ8ӆW=i����𵤿������/M�|�7/�z�t�c������\��Zwz���ʧ����+Oµ�a#��A��42��R�~#�?���:&X��N�Bm�+8��"Tf���3cCo�p��n[W��2���w�TuE`�#Jk�	�"���u_�r?)�:n�ǩ��yC���c��|4�	{�'`�?��GQ}�2�u��$���x��3)^�=��B���0~m�l���]��	�rz�g�� ����<ƕ��-R����Wc�u|l�*˭���m���ؑW)`d��Yi��r�2�J����k�{sA��_��K�8��n"�<'�#�?[%4H>#H]~mP�ۛAN� ��H1w�m��)�%9?��֤����7^�;��U{�l���K?�2Z���#�F�����C�S.��N���P�nlU��޹J>�ok
��qL�)��I4U|�m������8���G�K��Ø�����R�H���X�Ƴu��\^Hlqʁ*T �jV�J�"'acN�W%!#���%��PT�U5�L.���!��_I���v?XnH���p�B}��N�[n�Ko�lL�4�cͣ��r2m�P�*��<#�@�
+b*�M�CTZFOD����C�Ԗ�V�{X��v�2�-�HE-��Q`�-m	P5����#4�x����)�0H�Uly��7G�G�5�|��L�T��k���p�she�P��%�|�~����-O0�������+xX��q�0�J�����ظP#&&��Ԏ"u�ν��KL����f=�z����p��;��۬A
l8�co�98�;~q�Н�_DA�WƯs��f
�}�,{��H�];�M`�J~��vj��6�ծ���6M8���fb�p�<p$��S���m���,9�~!j6�{,*�i�L���T( ��z��D	��� t�b*�Ըo,��P�)��qw|`���r��V�l�%,I�݅��)�XA�?�[����eX�M�E|A]K}2���vsZ}j�_�����#�DW��"��+���< f
xX���?}���h�8Ҏ��;39s��f�1ʟ�6��A;��7״/����M<4���R���Sꡍ$��k%�}[k�9�����!`4x�6���fiW�^g����x�����!?q�*�S��hq���*���\}ѷhm~gOYP�iq����n�z��L�`���fZ��M��?EΕG����/�~��Y牯�(�FL�	=	3�u@�[|;]㋳(s���
v
��W�x#�c����n�_:n�6�(�b�H���I�(r�ˊ}b�����s��oB�6���k������9j �r�s7�iC�
��\AXT,�iCF�ߓ	��� �5��_�<z�(L��AreVbͽY��?Qeq��=M1�'mכ�F����s�D�d�t�*!\[�D�	,)*&8����̈;j�rN�e��S㐾P�~ĺa�[�)��=��vzA�!�6����*ݰ@.uϛˡ9(�u�M2���^u��zJW��cX�!ݪ��Wĳ]E�h�^����� �!��K��������N��9��9��n�ػ�u�	��	񼁥���.§^�G�l0�";n�'ţ#s����+��]�e�h��I �Ǫ��6�<Y����,U�eB�)�!?�n�uT#����'��-̾�bԠz��j7	d��v8���Fcݮ�B�x���!d��In��6����V�j��_�ZZ��GBbS�N�o3	0.�DX�LF bg�w���t\֏E�l�aQ�1b�y��W?T�� �Ć��_���8�eM�}�P��^Eߕ+����x|;�@��)�&D��W��
�j!ZX�f���0���%iç(Ċ��"��+I��־�+�]���}\ݥ�I�Y��E�s.c�O�`�(�2�a�Uqֽ8.��04��o�]`(P-�(3;��S]�'k+Ե���|��s��f�I�1{w�5�ӆO� �6�k�����/��KF,�mל����%'X�4v*�k�w�X~�N% �\u�m<�׽M?_]#2�;=��-��o>�q;9V�-�d3�>7_e�0��۳l�~��w��y��t�@?f4�u)��=�I#��cީ�7��e�:���kCng[��n*6�&��(�,1\�]8Ô�A���o�d�tT8�D{�[�k�א��j[��5��Ҕ�ì<��Hi �Ŵ����^"C5���$w�O>$�u]\���5y����.�3�
�T1��
��'3�����Vn}=o�y�_�8
����n�u��`Q1:i��y9�fuA%7]��ҫ��	&N��lB�;���M8�0���~��=H]Z����S��h�gRR�b�(a3n�BC�<V�I��6� k@�}�yV���	�-�%�G� ���D�s-~��o2#!<���ǤqD�ӵ���"�����VКE�:�a!��L˝e���E��ҐdY/T���쌌5�RN�n�FV�>:=:�]mE��^ t�2(����BX��>�?|�~��ܳ�r�x�&�< �����ֱJ��=�I߈e��q���=#�Z���q�O��p�*w�,���i��Կ֞����+�.�Z��=W��j��2o.�m�o�����I��N����g��5U����ܗ$N��Oa:q���_ά��MV�>��ͮW�QA:�{�uV�2M��  ?Z��N�T8Y�P#�����?�[��I��͘f��'��(�G�����M��B��!�����'��le5N��-�ղDP쁲�iB}o�5ͯo�1��p��w 6��;G�GF����˱�'��}Â�?��k��e ��A�m�D��sZ�&�>�l�9��+!IЙ�+���������Y8Ӟg2�5ز����7��n���O�	��&m ���� �Z17���[@Ā�W������Ƭ!��/���}uY��s��_��#A�Sᩂ`H���~��\��L=6�]k���w�]$^��ԕ�u�x66����jq��`#�ߠ��K�b��Rh�N��2eX �0�M��@ p!B�.��whE���>	���:<�x�������0߼��e|�����1��NHr�?��~E�r��˫G�_�T0���7ɲ����ґ���K�Q��\W)�q/�=��
��@�g��<�h?������{��l��-b��1܌58Y�365*yy�%-$�o2����;���T�H��L�_�ɰh������N�믥�X3I���t��Bw������|3�l �X���]�AMh�ٔdf��"GɱZ�iцڸ�_�}c�����(�@��C]�JFᵝҊ2�$���f#)�yw� 6�ļ���I�x�%�oD��u˰|���pn�"�G�W�L7�e��i��X�������Sy�h͘�1����W��m,:d��ufg��A��0
T��hKu޺�;�P�����q�hΈ~4� ���QI�P��s!_��Up�j&�a�T|���#=�="���Q��C:dLBba���.�z��w!�!��F����v��ԫ��M�v~���Nֺ{�7�����R�<�G��3Է��i9�e{:�,�%ei�.�Y�&���_#BۤJ^E�G��h;N^�P�^3�Z#�L'�x�AG1��Y�4F��}��Q;�X�'�-qG�'(��j(�&�3)����U������U�����5sKò�S�<C�CD�s���M$ �����Y+{t�r~tv	d ���#?]p�2���ڎBXx1����[��L͓�Dh�I��Զ���$R1V�t%X��'�J����,k���}��j��޲zJ�`�u·�ۻ�aFC=݄0�����x���1�uh�F���V�q�}2�{���1�� JC˜�$<k���,����9�5�(tNSJ�M_��>)�b�ox��I2I����)�[)������]騻���'=ˋ��f%߁�����}��Zq�8��Lyb�Mn���14"9����V���H��D���l��>v�؁�f4sRk�?5a�����:�s�"$|#�U�L�Y��z
��8�I��4W���O�d�lР��:^��#�q��[�I-&S����tr���l�{�P��n{�5�B�y#k�ʳn�RO+��a���|.�>"�KVD[]���At�rW�.l��M��"E4�o+�_W��L�_��s㊔�Q�(���-6��)����L;�ߧH�yXK!%�W�i9H�<�tCc�\�=��� �	��yE���~�Ǚ��d0���lW�
���YTD&�0r�b�%�@&�%�����Zh�눺�B�A�e�?�/|*b��Ag� Y<G�k?��dX�0&��l���*��]_��L�	�ֈ�D!�����7	G�^���(��l���ty�A�O��-����A�=;�7)*/���ex�ϭ� �;;�Xz�OFB��lw��KY�>EjgH�ojN�x��T�R<3p�o�/��|uÁ�24���/=�!�]��X�vLg+pb4" yO��6������e����������O@���3�ޡ�5)��=|Mzl������)��xߖ	z(�d�a��YEHa+�m�d"/[�S�;Z0���PZ!Q�T+ֵdJ�X�N�;Qsk�맡,==s�����t�	ԃ.;�´a��?Ҩ9j�ö�D�*3C�w����U1�=]��?�==J0��:qzر��øO�yvA���N�������+�q)�Sz%�ͻ(g�R�v��~2,��,��i�M�j�O��%�r��CT�֙Ϯ���Kv����o���@���hY%���m/�[�|�K��	 ��{�T`ϫ�̀�����#�M��0Q{n⁄�d���it���U��6 ����@�qWNɾ��uX�_� ���4{�͎�Q8�i��xMl2��a=�	�%28*�6�'5Nhd�{9�vjڧ�����q��d$�����xe
E�+���yw�(���a�]>���Y�M*��ֻK�&bL1��\�<(����l���9%r����AELC����T��3QRuX�������(��P���������i����d����Ѻ�!�(ښW�gǸ��D ���}�V�y1c��u�K���S6�-�$=���±S	�6{g��Ru)djy�A��z��ޮ��%G�煗j����D�i�Jz��z��ĩ�:���{��Bxqg���M�}v����{7O�,�I�c��_ո���{g�n9T����-	�$+��q�np(�1,��7�r��[�d������XS���ox�N��K�8�����^)�$ ��tu������\��MS�38�1<!G��x"��E��	����i7h�Z��.�euJ�=)#:�]K��Ǧ��1*p|)�D�u5��Xjλ+4�zq�)|�����lM<7���������3߫b��+�����1Y=�^Hb�C� T�5;
�W'��䮌 ��i�ϟv�f��mr�܏n�h�Ҟ�f����������Ϊ	���Bw�k�fU�T6(���;�0�����L���z�����
rheDp��{𐻮�$�1εP<�>uòx�$��q��P�k����,���U=�@u��5����؀�5�K-s�G3����d8R[�PRo9w a��+Q��$�4ݾ�E�ˀ��'j�~�N�^'��Xς��=b����m���ή��"-d@�!�m��z??�s$��a����.�`׺�}���P� J�g�ya@�-�$y�qg+�N~J�f�@B�Ԍ�S�k7�uǄ@Nu1DqX۾j��`�SiZ�ş�Q:��İ�+�qRi^+��X��ysX��@��1I���g����rt��$p[H�6�_�D��+w3u�i��!C݉%.�}��	�1�"����=�'�j���a�e�v����r{L������|����Eg�W�n�n�KՍk朲׈P��Gĉ!�1g�"�I��)�~}����ݧޫ���T��U�u����^*��������y�]�����Kފ�v�Zs�9u��Z;�!�%�X�^�A�(py��qέ=��"���Tx���9%�ǭ��~�R�[�v���i�c�J��%&�c���5�g�
@i��5.�;~[.��۳��~z#�6è���4�OdJ�l��3(Vsd�K{��˥��Ą�{�;�~,g��W~���gvԑ�O+;т��AR�E.�E���x�Ρ����qk���e�����y7z>��7���o���K��Q�hx�R�Z����w���%;��5�/"uZ�K׮�e<!ʄ�`г�9wi*C7�b���
ϛ���pQ���D�>�����Z���cR�ۜ�ƈFdg����pc����&�⦜�������[O&r^�T/	A<�L�;�<{tz�l�Qоy�W����Ԯ�X�V��W�ͨ��Ŗ��/�b�w&��ِh�$g$C�ױ�m�U��rk*f�C̀Tۦ�%&���0 ͍�bڄ	%.��S2�@�Kp��H���!�[�DiYf�b�<�jqcD4���#RE�G�Y���3Ցy��\���i@����)���a㷤Ԅ�(�mm��Aj\��Pr���,y��)PM/���.ϼv]q͇�TQbQt�9������Ή���r%�F�B�JW�x'�����@���pC膔��������]y()fM��_g��F1FYf�Z��1��ݝ!��xۈ����
d�Z�9����,MQ���^$'}%~-��H��1�j>���(*�ar�
rs,썼ܚ*�+��3�N��M��?�;x^�5N7m����O�_�	�8;7#I��}�Jw��o&�~�$�Vzgn�	Ө�O�R-Hu������d��5������i�m��{q�2�Q�>�6�
����J,��r�������EZ��Z-[�`:�}�쫵Y(�t�_�&��A�P���*�C�?b����ps�&BK�����}�g�}�+1��8�q � �u	�����eN�c�� ���!+������sᦖ�n��w�yM4
�E>+��� �C���=�j��Mj�ar�`��_,�9�wI��v�^ �;��(�I)�-��(���;=�9�a��I��Tp�����_�}���L�3�6�u����������p*����׋�?���c�h���I��d��A���2�2HG����L2"�����l�^�-�ޫ~�zd�E��y�r5d!v�3��v.Aw0F�n�\6*<t�!��/�M���F�%u6sc�	�nK����X�{���ޚ�ʿ٨K��G�U���P�v��c
n��G�j�gA�E��k���a����9"|ѮX��H$��7�������[������/F��*`���a߰ājJ��0hOLWQK��SwE0�V��ެ'��a��SI�O��輡�|�'p�'͐�]��TeῸ �~iZt����r瓠���{��JGV�D1Y~���� ���'�d��A��ԴE��s���眹��e�P\Q?;_�u6�p�:�_�?��t�)f��s�<�-J�Z	V�)�Hݻ`P2j��-�#>�N�e�$�.��W���jc��,�!NV��IEu[Zm�]���خ�$�+�̕��#bK<� N�z5yk�0y�ot�@Ӱ�2��V�<B�����l~v%��hW
��>�.LU�Y��J��ax�wj�;;�Č��L�T��0O�l�$��[���
�wHK� ���\%P�0s@o+�-�L}?Zk�;�O�M]7�'�9�e?[���QtXDQQ���f:�ڮ�+N9�=�����)��IG2#����{�+ƞ�U�'���A2l3�+�+7y�*2���<Q���^��	��%�ru�5P�M�x��N?�$���Oi�VS�ݼ�&��u��"�&�x�@c%Ǟ(�p>>Δ�sQ�p���	����;41��K�)e�������c��z\�i�T��($�<dr~G�?f��*��kJ-d�����8@�D�0+D�g3D��E)�/����j��rw�Ze:���3?o�k4�RfTT��c&����s�"���YJ�\�G����|�k8�+e�G�R���� Nn:�?�n+cosR	E��T|&�X�ኩ-GJ<����Q�сd���$����]����,���R���4{�珩����,��0�<�_��Z�0�x�X�]�ݪ-�T�>��O��(y��)ۦH�@<���rc�A�^�%��D��q�aZzi t��4Z�/B��|GY�+َ& >��IQ�� -=�p�.뵂̳�5�Dy��k���W��On�?��~`�bW��w9�O`Ѧ��bp8�+���]mP|x<=��8_0�I?�-lA�k��d	RX�%��xz�79)�G���ds�N�i�9�@��̇x�׮LD�a�ϥ�
|r�,?_/|
1*�T����^�w�?�������G�/\����z�(�V���c�|���>�_?�:-2�b� ���c�J���
��E�jIN}|�]�i�_�$�����bm��Q�(���Ʈ�C�գj_����X�縹�	_���8=(1ۿ�3D�a�R�1�d!�7Z�Zb����Q=���C�,���������UD�|��Xv+d�D�Tn��O��mf�o�i{]�Qt1��`����U�E��`�������>��?g��%(i�K�*�z��F��t�i�(�u�;ڈ%��G�{+�|��(���t7o�dI�*>���MĨ3p�?گ�-���9�
u�G�ƺ��נk��-o��+c�b���@$X{w?}���{�@w�*��ʔ��/�Q�U���b̻@v5�_��ɞ��@W����@L.c���J�K����Ւ�`��C���J=s	uu�����y����cu"V`{0ft�Ν�I�I#��U x�_�b����5��s��H�	�Z�D�`w����t��s�v�A���)-���>3]v���9�8���	-�b6��J��R�F|b�9J�w\�:�@��S�����y�X�8
Q#Z��2H7���ur��
�9}��uꎮ��|®����*��g$я�]t4�ӓZ�~o{�t�E�x�F0W!%�Gq���ѳ�|n��"B���NIm��0����{�D�svg�[�_���_�v(nSzV�įd�$H��?Ԗ�{�iq�]%���J���5�����T���N�Ó]���hZ�	|�4b���I���g#���M(=L6�N!��a��z�Wy�K��Mw�UU)�\*}f�n*��+�.Э�����D���17��F�.@Kѡ��ZɛJ�n�����YMض\�8
���?�
��!.�y�}?���ܻ��WԂ�m�/е�?g�O�"%8��)��f"2�y��y��ǈ�w��E-�5.�v��ץ �tH�XkV�����4M�O�f�}���7�&~�M1��@"����6�fb�D�<�#�
k �
h��(��$��22y�h�-CYdk,�u��Y}��4@�h�=��	�k��Ub����N0��br+Π��hF��jU�[Ē��������X¢s��s����	׸/������Y2K������6��h̾����"2HOC�SD_eD/z�&Ik��d{�o�K��R�"�U�,���n��tN &���R�T�?��U/�!��8c_�/����;�ܨ.��oy+���,�Dm�PO�ٓ�mZH�2f����RDޜ�⺢w���@���<&�lR:B��9�=3�=ʨ��锆�+�r�)���S��?"[�����6x�l6!��x%t�,+�0�5���� �.�5qnCiOE�)�	��m��>g u_��bU�J�Xr�	��\s��%Y�����^o,�r������l�G;uD���l%TAP�D`���)Cmc��߸b���79�f7�=�-��Y�S�oN�̝ؐX�;�GQ_]�,�(���m}р��:L�2��$� (�{�,女c�M�x��n�%��BT2��W)XU�Uw�j��~ J�k�`Ne�[1�� ��[TwM�*���r�L(���f�u�j�s�l�����8G<vt�o��1�!�[CK�ѕ����	�B=�8��b�o�����	���S�W��dٿy2���R7��D8�jwD�*)� K+�d�DX��gI�F�#T��֧��3�@W�D����fy7N4կ��0�ͣ9�\���0�����v"�9���]A�������	2�;��s�����7��jj-w��x��'�Ob�wA�~w�]�]_���&l[u��G�-,,aS%V��+2��_�@�o�H�ET��ն��B[m����[a5�b��Р�P��҇#��_�1�����JHhWT2�߲:�%�*���KY����dc��<�D�_��w%��1!y0�������C
ު�*��/�.G�h��@�Mhˋ�@�S+����c�ճ�x�����
e��ذ����g��"���V��V���0�gt0�?8 .t'�Ҭ�!���/EԳһ,ηNh�e˧�Rdl�w��>,8[�l��X�Us�Z�P�l�oK�^�C�U�C(�2��l2����iR���+���1u<l��SÏ�I{̭&��z߯y���6�j"���a}|���^����q���^^)F�~],\2I��*��~�^�)*�.�]���n]��a��-s�C�bjS�@�yb�k��^p��p�.�k�}��䖍o�)L Y��
�;T t΅M��>��fU[��2z߽�3$ h�T��3��.2�E����ɰ-�y�f��_ȫ��*�lT�s�wr���׎ )�5�u��h7��7��t��5�%R�T�D ��S�%��XX+p� ӹM'P����`�s��$�͡͝w��׭Z7�:)�#��R�|$��N�K���{*�=�{y*���7���'��S��oQ<���۸@�N���Y�ԧ�j���Tx����0Hn2O�԰�;_��x�S��
�E:n��^� f��!%-83�ت�Ƀ��~�4����.����r����;ӕ˅a^��h�h�����T ��K������ճ�Hl�
�nj u	��_�y��O�gI^�ձ������ke���|���ۈ��<��:2N$�{R���Aq�0��5.�[T�5FJ�؛Nu�9m���C&)�E�wPU����K�{d�Z2(ȏ��5}�DqF0"`˲OU�ҧҎI�eǰF俲_�Q��ꚧTAO��ZF��RTC02}��̲r�A�[�jn�HݱJtǩ3�6�4�;���\�5i��q�j���ا&5se<��DK��LRC�	a���e$Wy�$�t\?��bp�	ѷ��5 �e`ع�=Go��Ť=�#➬H�Y)JX
�y�����2��}���ԡn��uC��RŤK+��R��vr��G��?�H����=@ϟ���;�cJ�^յ�O*lۻ���wqfT���|��I��}x}fQ��q��������R��]�lJ��û��e|
���Fk:�S�;��]�`���ЖQ>ʫ���A�I�Ye[#�l�IuQc0KDi�\X��w8�A˽�@����_�r#�`r�L�J�0�z�Wʠ~/��~�ӿ��v·`y�<���mw���H����l��@�c�Q������3;��,��ƣ��H�����!�_�9����{~\��G��� *fZ��f�����>~|����u_k�(;�l����M\�č��PR>DZ���/����:7} p��γ�
2
��ȆBt����(�n����)�^��e���ts�6%)n)���ӝ�z��&`��xvr���f����m�ܮ�a��5>�î�~5K��h�T.��(�U��v�� w$��7ɺ㘟d�{��z��j���CE�R��PA��d&?��;�I%ި�qo�偐t��p��)dg!?Bu�j�SѤ���:��+�������>$%J�ea6�.}�ȋR��|�x�Z?h=��+v2w��'��l�N��<5�����Lu1(�nL?P��ϨU��tƭ%6����+�s���8�-�9��t(��%ߢ�J�#�)۽5�>(�Qɓ���ċy��4U 0rJ��Gb�\N��pÖ7��Fe���K�[�~�b�ީ҉����5s <;#2�Gkͷ�Ff���"��sj���6���ϻ�v�k�M˸*џA���T�H7�Wu��j^h;�����������J��'!�F
r�S� ��-_��Y,|2��$��gSl*�Gk��y�:��l����f��eۥ��Io�>^0�R@�����\�w|�c�_K��_�}<Z��Ո3��U���	��J}t�~܍�)/�+�O��~~�}�q���s�f4�V����n�r�Ϧ�s�,���_T ���}:-xa���z����q}��p������ƃ��Q�y.�7{�z��k�	��ND.j_�0��/U�'܋k���v�N��l�nW�(&V@S�h7��W}��R!��o��2@����je��S�H���͢��c1`���>���೑���H���=��P�L��W�g
���M��V�����+b���#�
���Mx����c�=��t�g{,7kap�4&i������>S�N�Y��8]P��H⻃l^�͖"�پ���y�0�!p��kVϊ�	��6�s�te��}B��:�Kڰ�tg���NU�,�K?��E``��㣬�r5޿�1A���k�y��h[��#�m�bjX��ܲf������7;x�7@(7��;�*!��F�x���f���h�c�l�����!k��uQE���5^���ey��t,��먬���҄�E��9z�~��U�ڛ��-)ꃾ$�T2ygrX�'S̑�&#߾ \��K{V�:��۶�j�tc���I���g�6�uj�c{R�~eN�6=^�:���a��$�*��q�i��S0l4:��S�Z��L���lƙ���ff�]����@<�����U$���O��#�x�(�rW+�0$*&�)�xf�^���]�ΰ|"t'��/�6b�fC�D��J���G����Zӂ�壛��M��V[fb��z����f86�ד��3�
�E���u�����hv�{��,B^�W��r�-`�m2�\P�]|�*�/��\�#��@�b(����=e岼֭C8'��~���%�����B�3ݪ�Fk�Ý�<�2��iz;r�YQ̀�g@�7>�Yߓ�����s�o���JP�O vc�5���Gv�q!�X���z �i��U������>nG����iVA��_� EfI
�w����J^��F�⍌�E�YXTX���jve�'���|8P��^rPW����y��������5?E���^������������Bd"�_�v�CYC�<k�"�l)�n�_i֭z�4��=+�0=�~?RM\�H��1
~��BӹM�F�*A�5�27����Y�9�I�_��'{���wv�q|���-:n���qS�ȼ5Q�k�+C]h~�E�d?j�kI��;��c?49�Oq���i9�%Ƭ��ĖI"�0�+�gÁw��G|�k~������7{�s+$��R��1U���Hb���=���LX�hrfZ��#`H��mjE^���p.b�[�q"T���4�u�d�j�S���U�Q�N��KQ1�D��Tt\Y���e��2�L�+��k�a8j^$�����;���L|$�8�r���}�|?+H�J�_		��g����'���:?�P:�`� �=�l���]a���,(�����1��B����Ѐ:Ȋ�PPm���s�[	O����dpf��N ؊��A��AP�dmgm�:������uV��7D��IQ]��8�3A<	�Hyת�(?���r�������U�6�.}�����Cnb�f��f��k�x�?�R���:
Px#�\/���Cyh�'ʮS)�<�\��F����2��I_��N,�s�ǣ �T�С�%�_��;L*N�Ҷoh�\vd�?qI'�,z�N�3*֞W`$�N/O�ݪ|��Қp��0��%�k�:�|1��MC��z���褬jp��>�O9���o�X/H �Yhu�\l &K|��働 3�^5Y(L��.񸣭�h}/���_��x�S+���[%n��#�z~��2��j��	�F$B�9������q?eǛ"���,����r�x|���H6�t�9#�FBkF��Z�X%��9�f=�~:��3;M/��c2�,*-p�jz/H}�gJ��*7�S~���^�F
��;�{9������3~%c��G�SX��c��{%N1A�-$�d�4��}#|�@�w�<%��0�mT�s|��ڍA!Y�!�|m~�a=�� Qy4����Rw���{�����c�/&6��m�2_뤬�9�q�a�:%8��T���1�轖���n���b8��x�����R��3�ɽ�&�Ӹ�ǩ���"a'(�����M�u]=�_)T*��qh結+�	}�Y<�I�K.k@����~uy҆��_i��n$m|�ak��W�Q:<_�z��V��WL�ސ�Xz"���V�E!�(�1 �I�~K6�����ϹG����M'��u�+׉��Vr���}k�
`�x�$@'�.f?C�O��������~�X��^Jn�&�uV�-b#�����K`�Fv�:_0���l�dc_����y�/�H)���^�k��T�g*����U�(ĝ���%E��Mo��m�Z56�vL��$��	����E$�����NƷ���Je�K�{=��-�9�rv�w̽+����x�tt��-��\:�
�nVGeV��T�nT̃���/�jI�+�9�y��������k�ɣ�������&�|�}��Ѕ��a6i��`Sn7hr�Z��ST��ʆi�느��R���6+�����(m�z[���{s�J6>����[B@�j��&?V�3v����km�)D@y�!�!,��<v�}V�;����8���`8������ ~�o�BF{B�#u ��ҍji�b.
���ϐ�e��~ՙ[����,O��:�'�)���b-�����r�e�*���?d*Ћ_�n���i�׍��o����,�}_���^��@��cfE� 7�}�6~岤���,;�2<���aG�o�Zh��M���x�N��P�X���Tz��Ś g��Y�ẻ�m�5 T��".Z��� ŠN��i�(�xG�ŷ:��Y�A��;��E�(�]��cNE�q)u��!r�6�V�����T.؝����PUP��D篩��9W� gs.F)m>��]bՔ%�H���1���72�_����:pЎ[�w$���uWzp���s���|e�s�I�7�QJ�xk_��F�P�ҫ�L.���+���0��`��rp��X4q�1��e��Yx\_�O�.�'�x��-~�{���!sTo�A�,=d�6���@X%9Ѳe���U�o�nLʼ��b�2��9�~�s����P�2u,(���I�FB���W3,}�G�
���5�1�u'�+��K��^؎��5�2����3X��|�w���Y�6�?����OҳubSU@X���0/@I5�����iԮ#�
a6�� 3:Uk��;�J�o�tEIp�(j����Xw�m.�68�9��X�H�t���I"���2T`R�_8-��ə�.�{p*��w��M*��4"(���v��(^���IR}���NE�Q���e�7�Х�6��+N�57��	��X��n+����o�G�̃,U^�pg^�����ϩaY����$����-^��6a2d��@-��wY������֖���Y�wmD�ê�(�N��B{L�(^h5�R!d,vXH��%��6y�|s%$B{����p���a�&�<`̧)�ȇ����8
 l��c$�	�&'%䫕��W��јE�gs}>�&�"{���������UYT�Q*٧�������H=?승�Yh�+o\m�%�oQ���nTϹ�P]:�s���`��1g�(���9�O{��T(�̠����E�n%��$%D\FX6�L4��PB򳌪" ^�+��������Jx��aH#���Y��̵�*X>؅U��`k�e����V��f��sd6����3M��Щ W)�4+�K�?�
Ɣ�pqu���/�I.��Dp�ڦR�;2��H=��3�|y�i<�g���3�la}���rkmD̂dG�����B-P�o�(W	1���H�	��v�me��
2y{;귧8���#�k�[D����:����[����h,���Z�i�0�y�M6��K�%��Ӡ�ܟA�p� �^>���w�5�"���)܋�����3�V����??�m����E�w,��2���	g��;o��O�A{>��	�u7ͽT�$ⶺqP4�s<m��746$!�e��Ǟ ���I� D?�=r�p�|����L1)",ƒ#^麭ڷ���W<�|� �V�˿b0V�J�Ԅ����y1�����|Db����B��F��gG@iE�N��с������v'���l*f��@,�gfj�I�x��E����"<ʅ�g�r��7���՟d�"�T��
�Dۤ�D��I����5H�p_g#��7��8-s<��X�^�1�HW���07�	���q����l�Q=57��ڃ9�Tt}�l�4�+Bְ%�==�EC{���E��R~\q����4s]5=�v�h�-�|��x��������o
YyL�������zm�:����W���u��(�����]��7�)+,"%���xQ�T�*���h_y���4���et%��s���a�NwBzO,��ꯝ�v��T�y�b�
72=}t��Ut *Y�����0'7�%&�d/a ����S_���B��@g�矴r��-��O6��G����1���4�B�'IQ��U�VL�<R�%�)��.܁NW��<�`1���5����K@���J���rqڅ�ͮ�FuXV�2-�0��,�r��x�umu��H���p���ٳ&Y��t͊���
�n���ۦy�f�Y_�g�M8�zq���l��������CQ�~k��� ("P7։�s��S�AxӔ�*-m�!~�NH��>�>-f:���frg��w��ۼ���S_��j��
$u�F`����ݒ��eZ��z7]d>��2�+g��UB��3r��>c#]lG��m��\N��R����͠j��l�J��>�o�*j=ƦY��r#ۅ�K����&TK��d5�H(z���3�bU�0w�$�'����^���z��V�9��(�
zڰ�(����K�nj8�F�jT9S�:;4��/�d����f-
���ſ��ݝ����5��)�E� ���A��Ds��3v��)#���zj�{�б��ؤ����\��@CXLu�����f�b�w�L!��?X�n�Ÿُz݃C��Mun6Rp6
U.z�!g�e�\WN�S�U����*�Yd�L�1|B���>�d��`"R�C@�����X	*�?DMLuqF	��dBG�f�PI9�=+!C&�Y�p�\kD�;�=$��iNs��z���u��P�t��̘\��D�S>����c� ?��9��3o,O��$�ڈ�C���	_n������p�6�P���cj�a���;>K�Km��ȷ�Ά�h�;Ox���mc���Z6�a"��=��]TĢ�Ĳ1���R�h���Z�n��7��N��s!����7UM.�[��TQ�s���(��Lgb����G?�S�r�ܼ1��@�:H��Vҽ��o0�ޖ�`�#5�tF@�~�c�n?�QS	�!��.���rbۘ�T-����P��Ә�<�j@�/�/&8��NP#1`ٔ.�L�o�&b��[f>��k`��m��mż�N$qAI��0��.එB����G?�&=_q�����AMt_� ��3:y������r~h���ŕG�g�`<����Ǡ�q�ĬM���d���i�P�\�[Bφ1%4넊��6|���<����A��;�����q�J����$�p���[�1�}}�9�?�_�&F���:/%PEyGE�gĔ�ڨ$Һ޶f��J��~[��F(�(ޝ�>�;�E�`�BU�DbW��V~�xl>��꯰�F�3a�IH�ӑ�z5�<+C��<{>Cb��{�／������)���GP�G�ʚt��b��^��ɾ��,H�5��.����ԙZ�#��a�XRH��e1P�}Ql��j\�tfT=f�X��}6!��z�J@g���NLZ\�x4��c2F j��_��,�#�I�S���x���0��Fp�G?�Ɣ��<g�����dO�8n	愑M�GD�������b�6�6���{�pA;�3
"�5C����+4�0�����-S�s2lc�7R��:K�����f��?��������f�
!�E]��~�6�d7G}%.���Td��f�р6Ž�8�8CM�뺕�6�X�!>] ����Ո��-6�y���y/�̖���ؗ����L�-ȭYl�j���-O��xB�ة?b���_�_hR�P �g[G�}�����"�o��2ى��҇.XE�[��zA��oJ]9�~8�+`�,udt�y���6������`�K2~}r?����q�P�:�eWH=�(P�nd��`l<�]i����%�##��i���Tz�
!�5�c�'�P|=o-���k�xhl&�쐼E5y%�,D����p:m�|��#D׸m<J�" >�+n��l"�(׏"Ɨk#��l�<���4�Їe/B����_9s��%B:'4�j�dؐ}�|��7�$/"�(&.6p '��Y�6x�{��r��C�(�1��q�m��Y��/J��3|�F?�0�����3����Q���*IrJ x���[������.*翩��(0r��o-o�]�0�ߖO�� iz8V��R�����-�2���2�3`$y48d�[p�	 ��:���`�3��e�ƞ�V���s=Fk��MeECY0k�D��qJ�Δ㙕NL<�ݨT��6���m*ei~������q��u^���ez\�B�O28/��:���c�:-�i���#���/�����nz�{�`�q��op)��ԃ��&����ų�}�F��R\��PZ3D��������25�e�b1�o87���Bz[��5̥���q�b�K��`^2�=�A���;")XN�Ʒ������CDB?a�`������:�"
�l��>�y�ew��0�y��'7�{�1n��1S�%�.Z��-�p�I=�^W�NFӅ7���<��A�%j�/��T���u�T˪^+%��yO���]�O�����74�[:�s���eۀJ��8v\{Nᮾnu�G�hJ)��krq���K
��� �i�k�W�,��Iw|N�j]3w�^�A"{I��D@"�ŗB�en>.�^��*�jsN�/��6�W�Wн�r�E]�Z���&�QkM��!��V�&^����.e]���BJ_/B���	r�^� ����X�!B_�ԛ�<�t݄��\�(Q�㌴�M^��@_o3��<<�(dr����
�̢�X�\O����'��4�#���Nb��X��7��n&�M�Ȱx��I���U,.���2�0�|9˸�����i?�y,ޢ��:��j�.Ԙ��zφ��9��T���t�T,l��YV���/#������}�҉�M9l��w� PY< ���ؒ���|��EFo�(�^�s����<QS�<���=�B�醔�ʒ�����ꘜ�d�4�_\YпVC�.s��/nԦh-�|��b�h�^)�>_H ⿱j��!���0��*�LVxN�?Y�;L�~w��C����D5�9���cUd�*j�M 2�6���I��a-p-ӷ0E[���q[ڒ��ޕaJ��^�b\��3��VZTn��џ�ԐG����]��eaS�J��+s�İ����7�k7�*�A9^����r��$/$z+ClUk�Y�qs�� NP���������(|�UN���m��R\(�h��
��v$�� ��,y[�_H��vR��Xo�s���z�^�8=$��߹���f6o���6S��5��20����j�Im�����d��\��7�:a���G;I��Z�������>�<p���)'�L��2�_L�z���X9��!�,@(��p��Ŏ�j��Qٮ��/A���YI�Rl�ߨ��{���#�iB;�������_#��}�y��.^�Ў�l�s��m�������}�#��q[kJc4d�މ�Q���¤����Q���+��=���s��P ��y��zz	R�]	F�w�0�zX)�#_K���nz���d��F������\�P-�!�ǿl�G�5�����b�>h���%����\��w���<��fe��h���o��DXMb�un�Ժob�'B�gG��I|q�d9P�9�؇Q���'rhԝu��?��Φ�b��@��������Mq�3=d�A�e���,����VX0�d��/7��H	�oM�J}����ZL��?Z�͵x��wsu.T���>0?����8MW<)��Nt�"�Q��e�y=�M�I��m���:���o� �h�JP�zpa�ϧ�����Qn\Ƌ�����Κ��z���vv5��a��
4	"*1��̨�`�h1�r��������V] �ЌI*J����;s����2�=�˽��Zږ������U��mM����
:�Α3�z���PΗO*9mMM%&�nMuDB��E��ی�P�� A��ϐ�����]:�+��q����K����T%�i<�cl�:OR��x�� [�������|�ǰ3�\�^�VP��kc�!z]�_}lۊ���ZxO��W�d�?�G�&��2�� �����ë�j�\�G= 
>���-�I�3�i�A�����!��S� `y�B�g(�R�#HEC�[r&K����$%C�$�-�Kw�����IP+��Z���&[��5�;�lBR^�^_!��s9`J� Z)�e����j%�9hI�`��CP��߳SE�P3�ؖ��_ț��7͎6��ݗM�Y�Ww�~�.��
*�ۭ�6�,;瓁��d���(F��M��Ң}���Սs�	����u�X܄�j9j6�f1U��2	�4�K��>D�U3�� �}I%�d�	K��P1H�b`��X�q���Jz�)�,b4�k|��w�RY��!�e$#����:߹4ǅY��.�D��RE�	l�)� ґ��?��iL��њ�k�VM��!���(E��7�6xk�K���՜N/�{�B���4������!o�:���Z�aF[Gx3�-���z��|�5�&��m�)2��0�z� �М��Ґ�^U9���Wq�h���z�ɅY�!*���}',x�7z�>�WK1yQ��H�ړ�*����� �#�qgp C�*��vr���-���ݩչ�f�;�	��l�s�hR�=���V�����oR]3XT)����x@ė�-_.!�1q(�����^K��#���ȿ��|-ĳU�je��3>���#i7��jsM�dFW�C��r}�|��g�מ'[LVso�ѓ\n�X��G�q丵Ig ��Vq��J��bl�Z���O��ǖ]_�{th�9��=����Z��ku��v��`uz���~��I[<|��EA&�X/�џ�_x��O<�C�SɎ�Mc*��Ev���@_�Կ�>���� @��2�I� �T����,H����xc5ھ�<����T�q�(_N��?�}��H�����g! c��j鐽g��[��]t:���l�<�Z�Ltk��Ԃ�>�Ε�P�$��@���Ū�Y P+�y����æM~���~ �j��UJLٗ�9�J�;��i��Ig8�+z�M�(���J�)9�U��;:�``�x�#��3Z0ps՛����i����s�]�/\8�%Ή�h_["��D[���x���*��k���Z�;٥}�ic��ޕ�G�6�x�Vs�9f��ֻ��̪m�c)X��3��z���_��Qq�g=�?v��e��z�YUEC�DMG4�Z�Z���#(�|U��ْ����~s5�Au0<��7�Ģ�����&$���y��<7��/A����^/D���Z'ۛ��p�S�b��3��a{��m��Qa��������9$�Ԁ9�|�N��]�v�[����,јr��/�E��px�Q5m�Kk�H]�����U�nBX��~R�hQ�:/xN�w�oA�j���G̖(+<s8�=>%�6�O3���=:;hFC{N�Ƅ�J��C�����jkd��q�� �Z�>��E����w|����{���v�F�[R�.S�ld�t����X��.���z����X��(�z`���&6l���/1ʆ(Զ3CmT��MN��I!U�63\��6=�|�b�tʳ=����KA����ަ�.���U���T����	�)d���7r�Zo�r����LC+m�ͼt��Uߪ�����~�	�����=։��F|��k}�3�M��E�¢^�'g�~y�L��K˷.��B��-:�5������~����N�^�X�
�ó<bQ������I\�q�@�r��NG;z~W��c�8mG��)n7a� |x�s��I���A�]J�{I&jSc�'2�쓧��ޱ�l,�(������Z�\��oW��5��3Uy���ݑJ�)�����kV�k-�j0lb�(9d�v���x6��x7�s�"�"��@���m'�����m{���7�z�琐>"�Ya��T����x*6^'D���0��R ��s]��)N�?.�����R�IZ&��o3�DB�҂7�8�*�Oi�v��ڧð�����C���=PU�<_L(��%����%>,���&��
�-�t&?I�ޕ�r�:Yޤx���}��*,�u�bp
�IgI��T��(񉹠~�g�����$Bᛩ�xq.d�&�����l�~}I��fչW����jd��:�~�;�4�?P�:@�Z�'[��`��T��̹��B��bd��,�l���U�o��FJv��b��I�������d	'[��4e�P9�?!�[�P��|U��A�A-8���k�.�N�V-���C�ėL�����9)��aN��+;�\|���3�-N�=N�g"���[��so���`�Z������'/n(X(QR�(E0Ɯ@������s@z�
C-���N�ƙ������� oA^��y��ہ;�[�گa�B~蛬!�-��DG�{@� H?����đ({5?R7��/8�ѷ����?�D�џ�_�^�xU.2�B7;�)�����M��mJQȲ�n������f�"~P�[v��w���ۨ�|�ȓCX80U喐mK�#�.��U����A*g� ~^d��Y&x�8���{	/*���3��J-�\:��5��z�2ڡ�`�M)^7�Dh�%�z��� gR���8��a��|���=C݉�ܸ��T�����OM2�ӵlZd�К���Rפ�ޕ�����T���;����]���~ݦ���j��l��JfYг~B��a��Z��ȢN��0Ca"�T�=<bne'�=�{��`!;\�[weyH��z�s�aJ���oA�Vm�zU�����{��;��kA������.|�IWF���l�G�ڞ+��-W��(DDhe���Ș TEG���E��JTj"ؘ���o^@m�.7P�z��k�6�.c�y]�k��w@����̔2����i�	�)V����x�-�U�R�͘j�g�?N�Y}�����
����^Դ�-e�zV�hg$x�nگ�:�X���C���%�p�>l6tv$��JUx0��x_rn�y3!������������yG��&_�5!�\3Rm�o�n,G�>r��}"p��xI"1�i��gpJyT8���|esbHߒ�{�it(�zn&F�e�5P༄��1�Z%y�e�׾��r�i�L�NX�&1�V�h�
�O���3��R<�(BP>[\�~��ή���ԏM�}#�de��Ĩ�f�k��Yii�|l�2yf�&,���Tھ,ky^�kR�&��,�{�ɩQ����`��ȧ��;=�
���.+��^�fEH���Cn�L-�n��V��9ds{!�x$2pHǓ=zN���J͆�:Sv�B�;��%�Y�
#�>BS�6o>(%唸�z���e�Q��Hr�/ݓ��H�p1���|�L�p��D���X6��|&B�$+�S�sʯ~,�^V��о���n����}�!��@�T44��»$�;F	p���6�q���_ͿA�a�Av]_��N-�K�:�-��8P}Q�o()X��w� o��%̃�����	���.ؚ�����BM���Khw���E�*�\)m�$��.x���a%��dk4����h��D}��Ј�&�X��,97u�A��ĭ����NS��m��\�Q���-��|-�l�����=����,�n�l!Y�vزHk��i��vP�����oV�)�yַ�=����5,Ǐ�s�$GkE*�s
rH�䅺PF]5��ǲ��7�`����ɿ�����g���vmL�����4BHr�Ǣr!A��������w\�.�����r�/2��t,��5$���Y�sF�(�k��㮶t�HjBhwG嘥$�P�UE���P�.M������D����,�׶-0N��&
��e��+W�"o���e�
!�h���䁚@�����@�@��S��<��A���H�2�����5�d�/��(�
Q�f���:�v�m���$�B��/ {��a��,gwkPϓ���:��7����nF#@��W���g,�h���r�E���%��ep��FS���{� T+�LD��L����%	��YE��I�J�8������=�%�!�u>�w�$-ŗ�����Iǒ�Z���8�3[���P|�0�'9��F88�}q�Z��$=<XC#S�~be$�:i���4�g��Hr�@��J��F�(PO)����sB���S�T����.U�P��s\u��?to�o�$�B�>�D3��ER�@<&�2��؏L��D���"tD`�TWh�.E�}]-�.�E�[�3���d$>IM�6���{o�W~�,���#�^6�$jX�A�������E̠��p��v�
�!�rz�EPO�j'�!d#t�`�w�JMG)w'|�����[����A���n��D�B�'D�b��P��T�F��&2�3��4E�q��g��pN�[[lrt�!�gS��r���:�q����*�����p�#��l�RH"X����i�g���TnYV*'<���!�v���;�Y��=��Mݷ^Q�if�;�������Ĵ��	`7�N���M�S�&��f�����6J�������;�s���U>��~�1�S�}JG�%N )���Cv'��\�s�LW=PN���	�m��q�M��/[��ǖ�A�������+��EDژE]�o�s�͒=��x'�Ê����	�1�	��7��+�-��0�s��UoE�T�a�M"��D7�����>���z�j���#9�ü���^�-��1AR햞�M�B �����L>��+_�sj���O�R�
m�-�*�����ܾ���7����-��i[a�0	�w����,=EuL�OY���Gw9"��#��Y�:��pY�W��dLB���?K-����@��:���ؿ�%��M���"������w��	 C��ʘ(ϊ/h����^�����Q?���7�ag�0�bqj��ɶ��	=�\���G	P����l� �=��� キ8O�!��<oR?�_�h�����	�C�R37�)��p˴"R��=д(�ǘk(ح D������`&�U]�}�UǨʢ]6������d�ZG���޺p*.��n~��C�F��Qu�;.'/��HΜ��m�G�4p����5�&|G
͞�%��d4�kD�'�e�&:�Ds��	�la��%�߿%_�/"��5ј�׌+��IxRp8�[&����_jug���N-FWSF���wI��.�)��t�����������z��K�9_ G��y<�����j���=8vU��<����L�ٴÑ��e��0�cTU�������#��Egr�a�0��5ṉG����\�n�T��6�Â��:����r�_(vU�Ҹj�}rPޞ�(!�������6@�pz�؃�tQJ*�����mk�W>K䬕% gMǸ�[�y��\��l�ԯ��0�D�f��=��>0_徥I��یk��l,�QU?�qJ�\�s�zS�_���8+��9����� �P���ψmS�E�&u�v0�����ڈ}�� 8G������@��1����a�ɏ�C�������ӿ*��vT�R�͓��͙�}euت��֡{���T��9i,�PWk�7dCB������yx�coG;�X���ܚ�*	�9}�HN���������`Fw����{��\��O���6ZzT3�I��{�F`�(�?|��j���zK�
 ����	� ��_/�*�7&k:�̅����;�*'�&F�E	��fW�>�k�n��s�D�����Bf:��@_�8+�8O�mJ3��CMqH����6�Q#1t����m{<�����UL���=�i�:��Lr6���ѳԇ{��r�ҕO�u��o�+'I�4rB���JմP\��'��L��/��M|�H&A�*=�2*W}�Z	���B,�5���˩��=�ll��m7�7�����]�*�i�tZ�� fݞ����;�OϬb:�E*��jz���Eq���Q�n�3��|�zY|���Q7�}S�Sw�fE'T�G�U.1��9�a%֜�f���	���]�8綽�f!��C�T��ok4&pX�X�p���(5"��j[:������@�,X�N%�ມT*��U�ڑ���|�P�z�t"q8 bx��U���	U�d{v���;�����1Y��f?+����@E�k�}~=����4�t&G��wkޞ�a��ʘ���TɱW@���͚��6��#���Υ{�������-;���%sT#Ƣ��1��I�<�4I�K�KV�PS���`j0P'{8���!&����\A��1i�P�����Z��Ĵ/;�gA�m���(C�y�>�mJf�9�2�ȁ�֨���Y� �t�"fO�(n}�Nl��;.�\��u񾾪bZЀ�q[��lJ�!��li��S��թ����BP�A��×A�2���Z�x�>:x�wя���XB���}q�Kq�גPy��$�Bm�"?b;���a2�od���SP��w� �^�at�x�d���O�Y}b��b�>�S��J��� ��M�Ev���o�&W/^��!A-;���! -V	3��gx
¸/��Tq1+�x2bF0���!��6D0��{�hL�2�"������vT5eĊӪ����oG������c|vȃ��޶�%�I��46^�q��]�^NZ/,m1Z���)�=�i�Kb.I�:e��Y�$���V��Zu��$UE>�H��k0ܙ�*���rn�`�'&5���T��_DT��T�ֺ���Ǔ�I�fL�E�@в~��W�Tr�w^����� ���B���m
G����6Ԭ�ooY*��d�+Oe��T��q��pﬦ7�C%D`L:��L�X�/����"85[�E�0=�)]�c��Js�S��:6��1Ϩ?�;儦f�a�s'F��-�j�e�"����j�� ^rry��C撬H�����麘R�1[��ݦ�Ւ���~�V7�����mLaG]w}��)��N��cD�>i�N��a�#�=�H�{��1�!e2vҊ��.��7�?
HD��|l�ҹG�I�Ž$�,�3S�w��\/���z���P�L{s��Tb�\���m�������ΰy-�DǙߋ;*�*���[]kHGt�p'��P�9o{�}�����!��r���B��r��>���J3�M89x%5�]:�������3�(�Y�5[( ؗh�����S����4ޑ���7�D�K>ſВ��zA�
�Ls��ͳ7�!��V���������B'�������z����iRkb$������3b��o�~$䆛+�f��--�_�?/�vщ�n�R=D"�
D<DXa�~���z��6��m]���/(D����Fz{��'�f��y�\�N����\Y)��K|��I+3����.��/]��-�bf��?oT��}E#�E5��� �K#Ou��y2��?�_v'��;�S_[U�(��0(�9�b^Qu���r�����ٺ�C �'/S�V&w�覆�����X�P4�:�H���m��#�%m�BM?5g
�%)oט�k5����M�` ��%���5��J�scλ[��6'��냆�[q2:�bZ��)w �}��cI;�}vݦ�D�d,^Y�$Ȋ���D�	�z_w��kP����D�r;�Z�( 0�gע�
���1]{y�5N�y��U�DW]�H�^�m��,k�|��J#r��(�3���w��[�AF�������f�����X	���&���埆"2u5mSz_�Pqk6;��6W�p`DD�=6к���l���e�gmnV!��0�d��D2��1g����訋5�%oM/5�V�db�7~�?i }S&�c�!j!�*!X��2i_O���#�#��;���� ��)���Ӡ�n�t�$	f>�(���/�r,�7�2�z�]���!Q�Z*�.�N�d��#+d���/?|~d���x,����<1��^����L��?j(ahY�I�=)������_��B�a����a�]������ ��$�V_]����KIUQ٦gT4�C�� ��I$�A9�Ӵ���&bj��w!o��rH��=("�ߏ_#Tc;?��8$I�W��S�>K���ҿgc#�Jނ�^���H�쐅�m���8�}Ų����L{�_ ~8^��;vن!�m�pVB�ӼW����B�e��IM�v��I|�oK.���4�����w(��b? ,G�H�����䅊���ĸl2��1�_Fϣr&9�㩂'Gu��Ϫ?�Ͳ�#w��0!���ƴ��qvF�E����u5�é:���6X@��#,so�[T_V�	RG0X:B]��_������c+)�Y>))S~��l�ܻ ��@��;�Ѧ}���C?	��r ��
���~گ��y`	EM��ጏ-_VqL&!qZ>[��:ۢ1Cu4)_%�������t��7��O���Q�ue{����E�
싪��!���iZ��V�(WBh!J�g� ����5	*�jF=��y6�TdX`���˅J��J�{!̤�64�p�ʸ�3��9�8`����O3����;�+1���� Eb���W��Ͻ�,�mM��=�E���V^�)!$h��6-�S�È��J����
��9$��������c0���ȪA3fՖ[�8�T	��Fr'Y=����!�X��d��$u��_�$''SU��{��+O���3��=F`��~�ՏS$�D�yn���}F��7���C_s�0C�_%ь�9;�1P,��@v�6(�S�t�ш?�u��?�jc�	��̱kG�������s׵J�:� Wé-u���L~��TI3����p���-�^S�s�4�z����n�#2�}�,&�N.WU��@h)�-$��|�WΡ��奍�-�޼���`|6K�� �Ṣ�ҋL^L���ukF�XJ(��7m_�u���|��>3w<�1�Z%���j(1E�Zd�7v�iZ�g�^�k��p$E��o�qr�PPmũ�U�,l"a�_Ԃ������(!_2��b=`Ay�?hG%�1R�h^p}s�(�B�9I���Hp���nRq,7"��BɎG���x�R-Kښh5��@�����{=�h��D�&�����D�����u���u*1�|��2f�n��Ǩ�s����d�(�>/ru��BK0�T��b�+��J�~(���(�B�̳��9߯P �w�o��̿�W��&� �^�.V+�����wȈ& "��9t��e�Ԋ5�T���<���m�]}yx [�ޱ�I�Jb��9�!��H|z���Y�/�O���h
�m���ذ/6W]��0���g�ًC��	N!������+/������ҀSwb�dn�A}r)��
ʚ�yo޸�%ND���<~n��qZ��𐘉/>/����c��(�4�w��R�0�$&�ԍxPߝ9��L���;5G�X+�8�3��H�|���O�"�&u���v�ɏ��F�ؓ?\�!~1j�[� v���EB5�]Ɓ���ec%ʂ�PȒ�1��v�F������^=��|���d��f
��Q>��[(iX]��C3lޓk�|1$<F�cH��E���u!X��Ռ��� w�Y]��~�Le8��
'����P�=��Ӥ��3�5����Gu� ����R٤Oc�A���8��>2�mf����d�`,�:C�c�!4�1x[�����X��u2�1)sg�~�����('a�����u��\��e���
�I���)F�i�|w����_�^0�Z�QN�	��4]u�j�
rL�@��tO���.�I��.@��^}?��.z#`Ѽ�;TZ\��F���a�i!�����,�j�?ę�0��o��~a7��Y�hkdN���W�P6��!:Ll�w ��Uo!�e!y���� ��5�b#y��V��'����ڴj����n��A>Q��]�o ����95%��Z�n�%�S"�Q���Y����us�9�e,����X���55�y�J!����qݨSW��-�*�,��'G����BlBɜ�B��Ν�&Q�Lyϣc�҇+�X��C���@V�4;!�_�! {������S|*!�̴Y�ƶb�t�]V�������L�}�UH�9��`�P� p{�Fx=�_U�8���5Y���1C5���a8M�Lt�ǒ(Q�QPu��9)p�k�0������������6h���R�H�?��)=��=?`����>�Lj�bo[4��I&�|O'-�J����	RX
�"-����;?(�����"����h{��`3�Z
���n-��[�{�M��:���9bn��A3=������AOt+XԞ3ay�R�s�?����:fT��ɾYՕ�ƊA3�ʭo���q�tM2�ڜ����&�UӤK�8�[�I�t3�d���Ӂd+ȏ��Vό��a��X���>K����-�G�O�YC	(	����Q���[�N�Zd"���4
f�MZ<ӧ�?i6<���)P�bx�ct�-yi=�H'�����f���ݔͪ��x�0gC���%�>c�a�tR|6������G?*y	�vnw��Ғ:�����%�|�`�J��Ɵ�Hw_��g��=�d�auӔ���M��'��v�(B%-�����@�:��塪{i�F/��bV����bX��F�P�wѸV*S� ���~wJO6:���r�����|M�[�q���Yȣ�G6�	`�"돌~^�o,pV���o�%1�+��vȾyB��d��Tߥ�Ѵ��\��7^�7Bh����q&��mY��k2A�y<s.̞�4Μ��)�H�Y�eM�M���\ڹIؓ��	�'�o�rd�V��X��{�!CB��ǤA
L�;��I�M4�}FAAc�<���_91mX	ʐ�T(�@�(OG|�%�]������1�i�v�D��
��IK����c ��D| �����v���x��Z�׃��>�/(: ��D-~Q2� �v���7o0�4�GVT����@��Z<3�+��rY-�G���	�J�»������2����yd��Q���Rdm�EcR��C}���o<��.Z(r�ĕ�e��v��]��{y���԰T���ZBT��<J8���p�ư�H��mp̶��w"�Yi�������Yn�~1�h����H\���#��'���4�A`����%@�����{uv0�`���R�M{D�(R~�f�:*��#%1Lp�(:��K)2P�p�3�I�w�Opct5����
���R^�AqpY[
��1D����t����`��2T���?6bMZ��#k��F�Ls]��,�����/GE(���6��$�.=.�{����[�L��$�{� �Dj����`t�=� �:�d�X�&+�6��l��{�cߛV3�Z�ק"�=u�D'j����׵�l������Gh�c�.�O�Okepa�2�:N�����.b�G�
���I�v����BH�|�;C�%i���)��n��*�2[ù��t
Q�Ќ�����y�Y�;SS ~�Z��r\���I�	.����3j��ڷ5��3sGm�Ӥ�m���9Z78�`31*`a]�Hp��]~����0.�mvV(80qt��Y,K�*���e� |��6}W)�n`&�4��6,w�����.��)e����~��ƀ�&9^�Y�//��������P�T��v�s��T�j��W�{��vgC[x��G<R��rr�a�;�j�)�n���-��$���e��X��O�n���M)�^@�0D�u�2��4Z�J��z�dFͱ�x[�-]o����z�C4Op[�j��KJ�� :��#BBB�����������-��]v��	�^�o���m��t2+�꣓rJ�<]݌T�Ⱦe�+b����4�|����E����8�}�[➶s�1�o���L�����>j��OD�n/�%T7��x/��9��^_w��w�ц:a/�'~)��T7B�y��aq]�rZ��� &��{e��Wa��v�;u��wɐ��k�W�n\�+q@��u�9
^GZ�^=ʗtZS��8�a
��7��\���6���c�&�Ķ����`�b����M���Q�Wc��-_Zkyǟҫ8V7|)G�����Ԛ����tH7��
=�.
^�;���;!�,��3-Jrۚ��K�&���7�br��H�k�e�#-YwB������]��ʁ/z�p8��*tgS�u���ml����&LFH=�:���$��Z��ɮ��6���L蕾���U_���R�)����+�~2��b��np���[�+q0-�2�݌ �N�Ӱ�ʓ�i��"ғ�����S��>�Ԡ��*AJ�rĶ-��&��As�g�S��gGN���&��.l�^>�u�>}f5��L�	����^!W�3s3z=B��w��+8�����9����\v�����gE�V��Q'�Тb�AE塑w��s@�	�&9WqX����߽A;�0Ha�0�:gy)�/�W�(d�l�m�G�"w��A�̚h�Z�=�����rH�.$$"��;_��4�K)^K<�E���/2\Ӡ�����^�`-�gI�U�W�qT��օ5I��<*_��Q],�-�q>�2�����R�/�ҙRkS=rH�\�(��a��G(�J�Wӂ�; ��O�C�z���q,��,o��Y��<�b.f�|Q�ܢӋ�CP$�B+ic6ZJ�4C��uq��tאQ�3��hh�vU���J�o��o�/�_8������MD�5rſ�W"v��L���j���i�P#Q���!�n�/ �@{�߶ٯ�L�����{+�{�<a�2�_��	{�,��4��R�8�u��3�p�;X7�Ƹq'��ko�_~[�F���!|�װg��m"J5��4:Ϙ1NE�'�f�}�1:B�$����`��H��Je��u�oq
��i�`�o�G���K�>-�+J�2ρ�{��l��J�U������m]1��a00s��oS�j7����C�/�$�ȥ�j:j��=2�d(�.�`�+ᣚ�$E����������V�����G�w��Bh�:]i
�?KܻY��F�Ђ��k�U��}ֺ��Fϋ�/�o)�x(��!�^Xħ��Y:a����<��5͛}��p=��ַ_�����$��:Nj��o���(�v^8��4ny)��~CO/��!��Zm��9��TMw|�&J��CqNfc�uu[�P��F�$Ha"�F����xϳ_̸h�3?����K*S����vda��������B���+n�Pwh��&׃q��I���^�ԡ��'����,`^��h��X��5�1�HѾ�ɷ�q%�����~�$���h�YV�����PO4�m�)��=�L��K�@�>����`��g�����&���Q���Ab~m� �K6��cͳ;
�G�ʨD1#.�~,ߧ�\j���sd��P&,\w�*ؕ|�\�q^� �-�%���Iuy��Q�َ��Dd�t�����.�3aOHI�/Y��J�P_Z&��C~�zb�?wxcQU�j�Y;���	�J�?i7gV��t�̫pS=4��!2vh��~��y�ZB�D!��,�v�J��$Z3�1���Qߖ	���ggmc���x2V|��P�� f!E)M@���|
/}qHMu��]la#'��,|t�^;t+A�Km-��E_�˝��}2sϙr@��$�HJJ�8pZ�h�BI������0�;f��H� ��_�R�����w�Q��rԋp�2��u��y��%:Y���y�`$}��D��
���^i\���&�]�Dj�g#q�G�  V�>-���=�O��Yfp�R�=�^���-bٴ5��.��_̺Rf)����m�=�i�J�|BĶhf�Q�/"NZi��]�ֶ&A9�j�����Z��_�u V�&ĖZ!��N�ۂP�aq��Y���g��V��jhtЃ�+�鬻X Zv]�tr$K;����cE���������/C��v+��ndF����A�n%���x�{[��&�~� AT��e�ӵ硿"�-�Ś7-�Կ��I�|U��Z������_'�߽s���	�~�.yk�ty��p�h.x�.�չtD�5ئ�J?�U��C���m�za���Q����[��1u��Dh�� Nq���/a���`�[���ܬ� ��ۥ�z}FA�Uɝa�jER��%B�?L[��/ݟA8����m�3���ǝ���O��ؙ[��v��1���6\4�厶m��12V6�o�RL}���6�P����Y�e�ꡌ�-���n`�up��}hu�;�b c&߇B���1m�l�Dxѳ6�Gň�*���֮�_���c"��6�L+w�ѐ����� 	%Bt	ȋ���t�#��vJ�G~��j��l��i5��>|�b�9��w�-�@n>gd�{�{jM��;�z̔Uʭ*'

q�{t*|��a�.=;��q"Ah�G�sfK�l<"���ǐ�d���+v�{p��_C���8nמ� ��R[���Y��8LԌ�yt�lg����[��^f���/o���Rr�u��$|�.~�����*}�#9��J�3�W�.t/���N��{>��yq;������qoY$9��e{�X�{^�k���P	I쩿��D���|y��s&�`DsLQ���<Bh�L���2�&l˻�7¥��̺#�N<���+�5�u/��h��/�h��?C��\��B!����_���l@�K�{���[��h����ب����Zň�%�����FL�/>�p~<��9���+���E_u�y�K��M�Q�Ε��O3�Z�����ۡ�����m9��9|�R�
�x���p��K�J�Iw�vʼ�\GI����}
npл�+���	�
}η܍���#��ã�}!P��&]�xſ�|���,�����2Ŕ�_��_�n�"CL�a���c�tO�˔��*zR���2 D\1�[-��H�E���B9����P���\���{f��K��v�|����j�E9E	8�Ɗw��b�tO#��2jt�OܑE~��
y�<A�'+��v�F# tg3Vapnqw���r��ЈZ3��@6��7�"mrd��#]�v�m5���,!����}`Y�S��H���z�*I�	�[�7���z����&.E�M<�,�u*)+�j8��2�-�B�S��8�?�����C�_�� Y�����P�sj��P�?�C�����$G�%$�6k�g����9�9X��Cq$<iZNC�a���lL�u��1Z�B��h���� �#.�I׀�2�i�@����!����q��)=��)>s�q�!�e��h�5G?�Q�6�(���c!/���h3�1a��J�T��|�u�[�楕'C��7�@7s!#���⎴���y��ȯ���P40��)AGH�g\(���Xؒƙ�2I4�X��?���۠���1��Xl��?�����F���f�%�*]?�$�v�}"3���&���V��Bpm�1�h|�z#	Ҹ�p�P�!��f#�[ �*|D���D��}c)L��\�Cn�&Q�,��?�5��s�[�o��[�JXU��sK����א���yQgw�`s��`7D>	�6��1����-isnk�{Ib>�?P�5l�hLb)#D��͐��i��&~7m�����;18���˨u"�~`�*W}7]ïLAu�8�(9��2� �
���7&����~Ȕd=�����ѨʅG@NJ��j�L'��9 g�k����@��{��@�+J.#�J�~�4,����g?!o�ۑ�N�.�W�)Dp7P�(M��'v���4Y�p>ͱD5�'�#�3|�	��]��G43����^��,1
R��$�}^���ԣv%���mYPD�w�>�,}6��d_�$5x/]?�'`�	@Ɍl<>�]^�`N��k;=m�I}����Lzɉ&�E��hK�lzvЁ[�Ҹ_�!;$�z2���A��M{�`�jR:A�i�/�P�F;�+��7g&5;S�ê���w�,%/+�A���4-&�c��"�D�Ȍ_�&����"�d`��C��P�CS���@�k
�����5z����_�O��e�(
�UD���EIP4���'LX�̙��q�~0l{y��MG�����Ց�G�y8�#t"/��z�`�b�@�c�8�Jz��FPS�f]��H��������0�֧��J���z�U�pN�$� u�&�����A�x�n����r.+z�#Y����ī8F��g�/��D���f��5��4L���m.ie��ҩ${~�	]"y��':��= �`(���cwk���s�2�#�&z�Y��F7lCZ�]�]���ڠ|�a:*�^������+��sF�lK6�RUO4.���f�k=�����L�l�1I��B�5G��v�"Ģ�� r='z�@ɍt:G��1c&�9zD�<��_i�?�ܣ�Z��E�'Ea�������;p;*�n;r�휚t%K���/�2гL�I��7w8�!��G����$b������tV�e��qP`zFǬ��4"z�>��JK~����Cb|xc��H�2�]����	�=9KX@|��-$b�s&z��0,9��� =�����N�(�5j��<CO:-�?D���4���φ�ǱU�O��S�e�Je�&`6dˀ�˼���7qf �4j�	���ԝg	
-�9���G�1��B�����wCQf��P"6�W���l�<�i�GTW�����X��j q��D�̎8*�k��a��h��&�y��uV����`�������PO�!{um�JB�(���Tä9��T1脻vY��WdfUZY�q��j���"a�d�
���|�E}@����U�
Mg+[կઘ��d�V���O5�,�a?���O"���O1�k�xw��s�woP����������Ӝ�Cr��c?mо�[��U#̓j��,��g�}�?Az�(���m��Ysx�!N5IZȐ�U��ݻ��Ґ����<���Ung'�˕a�cR� �۸���vk%c+��8%�g��N��y���7��@�Ph�r�h��3)���tVR~@P����ڒG4�:��z6�޽�얨�r�nr=
�a�5�ՒZZv ��7�t�r�T:/�S�W�/a�5�*�Re-�&û��}k�q~Y�	����6��w	�l�y�b���@����rV��|��s�/�f�u�F��69��n:A=w	��>���Q3&�*[�h8#�
��[T$1��.�U�$���c��8[�ढ़�yYS�r�W���p�J��~o����mb&[�B�C�r�Kj��D���E��Uﺑ�(R�#��lTG�&�Y.�K��Èsf���2��f>����Cūg������&��N�V-��ʗ�Ğ����&�������rF0�`���D�N��ebXE����r��
w�-��z��'���~ބ����'�R�?G��|�!����[��c�L��^�'�q���LH)۔��US�9�q���X_���z5���s~uR��sY�A���⎶�|(��`�F�|��e^/�_�{"�d�%l<�F ���P;twÏ�|W aȰ�Z�K��.�7Awrͱ���G9�Ջ������f�lˣ#(�M��[Dt]i��6��oB�����G�Y���_���ooɟh�����L|�զ*jV�� wĨ��E�����ߏT��ޫq��q^݋�E�ݱIMب���em�<�@&Wq�w��`�x�5�#��`��"����{��/[w��mN��P$^���Wt���+�#�,��x���0�A���f{�w�1d^3�~���4B�$����#.ӵ$a�����ZN���^~��&{&pȭj�F�P��PҒ�*{��l%D�$��i �)jk,��.Ve�Ѵ�č��ḉQ��5�aN������G�{�l����s'q��1���¢�2��;�%7{�ƣ��T�Z��0 rf�D�����RO���}������=��{=6{��H�D���?0�ޭ��o0�����ʖ)�d(��f�rDf���5ģ� >�z{r8q�:���j�m������� ���Ɯy��[��ѻ&���=�X��M;�~�Bh���S��3g?����X��%�7�<�'_@��2��BmW�ϔ��๯��:�6ƕh�t��8�,��c��K�d�k� ;��
e�x�D&�K��|n!h�b��-2�UE��t��p�����uvdIѲ�L��*E�'� �M�%H�J���ٰ�� i\�=}M��,+:Ja���o�}߻���JZ��E�}��s3�CT���9�r��!�h3ؽ0��ʄ/�,4ià+b7��ڳ��[KÕJL/��[���x�Y���`�C��K_\�}Z�W>LgEZŉ�n�}}�鲡�hh�u8�7��Ղ��������I6�ڬ�����W1Ax�<��B9e��BZ�����E��!P(в�;\0�lk5+�����TM�U:@���FA�h������~d ���b�.�<�Fqb��q�d�1Y`mʢ�Tj:��h���z��*��Y��yL4�\���{vTZ��~�IJ���<
���W�n�?R����V�"R���|S88�E�����̅=����I��$�Ŀ�����u�s�%A��m[�c���y`�d�D����F��Fr3V_��f䃮YAf(� ���1,� �2�y�oR��2��")y�����uC$=��X�W��4��t�7V��1������#��.~��Gܣ���W�
è�.<�$$�o"��5;�G�6��C��5�e��*Z��$��g3\�bM�md^�U0��RT����6�U���~��������"����*��Q�5-@n�J�m���,����|nek���^k��w�5�d�R�cќ�1����a0]�ou��}�ר]qs�w �����������L���G//)J��3>�����y/Ĳ�p��f@"�E�z� e�s���>5{/6Kw�aɡx�����p�0p�= �q��Y�&���+���@ņw�J1\WM�ǒ,�X�2�:��۩�.��X��;���#�-��#�1`L+����@�1�g�|�r9���=4�9t�� ,��.
��˱fS�++��8lSe}m�6�w&�Y���"�*NZl���.�p��<9: aZ�_�l�wv�r�G�����p�iquV/� �n_�~�oE�defX��u�R��*�H q'���n�����xD|�\o�U�/��U޸�~3�M)��s@�*δ�I{�v���G���֪�	�F��;�ff�_$���x��>�0���\}1	����Դ?����� �qc��|n�������S�E�?���ֽX����| �	_߼��J��8q���1"ł�P�pp�>���@�B1������OD��ψ����/�.��4�U����s
"��;2�2cn�Ke^[KOnmM��R�ԉ��S��Wt\h��u$�`��h6}�k���)Q��n/ƝY���Ҭ�LT�Z�(��P��8>Ӓ�TV�����
R9IH'^�u�J��������\r�*��d;/����o{M|0/�����$';BݍjqO"�]ζ���M�(՟ǭM_�ɟ�����S���)��e2¾A|��q��>z�GZ˿\���8|��[�	]R�B�v(�Ʃ�4l
s���џI�����B�w{��]��!+�կ��H��m_�!�P�D������i���Yh��<xd	��D�R�X�x��oc^������:j�5(��Y(��X��ՠf(�h��_6ǖ^��'�G��#zf�X��z��!�-,pF\��5�-!��6�X{����v���^༚�I[](�{��
p�^�.�F�zr�8���Qׯl�$C�� �{p��O�{�$��_1�%����~��ܿ���Q����s���II�f~��å��u-GOD��P��jh"��Xi�S��I�I�)�a��Ə>
��EH��=��Q>|#�.�� ��\ێ��3D�I�� �E&T��N�e2�3�c���KK$�4���i�x�ME� B#���b����D���G��A���	wrSR�����	��sP(�~�s��l�@n���b����S֬��"x(��B��bt��~p�z�ϋ&	��Y����}D&�����b���3��X�o�'��{NNOsH�ȢC<���?�|�!���8P��,DjYV��g�C�.6H]>y��㉔¬��*���#�fB� U�U��8>U���� C��/UT��G�He��۠o�5wx��F�u#S�����)Q�!??�0{���G�:5�q���Ҏ��!vO'|y����$����w�d��Ug~bc��2����e�KH80��9h�x�p��Aj:78��h\�_P��N����{D������#�R����1dTs)��ٞ��*QL��)3NZ8��H����w�h�˓X���:h#�� wE?�����ڿ���܍�2`��G&+h���~Z=\𱕩�ߩ.�CWo�y�m�>	^���h0�r[!a.�P~���L�6��f>��9	��*P=���9d�8!e�g�mbR���ߜ���X>��ai?^��� ��YE����5)��<��_w��^=d�����A�}���2MK�~��G[�QL�Y���ݤ1���z����6�K��f.�Yi���YKXu��$3�񾇯�6��>�b2vI��r���RQ�6�L�D���eY�,��n,L2��\�|A�2�0P47ZL��8܅�����z���S�w훖,��4U���~Y�՝ol.+���+}4`JU򣵁%��8��d������Hi�,5��;9�q(Ɓ��"�_u�|!@�N>In� ��T�����4G�V��i���&�k�>�n}H�=R�D�I�[3�m���;n%�ֵ���S��T䕯��@��]���&�-�[/Ͳז��E�A3�T�1@h{$�D����Y0{��J!�诺W�:�^�Ba&�W���@zsei�a+�c�9�x2yt�-Q >I���{�^	@O�8Ϻ�sHy*"�uN�M`�1��zVMk�.�,���\�}����`LA�!κS�*GQ�}��M�wB���HQ~���Z-x	 ��.���7���#v=�W8X���OhM_�"�1N|qw٠[�������Ȱ��Y��]��m����7$�v�\%$2��/���ս����So�/�2�딕��l�:ިe8�	�1��7<��F��(�G:jZc���5G�\H���(��� Y����Ԏ��"詮M+9��#Q4�'o��w� ���>_�DF&�f��	�*c�k{}��e�7B^׮�"����<�ꎐW�Eg�{ ̙��b�߁+Bv��~��'KO�On��\����X��!}^@��R�Q[�K�z��bY��6�jVO����	�PtUOi0F��N�ր\|1�@a��6�)9̺+�}o�A_�\�'�����DdE���j ��66���­E��$#P��Jr4�%�w��R��pMj�$wcQn����NbB`���}:�d����Ȼ�IEL�o����3�i_`��!օ�AOn�Ӷ��0R;_l]�DG�Ah����]jsE�r��
����<&��Y�����TKE[{sϐ.���� �
i�
e[vo)��T%���Ú�|�d�p�U$��%W�֙
�v��(��cP��c|�~��)��Y���Z��M�,��?�"��+;]lq�~�~��eb?)ŧԺa�?V���H��Kd�Wd2�uqi8�GwѾg�ȕO,7.4�t+{���Yꆘ�L�^� /��;���	�
k&���_v�91�"z�v�X��IH����Z��c�|iÒ-��d��NL V�g2�A�;��� @� ԓ��_�qp��zX��N��k&:�5L^j``��E��R�>��T������3�ZH�CFӚ�auM�:'��p�����B���6\Q�TO3�߆ź�:>��Ӷħ� ���t�q(K�{@�������mZ�n@�w	�SAf%�ԝ��Y�h���;0�:�4g4�Q)��#;Ђ�1嶈.�;�t�5��3�L���ʼ�Z�ɜ�}�5��?��R��NC'b��������j�'�ҿ�0c0�
���u-)���?�Y�,���Ƌ����9,��G�*%��|�Q��YB�9*p�OUs?W%�16	��A4M�c5�i���έ�����~+��Gp5dGῧ��L2M�n���[��لEdzmq�M��ȼB�5�(7e��c|?��d�8���j*._ ��埁=�Wi����q�Z�Cⰳ.�V�w�-7u�.E7��g�Eo/*�RD�_� d�"z��}�ÓW!�ܧ���բ�[;�D���k��(4{}��I㜿#� W�@W"Q��9Q�)�^H@�#�+[�퉰ڊN[���懑Mb[�A��ڥEAu��~�aw�p�&S�2]�GwfJ����q&Ʌ医Ñ��ɛRb��� �t�f;XJ'Eq�9
�N�Q5��$�	9[�+ -��g�-�Z��9-�����"7�_�uu��&hG��id%�^�,����0��.��8�K#�p�]�Za���9�/˛U� VY_�-�r�{������`���nb۷�-dW�5w�L�F����ʆV]�0c��y)���H�C�+��W�wθl��ho�rĔ4��Q�2Sx���7���"
��	�"���Rۉ�!�@0�߇EP�E�3�M��H����7�sw�B��1eg�3����WD<,2�6^�L���R��	䟳A���"[��1n��n��S�m��զPo���N�)�)g�]�FGT=,�H1�:���BG��F�4eE���]3Ԍ7 �؄��qÀ��Ug�@���z���\aO�`+i�i*��le=w��� 0�-���.��l&O������;Qܦ��t�~ԁ�>�����х��_��	�ܠf�t�_ת;R*eG;G(�PW�e��xw�vnY�&��ct��WCl�2��7nB��i��7�A�h`�2W �D���t͵��4�8�h5����)J���<v+|��`^0�k���c��G�vy<Q�o���8�?�>i�l4o�wNT��,�,�Mc��Ia�Q�A��%�������H��X�Mwټ�O��r���u#4����vJ$��u1���o�$��|�h�\�D�Pn��Ȥ�-��E'�bu�2H��}�O2N4:%��}�D�H�����99*�z�����}�v�)d�i��k�Y�*�H���'��9_��½kx�E�WE�-�����ܘ)təݪ��t��Y��|��.]�B<J�����:�<!Nyo'ײ�]�Q��ч����5�����)�J$����z����s�w��+�1k�NW[��q���b��"��	4%��䤒d>@\����g���7奚��Шh�~>t���twΨPQ�QH�L_�q�3�����[	"�hl�-;nTΩ��{��n�t5�����V���a�;#�a�V	� ��hJr��䘒�J�e�)��sP{*�F����ד��_cڡ]��8cA�Iw*ӵ�aS4����0J䥒- ������]�eY�02��ۨP�d}��`���<>H�� ��^Q��k=�Wk��W������,�>��I�<�8�p#�'�I���cA7s͛�am��X�:ht9*.�4J7�d:�W,�� ��5�[!8�.}�
�WD�jҕɱ�!�؋R��u��<���n��,4<+5t4�:ğĻ��<K�?&z�>pE��ߞ�_� YJ��i/#��9>D�8t�)�U�+;�����_�]��X�0(K=��S���P��֠i�� ���.�[l�w�5��ŀJ������d�m ��A��2c��.j@���T��t�v)��_,1��`R�bj�2N��G�eEY?D{Zb�!~�mq��IOht����>z6�S�'U���,��٬�����C�O���a�ޡDX��=أ�Q���O.� 't5&5�n�
%_��P�sO�g� ���2��#���ɚ�Go:<E���\]��+�,7A`P�}�t�M��-��D�ι�s�����C�����%�"@.�g�;,}U�XAE�7�<�y���c
`5S�@��7�j(�.h�|�_xp0��=�#�����em���('q�M~�[X�gC=pb�8����^�&O�����˾���̸uJ�	X̡]=�6Dc�0���Q��#�"49��Xr2]UE�^���v�u�I	���eD�E�hרUXp���Dq��>$���T�XK��p�
�e��҂@Y�Dx�uDAC��
��v��&�#ٔy @ceqgPg=�d�T-(�	Q�͡�mk�H���x�_fc
y��F��6wܵ�Dl��}�0�pg�t�_����s���_=3�r`�'���(�H�� Y��T�x�e��X;\ԿP��
J�B�靲����8��)k��,�al�##U�m��v�(���Q�"���p@��`R�g.BG.*
����S��t��<���c��r���l��R���D��ʀ�N��0e����	[�:��ɝ���)oiP���ʇw�Q�1��h���E'�p�E����p "��,;p�X	jEu9�3��3n՟V�x5�:Ӭqu��ώ��'_�my��Iǳu}̳K������ p���x�YE�R�#ԣ����]R����}��#��)88=��s�4|�W�-�����[��P>�&��~nxzБ�U��E�Ak�S�ZJMFe�>)~�1�zq
��1��B�_���m���&�VL��- eBD�j9�oa��'g=��ߩa����K�b7�z����l5D�-��4xO���_� �fF�$�q�y����Nn~<�����ƾ�of�Mg�]-	��#���o�T��,��!�G����pw�0h]k+i��ġ�FW��M��֔�Em;s�k`P�t��)���ED�ոs�裄��<�W���2M�6+q`�eq_�q���7�fà
��C% L�w�����q���p���S��}V%
--Q�2���DFb�X�����n��ۼpƷ�U�Q����P���/���`xF�l��_u��%�]э���ii������K;X�P��_>År��m����;Z��ܓ&�� Uչ���5�ݞ�
.���Y������e�DMO�\��,QRL8�E(����D-+ޖ�����2X#��,O�,��;��_O2�}M2!�|o�~<�hu
�5��%���%cl����h���Έ�ßy��u�p�A�|�[�W?WJ�z$���z�ۮ'�a% �x��^����f��?��W��l�Ƙ��	��̃��ͧ�� ^j��5%L���Ӌ��dd�97��IǱ��IJ�t6A,�q�懳�u6����c��5��qb0�=���3E�C��Ų��9�gd�K���|]a?նOw1C�9�!�ɭgJE�iD�(H�ĔD�"S � <�qqpl���8p1�\�u�pS��
��R&O��E�"����n�J1�t��?@ N�䟯VO���+v+��r}�T�C�(Pf��Ͽ�!f�y�<K��*Ix	���w�q�1�X	xi�#�
��U����
��K�n�@�!Nu{��S�����bG�[��Ub�;��7W�פ.r�c耵��fe:d=�*�I����R�_$�ղ�&Uǣ�,F�Q_������f��5��gC����?w{����%�Es����?�yϙ��nK��}���� �7����0`������(�zd=������׫5���,��y9r�.�C�sؕ*OQ�Ah�����g>�/�!/Y�6���н���l\
���]�m��A�m��h��G$�)H��V�smwU�`F���Jg�#�g�F|Z�㥔��ʮլ{���;9
H|wb�&\�u3u�G��nW�����E�����5�^?S�Y��@��x��-΢����*(�ԿE ��dn��=O"]/hO�ZOئ9Xo�\G ޟg�Aa�}��o������'+��z��;�=�Z��Gl�/�}cq��������C��AI��z2����� Y��s�JjaQc���H���1�_y���4�,h�;���-I?��C+�z:cF�b�3
�[=6µ�P�"I��4jWp���7ftn%�*�j�}�yH�$ݕ3�ϝz� [�<:�ő��8e�-lr6�xKB�p�:�o�U��w���9��-׀t��Q���������֙�5�N�l;\}���u&�oLn���5��з9�s��������Bt�>��w�}~ۛ���Q�3vW��
н�)�Yآrj�r(\�|���ZWzzg=���p�c�m7�'>��&�ͲV� ���g��jZ��z�����s>&\N���G���������B�g����Zx��U���?E�p~�s��%s�������iBs�6�@	zKs���iH�Sm2#ʍ�����b��b�o"j;�v���3�>�7�~�2L�Wo�%�8cK����>�/ Z������Xb%;r-u?������즡�vF�JMc�c���S�������3�@�ާ���d9�5���I1#� �j�|iU���[WrIz�����ǝa�v��>��Q@�E�s�_s�$!�^Н[�4tT��~͎σ!˷���4q�+"l:Ə�G�rĽ����Gs���,��0�Q��
�'.��w�/����!��J|]�G��m����ɞ)��m���u�A���,`_g[�y�:Ƨs���>��v�ao�7���J�{5�f��/P�o4Q�nP.�� ��E� ���!�pI�yc���;��f׾��t7�=V��
� .�&;ˮ��< T���� ���+�-7���HPr=vl�<=w��y��AH�D��ȏ�j�{��{!��t���_���[b����@�qĩP��+f�z,��$\�[��蚒�|���9�?�K�ү�� |@(�B�le���6Y(��ײ-�<>��hr���PI � ����s����]�Rj
�r,�E8 �mߧs��F����}ՙ�9�)����n�l}����X�'�C�e�D⌇��[��gC�H7,��=���BN%z	�)=k�|5��4	���|k�P"4S�'b3͙��xC�'d|��)"�!;��m���9�*��΅:��Ք�&2�
<0B"f�f��mRv�iF	׮�����_/�/�Y�!���Py�o�
�2kI͚���Ph���(,	:�z� �h����5��qh]��t�^1�]��W�\��QtN������y>CӐ���)ޢ�3��z�,k���L�!jN���F�q�ҙ+�K�B��������7#�apw�5�+hC����$I�v ��F�\;�K<Geڎ�H��c[��5�j�0���)��j���K�%��ݩ1^lk�W�xi�����Dj'��ܓ�e��:�mr[lo�n(�ڇ޳r/>I�����x��%g�顢}�s5����)qߢ�@�/*����3���'����|�_i�Fs��;-�+V7^з���k��˰�/�(L=K[��]�&R�^�T���P\����`g���NU4�&��R��yϩ,thp�<��M|e>4��?�q��x�ȍ������+K2i�LgF�C���q�
z$X�Ps��&�L9�ݏ�3��g�еNv�����v:k�Y|)�-�M��=˫�*נ�*�9�Ḛ��m�JŋJ�6E��<�n�G't�7�=�w`��=��l�G�u�G���iy<���j��Uj�	���O͛��0����߮�?��&�FZ�G�P�?Ū�L~��^���������O0#�ljGy��xj�����R��"�e����L�*���	�Vd9=�`�a|~{'oԨa�W;������ٮy�+	�p9;f�0p�Ήk�
�'>)I���ٮ(�NhJ���/	J�c�ϰ�D�|D��!�|� @^��J#E[�+ozVHQ%+A��_���C�-��>��������+�K�>��nJ����i�g$��z߉rM%���W����2��eĿ�7z=H�p����
�!�7��>"�I��/���`����Z�&��0*�B��׿���a@�=��V�?$ǳ������բ�j�Rm}c��3ѷ��sys?��U�ϒ��£���]7Dh�UaXHl�.�/j<*K���t�� #X]�W����`B褷r*�L��)�V���V!��qujH񠋼Zb�cAm�78ȓ�Q}�th}� �724����!����NP��JɤB��i�oYh\6�e)����Y�h���RJ�� j+�*w7B����;ڝ�2h�3Y�=Ԇ�ݧv���^���B��<G� ��Ʒ�f�6�^o=�����J�4m{��6�~w`� ]y����r�	0رDl�L�6�z5Y�s���k��Y�?e�/9��)�5~��!��}�j�o1F\�
��x�����(��P�e8v�⒋����#��w�Ǒ�d��Ia���a�W��B��s����@��8�л#U@�I�Mo�� �$����Ɯ�6�auێ���Gi��E-���>݅�V�~���<�A����"Y��
"�������ϣЯ�� x��̃5��]�=�R���[5���u�9�09�`�~i�V��D����G�J�KũUjI=c�c�OKSc҆�����S>,�R�8��ob�p�o����E��}P/Ww�俞�,��dc_.��L:�S�OJ�>���<Ā%�`�x�n��#�)�.��U���Wh��9�&vy��U�w}-5��/��ᱨ?��;�Q��љ_-M���ڤ�b���Ǘ�%E9�]GhH����CZ[kT/{ͱ����`_~M^|a���$�X��IwVb\�cѤ��' d�vu���ۄ!O$=eM���U�
*���2Ӿ���*��!���z�T��I�)T`Wi�LE�׵�oa�?��v4�Nuܱ��^�Z�?UM���SZ8���:���rX*-Z9cm�C8M��*J
}6P�7�FG��c˘z��.�?M��5�Wʽ�h#���"�)���#����#���"���¥W����p����w�jՇ�=uIBee���p�}�:���v�Ee�׺q���k��aH�2����>p��\�$���?^�Ū������&�m�a,а\�n��v�$���3���N{�Y����z�K�=�Åz������Ub���UN�	�jaijl��z�C�����<�������.�}R[���(̎���˾��&5��K�B�gqhU�[*�ۛ�B>]J��m\F�>?�q�ZJ�������hک�u��+@�΃{qK�g�̣���.��Eni6D?&�1\���_I�A�piyB���h���=L���(�!r>�7~�:Y��c�W,ltH*�pBE]h�A	B�K���TmH�ua�˶�(/�*xVl�z @���_�����4�6��=׼afI�峛;�H��Z�A+A⦭F��+�$Ek���m��,�M��Ø�E�>����\��kOxJ5X�C��܇D H��Cn&i��>�����IH`�����Z��`%up���7�`Xi6qd��z����E��߹���_D�Y$@W�P?=�@��-V������x����i�]�7��CT�`NL���o�(F���3=DW�#*!�ƀ�1Æ䜷g:hI����N��<�&p��s���J�-��z���s�?���3>[��2�Jg�������\>mE��Z�86^��ϋrn�Q���?�;��d���s��&���\b�.�J����4�p��a���QxF�ۻ�c8�4ug}#��"h�Np��B/��ܽS'(1�Ƙk�*?3�e��-Ӏ�S�?3ֿ���at+��CP�$~#~i�"˷�a7h荑3f��d����jm����X���4�F� �$�9�=v�t8���rO��&:��U��3��������?����c���7_�%n�K�Ta;�V�}�e8��r�)Oi����	��Cƌ��	7�M<70�q���r�N{2WH�`� �x^�:��h@85����E���|A_p4��l�F��ފ�InY�Z-[�`*�V]�$3粍d��UL�Vd�����h�g]����W�+ksw�
�/a�V��i-����LG)	N��|�>2��㖬�E#y����Y�����w�ݶi��%�SB�$W<�@�X)8Q)��7��K��@����*Ɇŀ�B����ڑv�s��gh�j�r�Ch�5�?o��<��޿�k��ES!oh����E8��o��g��4���e)�n�i��$�-���t�Z�3�W��R���%�g!"s����s"8N���]�ܘ��@4��5b�B�-��)���'_��/ ���]��� S�����c������	@Z�.�|�s�$E�dUO �i=b�x�:�q[�ēq�|9#�O�P�D��&�P��5��ܵT�NR��`���i�g��
__ߜRI�Q��{�1o�n �n��6'p� E.&T��Q�>�h�������p�ڐZ�N^ٙ�++5M0�7���aa/Q�ut��i:�'�)����J�"�K�������7��A��}����{�ۥ:�'{p��cE�`c�wN`�h����&:����s~ �|O+��J��P˲��c��^���F>f��<����y�;�!�4�)2g�Z.�o�i�<��e��^�Nr��#�>�����	I�c#�'��zb�+���)����4���X8�bܰ�+�J�I�j���
Ea��]Ca�t%�����p������'��:����d�vZZ��4�,|��.�\�û"R�*��ޅ��ֿ��D갺^&�Xm~��sq[*�	�R�q�^y�EOKĬ�B)��*�w��[9�J��Q�q����Be���j���R���;��tQ���m�BG�|�1�����F&L[�n՜@��*�ī��}�Yq�q�9{��� ܺ�����a6��Dn7O�q��ɈK�l��j�pYG�KE��:��tF�p�,�iAAB��V+�_�uܺ��s3u��[��L�}IiF��c,�>��`�	�<���|G�r\s� ��ĺM�t��M]���B>^�SJ5}��s#X�X����Y8N��MHş���"9(gVc�����ǳ����\��f��	3��K�7�/��u�K9��ɍ:R��a��!p���ޙi�0�6�|fξ���ſ�,.���p/��%����d8S䷛P����)�5���1���z���5�Q�L�$o�
_������'�[���]T� ���^%�阮ِn=��\:��@�*z��	Dʗ�1�r�4�0 ��q��:�����RK����N��J�@���s7�S���˨g�����7vEG�2�2���&��&�ܫ<%[T�r6�����n �Uڠ
F��w��V��~P�T#Q�+$zSӢ)G։�%�;��dA]�h^�.�$�\�f�ں��|������gb9���%4��5^�X����ɳ�R�j�������ծw^F׻���
:�k��3��0���I6qs[�3��Z =����7�\�+�c����n���ຆ(w���b������g3������,�^˾�=!��ת��0� :�%�w��fx�[���m��H�j��)�Tx=Î=��l���FJ&�-�:W/e\;�����4�۲���
����|�ږ��$�^�ah�X@��R��vG�����c�rt����t@)�&c�ĿD: <��;�?
Y����m�I=!t̻�?=Њ�<� /��6szڈ�a�{�	Ļ��F�Y����4���|lx��)n
V	s2$�@U�:�K��we�?sb���>�ܚJ�ݖ����:�6#���x<�o2a������ի񆫩��)�l �'�3�~jp�������b�hS�b�QV�A��p��O�q=�O�Z{5�g=[��'��w�p5mв�l]��)rDL�E-���}���@N)W*i�B ��<�Q�L����%��>�<�40��p�a&Z�̤J�h䦠=�'`2�Z�7n�J��.Q?43|*�'7��2���0�1:�9�L4Y[=Ш)]f ��h�9�Ra2��zZ��дj�ړ����X�cd�ҋ�@�sQ��	���|���j"$�[�n
�,]���H���+?�:�cs_'�8����[��e�ǘtR��� K�5E�g�L��5OԡG��ۓB�����yD]��*-���!�.`���7��N6l�C�v��t���v�F������7��`����(�%J-S4�"��"�H�TyW��|2&�{X�랙�y؞����po�ÙM]@hTГ��BW[ٮ�K%ʠ,��1�e!�V //�$Vr��u�]:PQ5�f�U��=�;�����M�w�[�0A���+�8�Z0{�Y���^B��ɛg���NHXHx;�>�e�*^,R|��[�����]����?W��ta�y�s�6.��P3�4P���V�MMf Վ'���^�����h�#]�<��JM�U���3�$�?�j��t�%��]N6B��k<`'t���8��e'�R��	�Q�%�7�|��yO�+MS�������+�$	�����yU���8	!׌;Vri����<@@�V�,i�b�_G�U3N|�E����h�PIbQ$��R&�� �wa٨!� &w����!���P����5bRΡ���MS1@>�Y�b`-�O/$0�D��<�'�~ꠗ�J��G���Z�Qu��&2���嵌4͌ԮX|v�g��ż�d ��T��Ar�,�n����J������@J�1�SvF��F�<p����i��$5�dd���#��U1y��ɿ��P}A=ܾ�`=�d/H��p���\p��y�K���H6}x�D�Z�����?�9�����q�&E&Zz��9�*l! �����!�S���5<nӰG7����-��\P��Z���s5R�~
e��3r+K�$�b;GuP���$�ݛ[�<8]�=m-cu�8��N܋��A�U���̇���\�1i�9;y���!�{��xj�h �梨���>�����O�w.2�Yi-T\�ܑ�L�<y��w"�c��
�L��vW�(�q����wj��py=�WF~��
��k^����>���U��)z��VڔX,4�5�'lt�=��&�6�Ή6�/��7ߒ���]�^V�N��M{���Y�Y�v_�b��:X�/�&r��*3?�L�m����a�;.E�ܿ.��5T�fV��l"�Y,AO���.
u)�v���4&���3��4l;�S-py1ʋ��a�{"�g�T�[ʣ~F7`f�J|�$�\n�Q.�z�d�@�ȱN:g���,�%=E ��k�8�b��^���4=�k`ֿ� 2>�}�̢xg4Zi~�j�8(TF�5��p~H��۶��b�d��hI�^�G#{K�WE/��^����e>��&4B�rc�[����^�Ѯ��I���^6'"2t�O w3|ר���L��Dm��n�)8�`�������tr=효���ch�G��+���v�� Wu��:U���=<s�����(
��X���mƜ�͖P�W���xx17��"�����ԓ:&�$H�TD�T��_� ���ĂC������|����t�p��%щ%Z��U/����D3�	���1��%��(�0�,y�T9��&n���(���tn���������|�3~������T1���ɕ����f���H��g_�zҕ@�����޻t�EZ��ؙ(��P�%5H�95֦�Ngnym�̭�#�ئj�c�OS&�'82��[��w[���8�f0	ˑ�q2��,gG��K��Ǡj>��(BA���{S����Fz�]�U��>�J"�wx��A4���p�Yu�����Y���F���BZ0�bW�)s�Fjn
^��H��#}L��D�F��C���̏8#4���� tԡT�������V=��"k�U<K��]��x��lb����7b�jp�!F���W>X�l�-+��va�����/ ,��Qc\:���M['t��_��YѢ��C6{��J=��9f�X�rO_>DHi��zU�$��7	�Z�6��6��,[�ml�j��锪�hF�28n�$�2O^~(��%����O��Y!F�6�'��2f,���?3���Ʋ���)*�gBKUu�{h��S���sțn���D�Օ�Z�����6�a�iNzD��X��-�g���&�:�6�snX���D�ܔC�]�3�������1ϲ������K�uSM
�:׶��a�Z��h/B�I�{_غ�g�x��Tv�� d���e{����m���23����'�^Ԫl�TZc��(�K�MsTl(*2>'� ��� dk��\<?�[�Q0}���T�՗�6q�p	�h"0��w��U�xU��WI��&U�����^���A��k`��)��
H,ҫ[�����M����(��&MN�qx�]���7���^x�bԘ�丽�YU���>e�͐}j<�i���
�Ƭef��p�yu��9���xX�_im�t[@C�_A���}�_=K�Vت�#��#���IT�X��4�g��J����ox``1@�ܝS?\涘��5m����'Oq�43��*��^J$%�t&�mʠ���}R4&���K��l��1�V�y \rP�.�m#��7����X�l�H���@�w� ﮀs8�H���e�WUߝӹ)�RǠ�o;,֏2M����N�9�-/��#s��d`�1Ҳp�#��Z��Ld�۵��4�{�_(�Є�C=����/L�  l9�@`Lm���蔑G"�9�������R�F�F�K}���*Z��py�
F����<�>�TxI��K�x��PҘ���v��C5��9��r���WL��%{�t�T	��kF&�ib��PA]�I��Z�t�Q��'`cm�Y�Uƚ@F����i,�#Z_��r;�S75����4��i��F�d*��M��&3��
��i`��;�pL�����tg��6UQ��X#�O��;<�"9�֕�
� Q#�3V; ��h�^{��&�Ti9k���m���J5��}��ܩi^��e��`~5�F�ڒ����N����ԜxN9����Ҍ�>��X�~V��TFE+ޕ� 
Q<vgd�6���V��K!6�WF�����.����k�iGq��[�����
w-�~r�[I���������M��-�ڹ�ߔ=u*Y�ME�o���]B�AGCkc�Og,��@�Ӂ��!�C~��O����r�@l���L��8�v{Fn�te���oc��Mz=g�\�3�~y��<�� ���e��*��Ύdl�ϸz��yN��C�t�hB 
��vT��;w�<q-/v�c���'�G��tq.k�w5�-:xb��!c���y~�g�����͟��[�����OYjy�\����{S
L���HTV��g��*-�����t�2��-S�й�Y�H�*$�����4���b�=���"~c��W�%��}�6�b�`��Oc���'HzP�,Jx�N%{�]^?ZPr`2ce�2Z�t_���b�s�I����9��w�T�qY����6�.��7i�S?�Z��+għ�!�Cq^!'�x��|�|ˉ�fi���\�l;+����#��Jv��V0�G��Xt��m��@\�/�7�������T�kh�3���s?�z�'{�~�$Cѥ���'/�Vq�sI�wET[���}��9]�m(�F��lZBl/`0�ӻķ7Z+i���YpW� ��|��Ye����鍓|Ds9�s�7�K�Z�0z���+"�~�u��r��n,�����4x{1C\�F�飯����#n;�s?��Dn(��=��/�9h	���sjE��:���&����q���I�A<?zp����!��ݛ�L<c�"�����q�5:)��6���)�!��e,6�[��{TS��#�C�턻�����G����ԕ�eHa�U[��^�!�s�*�̥ I���ɉ2��r�y�E���1�Aj�"�I�r�+�olK�+т�����(�/��%��J-�3�Ι6��O�{~���^�7}�򵞍I�vdp�[[(�tJ���bMl�4/]ݨ�h�����1�VM���5�4�G���>�$��M��J�W,&�eo�_.ݧ�v����>[��6�����r�����U)��&����(+��\��M�6t�u�=qh�bLt����=?���$� ��œ�,���2�ë]����3�	I�e����/f��h���U�����X,�)�m����*�h5����9G�=�j�w_ʸj>.?�Y��pdO=M�3��͕�
h�t��B����.��[�������d�	����Itlg|v��7v� �t4
r��(����6���W���[�F���&g�Sa\��	�����8�t=M�6�a�~�nvϫit��D�t��pp�ڑ2���{cl��!�Ǖ��{d^�fIcqK�����"7f�]��Sʓ�r�Iq�;��^x���R�[��Y�%���C������\�� v�iw!�䶪h��$����P�x�Y0�3g9�<�M��[���-#�3"Ao���Rԉ�v�5�Ցk�p6~����wȵ)9��/,YC�{�����Yz=^��i'�O��/<��!<���u6�ͬ�k1`O*����� �%.f_�-�"!����r�=����λ�'�?B�q�����X׶<S���(���21{2dюm����Eٞ��k�%��Q��+�0DZʔ�����:�;���pw�G[�lp(!��e�7�UaG�F�F}:���;�^^L���a[7�b��,1K{x�?�o�� d�"O�~�����T��d���K�2+ͳ�1m$�Oz��DD��v��,vLȄ��Ɲ�8C�Ng��3�ޒ�F��������aFOeq:$�T�ק�� ��t�0c8]�z�ZT�A��T�<d2@i/X�e
�C����Mڭ�(A�_it�
3�˭�o������2x�}��P���Ź�3Y�`{����}M��\��J����)e���Ƴ*�&� PRN�]-k�^`G�_���5U�}K�ͥ,sSv�(��Q��ЕO7�������`K�ò��7lT�&����
#?ߙKOZ�T
?�>��ҙ����Ƿ�q�q���<sd�ץ�������T_����)A�y��0�U�
��Հ�¼Z'�7O�躡�����R�B_~����hī�� =%�W��`��!�EFS�|cΊ#�����2���F4�E�5FQ��Lt��2?�
�n�t1J0�̸A���`�F���yϒ��_�%R�M��V�k,i�pҎ�s5��@�.tce��L���ΰ���9p��L�2�ݺ���ֺ����X��y�6��~�H��6��\kՙ/^�x�ww~���L]i(�y�g>jo=S$�L]�p6WW��\#�|%�'" ���Gz$�-椄��~\������\-��Ʊ
(�;�=��0%3U��蘒6I�Cpk�nt���ܲ����S��~��@Ԁ|d˘Ӎ��?��r1췲�{
^,Ҙ80z�A���a�8+&�N�������������3�,5�_�8�{~�a�����C����:�|��L-��
J ��ʴ�Z�����G��a4��K�����~(��5��z�^J�2���4��2�J�����O��^��pm&���m������d�aK�P§�_oW���Un�Ca� V���Փ��BaCg��z�z�*�.B�Ix�=�YӵÂ?	Nۼ�|�h܌��_/T������(NXI��_]��)PF:Y(�_n���4�˟/�lOg�}�t§��&+���;_�ß�?� %y�s=z-\�T�e�9�)�\��T�}��� t��M�<T.�yð���f���� VI�j��\~�h��ǫ~�4��0|�v}�T�u5W6<��S�M��A��a�������T���l`�I�Q@�.��"� ?c���2E��_Kk�0����pa@�Cb�a*n��j|RϾ�nvV�OJ�b�8p7��h2�hD��e >��+���|p|�p/�䂧��f�XB�e��9C`"�fGګ�j�=7�)�H,�7�/Vq�D}F߱���t�"��/�uؑ��Co	�r��ے���>t�[p��������R�o �#'���^�x� z��溜̟�J�K�5�'ݜ�y�R.����B�@��c�tY������[`ߕ��(b��%��!&7:Dy���T�_�悁#��gz�z���>������p�\s�b���sӯ�R}'�lܹs�e,�źpw�.�5<=�:�N����A������>��t�����������y/jD*�`��nhK/�Qzk�R���'c�V&�����N_":�))�N6�ߋ-���9G7�C��f�Eܐ{I왑�;Uk�mm��qN��2�tײ�ѫ`�wh?i7�:�N�u�`B�o�!���NOm�*Z��6%��5iDTFcs7Fi2�5Y�6XI
���[&Ek�aA{�	�Q�3k�i�-~�&@��c(��Q�c�\�2�Z!�`�7�{౻ʲ��)�n!2u��V:6x�{�b7^��p6�Vψ����¡/#�D��-�� �P�a^@�+l��r��i@�/��܇Әnb&��$��؋g������K��C��7�}4�K�s�c�v�%�P��/}�2-_XŅ���jq"�o��q$nLC��kP�����i]b �� �c��d2eհ�X��ymy|����M��{׼lzK�ښ7�Y?�|��qu�VX��Ǚ��㚗:sML��i�TjJ1؊7����@"�É��mUb��f��Y�;L&\hI�Ť�"Ö��u+bV������m���^b�<ݝ�ڏR<Uh�_}s��L��wT�(X�0���$�����s�_[�M��{}�M����sHZ��U"����_/���#�U�>�ш�#��;�X=v:ﵳ��C��{�zu*�j"�(*_¸�JU1�1mB�P�������!��-�̨�e�D]�OL	0o]c�r�,���$ "O(��f��T��:���,H15�1��r�BJH- ��l��T��w��~OF��\$�dv~�Q.�
^+������XaꞸ����a���X��F&ː׊�{�qBX�:Gv�e��D�1q|B]q���#�o#��u�����W͔F+��T�M�u�2{�o1��T���B�>�>���7��V	58�ν�IA��͠�K����~�/�[�5���<��Wa��~}i:=�	Ï4�b��`I�ȕ��'������M�6�=1*�T��P�]b�ä;�?B>�P�e�S�X��͉^%��_{�>ȏ��`z�=��� �����$���G�*�Q�ɖL���6�L)�v�-o����y2IÃH���)�ݮ�����zLo�V:s*:�4�|��ILnhyHL���؎��|L{r���ޟ'ϧ��C��_C?�U�a��&�ӷ������:4 �H��]3f��m\�@>����[�2�E��4�ed\�F���0`��o܃�O�����,��2��~�Ҷ����f-~�^��	�G�>D�"r
���`z�	 �D���h]����k�"���ͫ|̞Q�-h��?�.y3a�f߾�����Q7Cڢ�<Kӗ`i)|ơ����>a��r�_���\�N#ݒ��!�E� A����@�T�y���4�̭�3*jnR��~) U��ٷ9�H5HP[tAݍ��Ǆonl�t�cesXc��\8�#nwq|��"�j�.��do�&H�$'���@���yv����,-8�x�7e����Ხ���4��"�^�ZR�j��y�|]�zX����`��/�ncv+��L�-�k�>ֻ3���@ �8\�y��n�o�(�33�3db�C�f`�'Z�LÛ���A<���7[ _�T�si��Y��fTN7���#��ek3�r�t
�4��/���W�m�׮�d�Q\�a���zT���{���wW��l-K����L�x���t�h�!��g�4���2�r[	�����T������]�������܏�nګJ$O�oQ��	̢K)�p��\��R}CI|Dg�י��ś\�G_Agg�����Pu���b��E��N;"5��:a��[%g��9j����$�,9
Gk�!��O�����m\�	C:
��N���	E��'�����G��5��|-��p���ނ8��^drBy���Wҿ� ��!�H(<g$�H}��?ذ��0�a&S�3�C����ι��=�8�E�_����&#yǾI���{���
�*
^�[[��Ee�d�i�����{:1�4mxn,:��;{�t���G��F[�di���#�X��i�f�	�kgG����i�,�;��l!�/e7��q�a87!f�����G�}��ځ�I#�v��]$������d|�b0\U�U���b(�+8/8��7����Uen?_�q�hx���K���ñd�Xf��IUc��s��{#p�	�5Q��\��7���+�����r�WcQI������CD7��3hs�kd��&����蘍�(շB�"$�F��7��J-j},�^��Ǥ�[%���q�|��I�Y=�=��8x}�GQ��Y��}�C ��L�@�C�ro~�����U�D>�Ш�H���8ep���t�j�V^ʑ��Gf��D(�~K�{�Jl�A��sS`���F���OS�VcSku�hZ�#%�Áۺk�5��K��.Fk��)�\`/�C�"Q9f���7�U4G�A��E�(5���h����%nK�%?w}:�8�K���"C�$���jH�N��G�����c"�}�,};�Tiώ��XcM2�d�d4��#lgX	Qъ��Ǜ��*��|H"��O2�"4�	{A&X��}�$��L�?1�Vl�:ƿ���P�Z�?���ｳ�e�����L��_�%`,�wh�r�'t�	�G�s5���T��Q��О;p���F����w仐L�G����"ŎI5�$�WPlJ<��!�T{�&�+�,��HM�E8x���/���T�*��@��y5e�N�@�W���OVX(2=Ik�?N3b�8�M$�����Nx�Z�q/���T��7@��I��Lj��e�6]�,�����B��J�dꁷ�`�ԛ��2��G������ $�d�����I:�	�u�`�a���Z����ˋL�l�Q����뚱��A)�;ð.�ٿ5J�p,��L=f��
��-��\��U�lѫ-pbb��Ho#k"b�j
"����8G����i(;����d�vW#4���ׇ0s �F]����Kʾ�&�A��q)�}z������3�[���(<1 ��ʇ�i"U�HY�y�=�13ߩY]L|b��)��Q*~��čy���ݤ���H ���@4�N�.�g�g���V�}�q��n=:Կ��_}�z��n:�5�j�L_�m]刪��(�5"	�g�����W�f���F�N�ҹ!��P��7�<�S��,�9K�����H���gj�3�T����&� ���Q65Jق/�Bq|Gx�G2"�m=�j" �������%)��ix�1[ֺ�"��n>W�x���u��x_��D՗�1���AsQ/����_�P~ϳ0� t,7Jx �α�}�q:�cp��9��ц"���a	����рs�2 �H����%��?����L�?�^cD��f�~%_!w���L�M�"I���՟2=0�gS����i�_xK3h��Fv�Uz����J�fS+,b�u�3�6����ݼ�e��"�b�C'�����p���h�ݏg�K5��8���G�%�g� AJ$.'�!G��[Y����s���L7nVHD��-�	����$G{���Mժ���o~�՛� �2Q`����na��95}��z���IY�Y�	x0��cx�K�a�9�k����o94��x�f3����۹hW���r����߆Et '��ƾ���R�Y[	�tx�1\;[�ӡ@�$�n�o�;E�y�ZƳ��8Ҭ�1,UE	&�}�S���׌7�p X�,v#{h��13 mAK,�-�Y&`FCd�C�ᒅ}�3rIC��R�ŷĥ�Ch!q�+�"�˯~Y/�Ѱ�o��o�,�(��_�7rz�4|��oe�;�� ���ٛǙR��~陵��ΒsO�eQ�M�܅��d�3��+�gQ�ܙ�Y'{W���[橇b�H�����kB�ӭ|���(�*qς�Ƅ�ڞ����"<aU*`�Ӗ�ί�^Js�yqHfH�@6�4H�4�`������y�D�.}�V�j�^��L��RSQ��|�l�H:���g�㏔)��@������k�CFS��y�eV�bj|>�O�
+�B�*�?\�
��鎼x��8L�g���g
�&"��좌J�/��6���$73O�����1���e��t��ϔ��9��ۗz�-%��ڟVN���m�MN�5,х�F؀����&�
x�Ef>v�D�n�ڇ��խ�������p�Ӆ��IaG�f��ZE�?8���R5@�*�~F�(���8gU�_J���5���ғ�x�& Ӓ����>� G�C�M�շ����S���i�<<7F~�17xtZ(��t&�a�i�ǝd�L�mmvL�V,I�)o�#h\MP�K^��ɨ������+L���c�Ui���^#,�Z�X\���[��$;�D��t�o�$��u��u�ە�4C"i[��ti�����G}�����Kg'�Iv~i�ݯhҁ�lU�n���Ζ�,K����<��E�N�~����r�G=Z��,9j+��.T�Ο�x��Yc�qw�����%?�Թ-X�<���m"���aۿg�l�i,9����q{g��p��p��.{�* �Xx�ܢ��(z�}��O\<g$�^ �l���?�f����Lxq9�;1�z�Mo(�̰�3zԁ��vx�h�ئ��L6��1��CߎԸ���,c# 4�����2���e0Xx0<�C,��ћ�U�mq^K �M�_�Z�h'�Uy�2f�G���@��`L��ur������J�[��N}vq䩝�3�"]ё8���j���� ��c�e�Y˥O��s=>y�ȖT��nd3��X�4����5i&Zf�,��)���oa�P �03@O],Q�v�\�Ch��"VV��i�n�S_�C	�N#ٱv��,+U���)��:�7k6q�U:S��[h��?S�#����]�@+����SAnw�����C�lN��Ǹb"61"�x�Cd�)8:ES���������Oa��%��KtRX-y�1^p����H�ׯ7+<i�o����]ݳ\bk�9 ��!���C~��.!!�~���"��9�>��f��W{oh2L���ƚ�kKwhɜpɬ�$IU�%B�p�{@��+�ejb#�r��U�����)�U�O0��Y�f"ܩ�D':π�L�DP�+9LY(�+b���%��1iU��)��~�&��к�� ����H
�>Ỡ�W�4�|VZD'��TJӪ䓡"��Gm����qGS@�&Ձ��6����H�`�8JN�MU��6��#�u�ƞEp�ha�M��i�vE��dPs����	|Y���*���k�Qܱ�\�ݬBF�ϼ�7$�։��P���i�FӦ	�f)9�j��d����-�w���P���H��=����o���<#>J7x�@zʴk�]�'b��p�m�Af1���~z1��s�Ŵ�〇��[4�����1 �a�s;J��C"�� �����S���-Q�z�؄Ou�K%�B�P��u���m��̟�]^ϸ#
p�dͺ1X��<T:����hc��A��*~y��"��-�Xw�3N)U;b����`��T2��������n1T�)R1+Ee+�����(�����y��lI�#��޸y��e~���ҞK`/��b9 XND�A���b�<';~����$������v�`
��.�����dS�c�G0qM"?׀N;w�u��dat)=9��j��`��䓖wh�ѹF�������ll�=&���躧����9D���"�M�7�L�N�f�[=�D$ �{(u5� �z*��s���2���FB¿Ɗ�h�h��mM��+���Z��� oc[�"V�1��;t���`��9���#��h�^�i.�Lb:�"�jN���n�e�եM��"��{�QH�BP+�������B��u&'���-N@ڷ2��zD ���Qj���z/.Y�ChL�p� �����=�9x��.Y14Vv�5pі�ysU}�	��<G*J��!���~1���e����]�W.I��1��诒^�@XT�E]u�4�3�\P:�Z҇�G�`�1P���O���py�����c��Ueߒ���}�
;�2Pz�"�"SՖU#����K����2����>��7>P�E������̕��\�,{qo�����1��娜���E����K�t��}(\_��jJ��*��)5t�&JD���ɣJ0c����I����P�C��l�gÉ/�Q0�7 ��
U�����7��z}�4R�Xe�i/���;3s&�d���L���1��0�
RE*1h�cH�R�=h�dؼ=$��`y�=��6؆ٳP�C���F�M������w���?0�9�=��̶��~�5��+?I�2��o�fR�BNv��3��s� �C0{�,�G�٨L�Y�.C)8�Po�_|�����1����Z�I��]K��<�p���'� �����͓RW.2�e������VB�y��d�)u�Y�̈l=��c��@D���T(}� )'�j,�6e;�����:��w�l��jT��d�WwێZV9;����6'��im�h���]Ʉ<��d�O/�C4��3�NLr`|�vWx���P@����Ul�d�@":�@>p+�Y��ó9n�N(��{O�K��%��]��	A�,p��sA��Kn��Ӱ�~�̗���ZAG �?1dPp�H<.����4V�+.��]�c��=,�8)�əQ�Mm��+�s����e�J�$s�?�m�Gzw)�1m�� ���*�)щ��<5����2��[� �v��L-
F)�y����sx�����'ƚ;�8�t���g��t�h��������WV�g�.m�2���K<�M��H�>@iq���@���9�+�o�^�$Ot���lxq�t@j��$Խ��"�xՀT^��7�F���9�c��'�"����2�e�\Gg�ڧ,���>�t&�R��L:mo9�٧p��=*9��ff��Jy��8q�c�N2>���ύfIt��2���0 �MaK�6����g{\�ve�T�⢴���~���X�-�0A�Lg�m����u�� �W�Uo�&P�=x| ��(�o��J��k(��4!��yL�	�����A��x�k�!v�mb]c�^;�9�~�I3�r���a�I%��7��������Q.P�O�� C~��һ �ڊdT��˒*P�|��ɵ��	r���	�bL�i�n�z)!6jd$'�=4�=0dER����H1d{�I���*W�vRc0|0�p��2�sފx�7�Lo%Jo�V?5�VL�W hv�ju��G�.E�0��Ҙ[B6��K|�E~9��,��lQ>���B�j�J�~)�7��鸚#�*	A��f$�ol���;���#��'�P�nӁʘS�ȼ�����`tL�;RԠ�z<&t�:���%�g��n�8nv�r) =sFу)�ԛ���_��u���=Waxb���@5���m�9#R6�ݢ�NŮ0�f����T�_�3��O ۀY�k�����%�>�	�Dj�p��%FP��<5#J3K!�v�bl�$�\�!9�.|���Tp�����?`��B2Ƙ'Y�AX�VߓC)e�7K��'xV��su������t,K0Oe��}"L��^4^��oK����y�#��.�	�v_E�4f�u8�q,�����;C�����0�IɃ�8=����xսw���ܴ{�0�q}�"��2�͹��>�	�a��Z��QߥQ�[0$T�d��F��OJUu~ː��=���%��<�c�y%R����f��%��C,�,���ٳ���(�\znJCi��n��uO~�Zs�8}8�z�Y�@X��4��0ٽ8�&��Y���-~��B��"���3�əK��74���q �$�q�`N�Q` }INˡ��\�ʅ�D���=y�A�Q��h�?�������$x�b�o����[V˝�k� �%��#K;q�~�̱f~ ܜ�\$���^�&r����9��$2��Ș�RtA��&��Xy(����)�f�5Р�4�������S�C�������(;���c|��'�4zV
������hW
��.�ˠ����P&�א)p��OrE�� L_(���`.��� "���O��\���M�� V'X���yhI`}X�u�<����?)g|���<��
X]y[�;��ڨa�Z5.�ޮ�RԿ.���Jb�[m��4괭oy�c<���c����+�(��ĕ�9�ΙL���S㻀P��~�(�BO��ɴ�*kH,����zF׵nn����V����iӧ��7�xU��sp�GhH��vC����!dJq��=�w˞�d�4��7��5�%��r������[�L��A�l �<��puH��u�E5��-�"F�	\ǩlF0�+Q�zh���v�qm˩��ZC���s�G���3v	o�*n�h��ի%D�hmZ���KY�$$����%�Y�w4�M���E��U��5`��2<�NA>����	�/�5�oL��l�h���䡁���-}[�r�+��M��������F�L�*w�Q�����
Cq_�o�-�иu7�^�s4���������D�����
�_�P��ʍ4 X�M㘊hW�:�ϩ��3Y}�P=	hHԜjt�l���.۸3���T������Y���򞰓��@�(o �'*Ĩ8"���v�a��X|�6�5�t������Ϻ]���Y�gq��w��zyZ�r��L)��WS�@Ǔ�AD�*�@8�����Jb��[�6�[ 4��dUt"3��݁aß�v��_�����D�ن��mC$�U���E׺y�8�t�����F\O+�Z~ep��p�EO�k����v=�Zl��D��|C�+��̵��L��������n�V����~���"�Lm��(v��7C�Eτ��V~ܹ�%�3���]*���Y'�j�����1BNJɞ`�U�GC�T�UȃZK�z�����RB���*�5�L��.�o]rݓrn�Xǖ�o���Ο�^y�Hs�Nλ���P�X��g��2��'6����Q�Y�1ؘ������!t�o�����M���{^�V�&Į�oSj�)�E���ˀD�Z��a!*�{F#
{����}h�s	��$n�l�Hߪ7/�&4]��D9�<N>/f���[S������{;�>>�'���*�fz����V�wtR)z�P!K�I	�FnT�c\����z�<�����v�)�����ҏ�(��N����P���PR[ea!�|ʕq]
B�Y�k��Hwja�~dz�@
��\��P1�|�6Ò��r,�m⟙�|Ѥ�4�q�����w\����Rqi�A�GeX�FYw�N2�Y���t�Z�;]�7��:�Q!e�(� t|�+��K73Ӣu�ݽu�Rq��y���P�v>�^W"P��;,�rY`�#��"��䛟VP�ZCH��B�� }Q�ằ��zvX-���'��O���_���-N�2DW��y��yl� Kå>�XFsP)�c��`Tى.�
,ls�Ÿ&/�t�.��usL @��>y����:�*]|��ڃ�N}a|����:�Fw�͝oE)��Ԗ��Oay���U>i�><@諨oP3PT�O*m�x��6Q�-A�:W�3�S����K��R^m�Ҫ� �	��xm'�3�����R�Ȥ*"���7��6k=��;�����$�4�m�fd3o�F�Y��,jL�p���V�3��'Ltq�|7�D���}	kcD�S�9�Բ�&L=#X:�&G�/�.ڂ"�3�㑻��J!�m�<+��n��<�#���G?�D,�a1�#1j��Y���ۗ}�w������{�H�����0�`��9_!g?��X����4.`M��9Z6��L}|��L�.���*��o��t~��OQ��� ����G�@�`d~���1A�iO��'��T��=@�#����4�t�b�=i�<��|�[�.s{����.O��_d��� �,��#��ic�����? 5u`>T'l���Ҷ@]~�,�151�x�L����X�p�W㌌;r�{y����_F�sͽ�QZHW��PC�캴O��a+��#�d��dN�'!�ʹe6�
<1���6��|�[�,����2�D�0K?��rs=��\�����q�^�@�I������<']hN���Qob����!�`�&�⩑;�m���L�i'� \�7�$]'FG�r���X�L2�$n����r�Ս<hwb�8��_��$N�Bt`������s��LI���O�
�»�T�YI��D���h�r�b�oo����3��`�a�4i(V�`���?#��y�*kZ��C�4�)}�,K9��%FY���|�e Y����𖡪k�8N���ꍠ(b+�ٺ7��hbe�Q��j�s��58"��B�wj{ꑅ�F��Qf����1f�8��(���]��L��aVi��ʖ�<���{G���`ٹ����=�F�A�|L6g�iY����v����!IBl2��������1�������vre(�� �߻`W�e�@�m��4��`�S$����"�H�(Z+��Ԑ�Oڇ>=�sWXg}�A���fپ[��B���d�E�؋g�c��}�g ���d4a�~r��u��{��}�����hd����ꯋ�*:=;)-��k�T����[�Cdf�ٔ>�i6��Z%-)���U~���5%/�)𒉣�
��e��!�b~�!�芭����+
y��=�X��xs�d�t����X����7��]A���2�soZ�n�[�K(��	�㏭Sw�uQ�Ã����aj ��T��5e�2�'5��)>И��`�R��j�D��芎,`f���F�(��$d��B���{fk'8AS�!G�eg�/btG`��x�����=?�4I�.1̸h�T��.�~d��Kͮ��L���3�Z4p�I[(�ͩ�I@%v�� .>��e��F�2w�wj�#�WݸE�2]}6h�����_;%R6�Ÿ����i�H}��c1�Ǎ��|�U%��kX�����Ja>u��C,.�Ǘn�����Z��u�'�5�� ��T:����Ysz[x;������o���6@w��J�~G�V��%�k	T|9�pg�!��81jU��-�l#�cd@�"��|4M`0E�����|��
��~g9�������+��3�tK��L�l�Px��d��g0�J��h��#�;�~�+����4M����H��� �J�a��#��֑�����s�.��.�zO�����z�]�gͥ�pd_]�"N0���0��ب�U����[��'�etn�G���<z����u��t=V�f�9ۨ�r;�{X{Pc\�ډ�x�&1F�2��w�6^��ˡC34\��
1-b���rɖ���q��#��Y���h
:�t��/
�|B \uv�J3�T[�	�/@ z�ą7��zV��_:���EB�|P�BB���铳�B%��$���4#��D+��2����3�TW�<�����;��f|�g���aA�֖��F[� �$�o��Gy���P�����"��Ϸ#���ŝC]��򢸠�uӁ�`��@PV*�o�r��'�������8���(�P<j��M��8Z����d��:?�%��V� �@Iр�Z���l�h2�O����=e��	+�jf��|�����Q�����,���:�֜d���OS�S�8���R��J&g�Sڌ��޻QV�p�l��F�%dK�d��`�.8`d�b�"��%�648���n�m�`��B�oV��7��,�1+��x�n�o�Jh_`>��n9ϼ��0����l)��4wɊ�3ɰ:�؂v<�Oǔ){�6��o8�r<�.J�:�粇��݋��t�f2Ʉ�A�L����{�E&�-�G��<p����t���-{�]�g�
����wi��(�,�b���%��Y?K���v`��lm��%�s`�g��X/��Wj�:�<�B�l��nfV�/P�-l��%'�u�.F���0��� N;6K��8Bo]q��\���353�r�6�r�3<����+a����Zz{�� �����L�zzaL	X�� 1�,5��� �A�V�_OKgr���ٺ�{����8���>���n.?l��72J/[����f{�t�vh� �[����I�ͳ�:~�����q2#�I�Eu�����`�	��N3W:;±����(;$Lu�`穀>
��jf3�O�R=�����`���E4��YZ��:�=��SYeq�6�Y��a&#��Iz|�+;��Ы�.[&(�%GJ�O)�5�U<y.MS����\�=���ќ"e�۪oȟ��d���>�;����y�tt�^Zp0�����ԋ�꾑��"��k�D;�9aF���g��
��?E���)�t�Xm�.����0�l�^��01��:�;1��!|�۫�6S���6�c��2��I1�������ڿ|r\M�Be�<Z����P��W|�0���6Jy�Z���;������ϊ��W�{ko�5��E�b��OKh��LCM�N	&�����F�}/mE�����H��)�zL(�W#-Կ�������h5��"m�}1ft &���j:I�DjQu!������B�d�Vu���&�Goы->sܳ"J�b3%T^@�G�W)a_��m�8z��~�ڱp���R�(�Q�����[2�H��r�;o��Ls���o�_����������6��	��&C�$��ս����>�����0�H*eV�c�$�]���7*����#���~�L?���E��F��r8>�F����]>M�x��b�##�5+�X��@rc�e���0��o$r4����0#l�K��_��ګ���Qϝ3ل��kz#c�t �$̀����S�7 w���zc�\��Ư��M^���������ZD�郛.���G+���D�i�IC���r����k�Me$�����V��_��B� ����%=�k��,ʉ�'�Q"V�:�^��h8��e��E��|V�</ެ?�Dym޺��#���V�3M�A�uoP��W��)���L^Cq�[��z�p5�O��5�C�W�S��E4l[�uQ�Ϯx�?��JM��
A�NN�V>w�X' ��
p��r_���MJ{z��	�sb�/�"7����9��҃l2�b�X�6���.,�23�,L�C�I�{r�����ޤ�����!���Trcn�yW�rV���v&RsԨ6�+�k�=�~.�\�����(gL��&��#��ƍ4u���ɕj����%�X"7������>���ʦ
�63
�]�j(t2C�i�rHw��c����9�Q��� _b>�ہ&�W�騭�h��@�#��{����f�a5�%E���2g���S�taY���DՐ���|��K�u��#qD��V5"v�ll�����"ۛhr�����Uǹ�f��;q�P�����T�b���}��am��S?D"[�9�=�$�g`J�8&a���½%6�]W��d$�h^���\J��7�i�����у�g)@��=��s�;��'g՘��D��4�xc+� �Z;|���Щ�A�SB}e��=es��\����-˸Lh�y�ظ����-;53;�Ӑ�x�YwAB��VF�A�A߭��<HI���D�9��5�Z`��y��F�sQ�C���5�����&�:�S���z$�|������jv��Tz�U�:��t��2ͩO}���� �G��y���'��`�ڹ��bХ�卤�f����,UG)Z��~S|7�z�n��]��t��ϼ��Hw�{ڞ�I�Ʈ�^���B���H�������+dx�\�
�{)/K�.Ѝ#����!1�sIP� �T8gv�i;5g���)��Ȱ�'����ʫ�}�.J��M[P�r����|��(��#���l��]+�T�L���t��s!>.�ɥ�[Z`��F��dB�B�m���9ͽөH�!���
aF)Lɢ�AY�A��n�G2d�}���_�Bqri]��]�?@~	�� L����d�㘺�PXU	�ET��+I��������5r x�z�/[� �$a�B���2ӳ��|��|*{�B�<z����6���:ce���ٶ���`f���cό������i{����j�w欄g�q�>�����L/�L�1lcC����������.��S5���x�_��Y��n���{�~-j�RA!���� �?�� ��*�轵��=��*:qߞo77�kx��D���)�I)O~��P]�� ����Mm��]�	%!;�E�)q����қ�{JZ�R!�D�'^�P��?<,Xs�=E �r�~]��m,:V+�0 0���:n�~�O��SH�v�����,��NDw������R�ER�(4����綜AI��=p~�4>��J �5�	�2ӔnW1)�E�~��^���^��c3>�s)��3U�bb		��"�*��4��	|���r���Cq��E��p��a�T��[�ď&��ȧVs>����z�&x^�X�@���֮�7�`�=�%��Ï���R$!9(#���~�S�B�Q��wl�Ł��龁�W��lr���VA����Mߘ?��yb��V��8�}�&�H�¢��gEi��.S�@*s�&���* !���c����	 ��)�i߮�~����p4u����XF�3U���kS�N	��a��J�Z!Zځ��)�i����1���epha=���ZF���ƈS�1_4�\�"F�'�u�	���R�I�-VV�fP�@=酪�9'�_�9^��0�ooK6ћB���p I*����=io~�!�?�q��j����-H��O�`/cKw����Ti�ev���S�fjGb3�s�<�XPW.����,>�H�<����n�3��.���}�Y)�����K��֊�U��*��n�����Y�\]-<gߏ��'�z���;��g�}��WM�[U���E�d�����(���3;�a���H?i���%������J��Y���@)~�h=ս}�}�ҭ1�vg���JU�u&�5���R����J�I0�����-�������ϼn/.Ϙ���|}��I�n��K^lYS�H���
�I?����2΢�/S�5.T�`���kC���Ŧᝳ���rP��2ę�)�rU��acsSG�a����h�Ζ�+e8�[�d#x��>L-���ONrb�P�A��I�����)z��U�i��us��fW*�a{�.�_�+j��ِS@�^n��%w�W�qW���I�C�$�v�pB7,���7�������t��e^,�������&�j�n�
��&�QL���s�x�x�T�OGL�C~���Z7�\`$�ԇ.��<���?Յ�����'�0 �u�(go��VF��SmC�"�f���`�~�h���AoP0�k�9i˥d�(l�-���]��-n���Q�J]�C��Nu$m\0�w���t�.qɫs����<����<�_������ܼp-���';e�yk���jQ���<+v1�����7��,|	�+~a-EꋖoG�u�	�cnQ.��x�Fc��+>���u���+*9�>��U���U5�\:u!23����Q��Fj%v��ԯ�̶�F�c�l>�e�$-I�ڕϝ��E�H8�7��r
o�ݐ�L�a����[�`��S0�a�F.;�QO1! 6��5�L4 �#�0�
m#��x*����GK�]L-�$��r�}��g��'%x�����A�;�P���K����V$��cO�W)\~/Y�٩sm���o	��#��* Vt�O�e;�Z��1��%BG���cBX�7��f
�ɦ�=dJ��d�V�c��b�H��HZ4d��_2R�szb1U�P]}�[�t�l��@��z6wjA�}%�$yҿ���RT���an��a�%:��2&��	��~�ռ�m?L�u)@4�b���Y���~��Q18M���DxG�}WdY|s��7~PF�X۰��ŶA�0��Z	���)�b<.@9��۠>1�'�طp��D�2��\i���q�Д��"�}M�ta�|��ٱSK�,�ki)�49e�#��b�L$e�r���l�!a8�q�=_`��T�(��>
��	kv7�[|ě�|�Ԗ�	W�$C`A�Bd�ق�� ������>�7/�S�{_lb��&2�0�G 1�b��F�E�i �	7)���T@�k��iX%9��>CW�w��b�PQt9�E,k4�&b�b�y�9g�1��$��t#��hH�<�Ug�j?�0:U����=����V	Y�I�A�ףی�v�a��vR+?��"���q�͟�����m5)��֊*�p
7 �&�OS]�n�V�< ��?�nMs(������E{�J�L��mX��]	���J+AR��]�C��B;��踆�/�z�Im'?�(ySCH�o#�i)nG����X׭�,��,�,G�K�/@F� �#A6��돊$S���'�=�_,�Y����wd-0 ���Ǻ���H�u�>6�V�]�♩��}ag��6й8������,΋|]��E�/�z��P�`�'�':�:U)B�@��F��p=lE�'7������w*6�8ے�#*~�)%?���{E�3@/O��Q��f�S�v�����Gt��@��X���-p��b��x�$[;�^6�=H��礈ܻ�3ݳKa��������ͽNi����L[0N�iaa�D��}�M�E�{�/'7��B$k���$��y+ٖ �� �!���v��|��I�>D��
 �>Oe�|�W��TVh��Ӯ���s�I֜Ω���\.������,��A;{i���g1�ii�G�"�`��H͔�v�V�(!�Q�y:6}D�b�qL�X:ݞ��t���z�`��|
�fP��Rt���u,%������y�c��d@�'�bp`�����Oq=�t� S�s஁_�fX����u5d ^��L���eB�<τi�vPl�om�8a|\(���ěq�e☰3���rԪ���_���I�ȇŪ�B�|�.I^�\~�8	�A����ҷv ]�\Ý��N�i�M��grDݶc�-��iC��b���2��W@�0SJ���P��"���,������]�����`�[u`|�z:�IÔ`����b�Wf�1�%��c�1m�a��5���/���[V�0�s���Y��7K����[֝���kk����|��KaL#��o_a�ܟ��Pv�ON���:�ִ�j���@�E���۾�^��v��y��d������ZD1�Q��ļ.���Rڅ�c���vС��RJ�o~�,`E|�i0Q����. ��1���Vv07X@ZM��UQ��~����)V�>��N��� ԩy�0hҟwϾ���-�4��E9��&��\Vf�ξ�L��a���]nm=Qtn��*��;nB�?�4����Q�f\]U��yM,I�G���A]�,
x�|�}\�a�/XO�s�Q��WQ$Lj	T�m�{w2��(Hg=�aH��'2�U���/�~�T�A��pVM���迡6��:�3�3��A���z��֡��-��ެ�:-��ȚK"�5�F|1@@��~7Dc��g0�d�"�zC�l�`����k�;�?<�2}��D>l��ت��hD7()����,��?>� �T7]d�8AI[wPy���!`�`��Sw������H"�߶�*:g������MM߳vY�:b�A�
@�	���6a���
B��̷���w�dH-L �e�@�oҴ~�� ���p �oZY���"7�f��q=S��S�dƇ;;�f��z�T�/h��䱽M�BE�Ei�L���ޙ`%V�N^�Ii���b���q�����V���x��'>���cֈ!Lp��EW���_�py����1(\�U����1���a,��pj��@j��?, �@���ؤ�_��=�8fP@� 1< }�Q�ۘ����:)�ҋ���6�=��ik0�g��w�?w��r�ܰs��g�%�)�<�(�}O
2ǁ��X�/M#��3�N)G���i�5�a,�o-
�͆MR'���n�S2��f�im��'��M{	:զ��6�=���5�#��+뺫�J�O�=1s�	Y� ܙT�e$�)>u�%B��z�n6�-/ s���p�s�@�\=`Kt9�+���L�N��ot`r���I1�5�,����B��E`&!+T�y[������II���j@K8��A �:CD��9LY��4!v�,+�_.��py�7�����ft�{��a��+�,�2��K1�^�k�A���,Q���nٺ@��K��q�?y����uP�V�M�o�t�˴ <��*V.����s���#WmJ�X伅�X#R8�w��!fQ�$�����>8Fz�P���f瘏���'����4�lݖ∳p���F:�X��W=X.jW�	<G�_�͓���V0�ɐ��������a(��a�V�t��3��C1GW��0�Hi`Hׄ���f���&����|n���W�����w���:;/����������N<ͨ3O�۲��%�]��".uvl$�˳L�2�F��:��G���淛�&�}��_�iL���U!�:bSd0m`�PI���|���x��N,�7٠{dF	���(�o���hG1�*VeL]L!>�	�s3W�U%<k�<���[�<�r{`��"l��)��W#��G���"�9��nw���L�TS�U�Н���W��9���i��*r���VO�r�Q�V������7��!{,��0.jQ�5[�,:�biM�(P{�>b�V˔)�r� ������Aqv/Rf`�iK��������.���֔� 	L�q��kZs $c5\��X����y�3gs��Na-�V�j��b���c�G����(\-#�S�el�W� �l�u��v�h`qq�Hs�%|i���vP��Z$�����5o�A����ۑ���p�����U�#JxӘ�I	�N��d����K�x�H.��"`�p�?������G��I��G�X���*��nAB�8y^��{ �5����ӷ���4�צrr�B��E#�kb�"���"�C"����͸�r����{ws3o���-5�h@���U?�z��O� ���J2��J�ۚ�ݢܺu�Z����¨���#�BF}�s��q�i�Y����~I�%�����3�?gi�z���R�#܅ܥ��IC��P�i'T��:F����z�]K�T;n�lz�ɸ����J�.4���H�(�.����hi)�[t�a�V�Ჺ�bI`_�_���LR�'�ПYL� c�Au��v/&���lx��DL�dn4�^���`+l�^�}tq�����5��w4�fWq�m�%uЬ5s{Ѓs�S
���)�V~��sw*'F-G��H��6�M�iL�QWoX�<:n�T'(�5��S+��%�.(__?�j62�8�ā�m6P�����L��p�T�y��*���M��B2��	�J�\3���<���WQW;u��0�Rhz�i�#J��4o�?):D�9�B����BۗF�`X���Q�d:h�sBb�SjJQ��)�a����U�(.H]�x9X��~\\6E��r������oL��P:\�T@�Hq�H��:����U����S��m��BXѱ�튾�b�Y�IO��65}m;�'I��l�|�5��D���R�hGK���`�f@;`��+��(6��G+k������	��eY����sүG��q��U��%�S�:^�h-P{�5HW=��Y=9F|�I�щͩC�SD�6NՇ�rQIx�sjG97�Ma��-�[�/���u�Sp_xgk{"�S�1��4�MN�+6��[S_8
x���m>���ȿk��	�2װ?m@)T�PwFO����7�7��YnXSC�+������s�fz<>����j��D�Y	�Gd�{�s�{k�p�᱘w(X`Jb]����o]�H(��nm-��4
�$p�\^��6��y �1�ˀ��UX٥���#ճ#�0�"�b�t��C�H_\���S���Vy�A;8�K?�A�1Hh�9v��ky�D����|���S�ﱥ�ʘd�1OF��FZ����t ���*0 Y�����k���ta�lqce�$�z}����<��7��H8�ܺ2:�P�aƇB�=�h�ԑ3�P��:�x���-�8��mYͭ3���d���O��Π�݋v>��k�'\\�p�|�U��BXw���V��gp�� $�7H��pK?R�k�b�v"��dyv�H���7�m���i�-H�[�נ�9K^�e�tj Bm��DH����{b��`��!�����'|���X[C��>��̤������V/�c%k�x�J!l��8�d�&N����fC��H��_�@��@���E��:��p
�����!�$���Fv�U�_��$&�#��z����75"�Ӫ{fH�n�5v�����}e��/Z`!�Q�{�iWE�!q��f��f5ê���� w��I��f���.yJ���j�q$��k�}�n�A���=W{}A=X-�+"�.�N�$�Z&J7��vx�S�&�f�E���f kwv����̏��J�ޚ�7S��/#bK*h2��-ň�[��0�%�9�08"3��]%uTb�b�`�j�j�@���x���7�U��7Y u���}������9i��.iw���FDqk������o�@<�������jK�z��:	����)$�)���x�5%K�1��qp����Wz��L@������~��<��G�8�G���s��AЁD8���)H8����X�V�*D�.���$+{��;��Y��JZ�+���e�������q�`�e���y�:���]D��pW�)Uxc����DS��	�:��"b�N�Nt5���U1���1Z#a�����v��������+7�b胫�F�ؔ��Yg 2��񜀽N���a��8`��t�hj�� ��$*-a3=C��O�3����)5�J>rʹV�KS�o[�П2�Nx]&5�.tNL^�Y��w�!�(�������w�����ao  #3F%V�^,}��02��vsd�f;�2��\��B8@_�d�[U��hBq��}����G]�J'U� �(sڄiz�_�z�5��:7���v]�@��r�`�q,V곬:Uz�Eg�f�ZnT��B����A�{_;���6[����|+��
�j{�[�0�m(����F�a?ir�As��钙廐�0#�=��f�"3����קgGPI,&��@<�7�?���j>\/A�_=������'����r��`0��z�%��l� z?C✄_%�w6��D*������`��F�8\�p�j�7"S��p4�p'�������*�M�S���`b��Gb'�KDC7u0�:���!�m+�|��CK�sRA:T�dZ�vbO%û7?'���zA/�%���� Q���׼j��'�50Qؔb���j.f�,sr�Y{����U���{#�����nOu������[�5x�C��})�ߤ!�9�_�(�9�o�8�Ѩ�� ���9�b��)���F$���}b�B~Z�p�'�Ǣ���u/_\�R�����ц-c��~A��G\��JЁ����e�����v._3����l׀�we�#?'���yy�|���B�����Т�N�*?��El�`�Pٗ��0'�����ս���lm���)�_�{q���ݹ,�q4t|B�;⊪y�k!�����)��*x��0������_^�Nz���VQ�����{o��*%d��)��$2��@��v�w����D�-�2�l���dL��I~��~RhG�a��w)�!�8f�0�E!�|/~qN�
��j}�P����4��JͰv��k�;��`!l�JAtdd�t���ɣ�0@�?����bj�p,ȗ���X7�|���ȣc�� >u�to��r0��o�tH�b�T���������j�_�+�҄hNv��Ho躼/�e���ߌS�&u�ZçA��*��R	�%Iv�e۶w��%Gd���F�^0%g�4�nC��yMŠbLJ/��*�����BP0�b"AQ����.>g��x�!"���o	�IxǠQ
W�yQ�Ys���Vފ%.��RJ+m&h��Ŕ\�����[�e��z�-3�{���@oc(P1�m(RǞx��T�4���8���3h9�fR�+n!Jn���4(��u��d,�Ⅹ��@!�d���W�H���[�c��!�c#�fmjq@L��
=1]5��@o�@Ԁo[L��ܔ9��U���n��D7��7��$���1�>!C�(7Y��)vw.���3p��>�Z�m8�G�xS �T>�WI��CQ��K��
&x0��I�w���3������].j=2��s�떕=�D#��C��|���p�_�!J�`����\��LP��;!��@ox�Gz�B�e	.�6���K��ݸ�t7b�i������?��o����9��4�ṩ�H=��ǳ$K=:2�
[�`y�1�h�ȏ�(Bz��r�	�Tx��"�#��!�x��y��Mc���jdJz2f��께8c�_����j�""�r֬��~����o\s��pWo���"���H��d����ӿ'�pgޫbI�Q���YL����[x��}���pZZ�9��������^��,�Kj�W���G	�e3ݜ�K�5q]��p'��Me�s鄧�)����=��]��U�B�ѷ5�0�
����(?���Jw*?��Ff������Z<�t%6�J4q���j�J{�VE�'U�G�/_�� �.��-0إC�5�����=섚8�m���|�!�٪�^�NWOuT�k����8���S{�������y�w)�kA��3E(R/a�����I���3X�@���D�N�;lD���e��8�`�D;���ΜWY�u��;�BoԞ��<�N1Q�z�t���9`O��u*c��Udg�w���:�Ha�,�I�!	���*_N��o����r߮�Mb�Cɹ���0����K��:p�_��C|�_T�c��*A�Z]��7�B皅��{-��W��-����~��փ�K)�3j �$�����Ba�~���QE���_Y��{��'l��}=\�ˋt���E�9�[&��<Z�j��m�1�OcjUO��k���K\�	9��8 }?͎lw��jg�IG�16˚8p�{���ף
��^d�ypl�FH�����3ä�0)01X�=x�b>9	��*�v����dr1�$#�<��t[[`��iڈ���`j�g�m9)��c��$������ 3����؛1��Ϙ�KhvQ���vz���o�j�yM�:e�h
%�$qY^P߄���ޤ���bc2���'���I%�!�QYt](���c���p�����{� b�p�i*/R��N�k�|��6-� �����E��a�.c��ir%��,�R��9$)&�z� �����+�L�~q�� e�ʠ���4&�S��*f&�*cǔ�ON;�G?���ӭ�H-���A�ǟ�![��֎4�I����9�~��,=�>���,�}������o�D��n^l�����U�Z�=	hy�U[\�kOi�L��V�ܞ����#�l(Be=���%P����Z���7W&|΁�/eld��:_�
���q�����3G��l�j���9Q�)Mu���!�aw���Ǫ+�ƃ%ɐk0�n�u7�h��L���`Sֶ:kr��e�z]�^T��@�aX�	Y-�Y
B�;�R�<�b.v�X�)�U3�#� m�h����"dm{#p2�t>*O�f	!�h���z]tIy���=5���/D�8R*\�zg%9�P{�~��8? �F�8�q��L��#KK�_k��=#�=� e�	����L����R7K�������;Zkb$y�:�喻�o���ߡG���������"�y_��fW�PiqT���A����:��eo[�=�ĄT��� 	kC�H�Ujp,=�(�R1P�v�[gQ��x]��������F�Q��o���@Vzٮ҃�"7)emLK��%)���몙�GQu���N�e\fRb횟z|b|Ĕ{r(�L���w֭Komg&ՊT},ZZ2hs��>�7��Ɯ��w�p�R���	�,���뻭��$�rV�3�~�+�l�����-����S=����qv��|6T��e��EdI4�D�O4H|��T�z�����a����R#�W�<!�¥�(Vw��t�;0��M�)P\F4�"1����+�������;7��D�V�*��������l�֙�2�R��U������t�MA���Ǯ:�m�4���HI�9J�S���]�D� MӠ#{���ڇ쑵qv�1r&�Qc=w��dBH��؞����P�p����H��W����` )NC�/�$cr@���يјQ��(�?p]H0�J�4u*�n���M��ܴ����0�\7��L�vەq�Hx��$=d�R���9��L�%�)�1�^��u��g�����F!H�2,:il]<��6�0嬜���%j�@���W8&�d���)q�v��=gF��Nl��wB-R���Z��Z�#�"��LG^At8��٧���0��i��ƽ�Ѫޒ�g=�����k��/����$��@T�rp�3���
��>����y��)�[#�Q����/1i��e�X�,Lf��7סZl�o����pdV��z�R�I<��e�y�GW7w�52��x�S8kR,��$|9Ϋl+r�E2[���pv���A'V�3���2ew|XPvj�"�F���)���T���Z���-�:3���8/��E�nu�`<�{�m��B��b��AY3F�Bt�>?xs�Z%�'�X��)�����̌7�k��f����sS���L]����k��`MV�aZ~��
#Q�Y��W��VA��BdI�&�D�k��o�/S��tM��т$d����	6�~�Yx�ԯ+����Cb\�:8r�-�!g����s�����s�v�;��b�I�IICtm�E�
�!���:�T��������V:��K�	ī�X���<o%f�<��mTЊ�
,sƘ2ܵ>H��S�97��mo����ms�����؝���X~C�K��+{�W'd�:U�ѝ�o�lt~�-�_p��h��˿�����A�[36}�����F��v�SQ�ŤR�<�<Oc�}����d�*�6��	Ȟ�"#R�J�e{��&�4�a0����爒�¢�ZAh���������Yt���8�.i�d�b�V�5���͇���g�Vɂ$���1�e5"d��N��cTz�� �N��m#Kd�+��b2f�P���`�-O��j�,����� ы�=R�Z&�s��)���q}��捳��S<�Oי�s�����,���#�%�m�rΆ���t�;Maxk���Z|t}�	Ud~��XۺFL_c��N"������YY���.]}�#_M42�������' ��-E�����G��!*�E�S1��T���� ��s��w̓��S�r��.e%���
A�r�躢���)�DG�&�����}��u���N̽X2&C�^�S��'DG%�H2������W��8�r�zG|A���&���J�ѕ��������O��~pD���wg�yNʍe�t4��!h����ϥ�M\��=?�-LY���h�MR;�	���Y%�vَ�|�{=h]򵤈�wq{%5���\�:l��Yr��&N�q�h%*�W�aa�6���1�%l��)Ҳ�J�{��Y�f���]�è$'�p���ݞ�$cg��_���0#�&�)���l��-ԍ;����Iz��/X�!'�G�}"d��Y=q2j%
z�k�	}:���		���*=�C���	�*�i��E�	�,˅�7�8�A��n1r�,8���! ��6�Yœ���4J��(V����X��lh4)�Mj���%��Q(\�%k��Qy�(����ɂ�Y+��F�AO�U	
heb���P{"����*|J&�D��	J����h���R�0���e�«-�½�

�?�Fvd"�(~:�y�P1$@tj�1�����Z���-�Xu%��E!��y��n�7|��O,N}�ga>�H��7�t�n��,�FM�/L�K�: ��[�w�B?<��5 
�$�}��{���7����%ͦ�艱K�쇖r?� /��>��"`�pnLz'O�Ke�%׽�h
EK*y�٦�ryhǰ�]�$t��s!gXQ��������'��0݊΃ƔTEN^Evu��2��T)d2�	����<+TpY��a]�c;�0-�y9����4���QU�|;������? O7%}�x����)I��ք��/Pmb�p�	�n����?	���`m62�F9t�Z���ܣ�
��`N�g��%ѯ�L֝�|s4�U�g���PV�m�n�!�i濫V��̣�M��!l梈@g"����Bʴ6fA�zP�&3�L�k돾�/,8&��s�� ���^T��W�%i�[04�JE�Ł�'�+�e�%	-���� ����w�:P�*���2�����^�_I��)u�_0���E�I蹫?�����ؔ��t�������	�)��ύ����:����s���۹�2��ͬ����Y����	�G���Y��Y�������v�Ƽx���^/_#N1�4�Hy�=�B��F�_{_�T8�:�7�2u"0��t�-�V2�0��הiC��E��V�,98�{����QR�6	Ҋ����v�&U��DE&����� �
�ز;z7�?�bU��I �osD� '�ɜ��CxնoJ��x���1��:�ͪ���J�Q�2r.J�j�A3��O\���2DI��L��C�I�}�N�����m��Ǧ��t���̊�=��4���GU�̑��ܣ"$�e�`���g�"���V�s���y-?0�|�d�$X2��V9��� �U�MY�!�k�ܯ> ���%�Q���1}!!o���=�0�������f�S��J�*4};3��[��r�_������ޟT�H��0��DAP�B��o��x�hq��)���nLz�M�uo����~n�1N�^`���&���� \jLn�[0}%�Q�"����_fn��1�n��[�@i����7%���1�E�|�BBq�2��1^�.�
�����S�5��HD�1��Ij1ԐvY�����$P<��Sn�Η��h�*���6;b۬��4]k.-�6��e� ����M�K7����q�[&F�p.�����G��y/g�/ $�?�A��c~�e-�,M���Xv),�F4�Z��X�Udqm���Y%cN��V� �w�TSe6�;�f��}��"�?�.ە��!ԋQ��g����@�qGh�ײ�x�x�a f o��m�w���t����u(2�����w�<�1j��2��ZtbJ�j�Y��{
'+5��5֐L�G����뺾�7�!�<���OQ�|� ��ux:9��
�f��ƹ���e`�.L�Щ e�_S��A��)�o4�\'$�;��)���T�O�`��E�S���$�������3؜4K������f���C#���V���{~���I�)��5���k�?ld��[��LO����zS[�
�����6���� zU_��D�*�ru�Nag�|J��$��o��R���F�)e^c�Z`��j���� �k�X���@�G�G�"�a�T#��;{�a-��x��'����fY�cҼ��r��9 ������WBeuM�D�?����%i�[�#Tm&�d��sO���gDƑ��(�4�����j6�c@���G&&~�����N��n�>�����r���J-���6��s�v�v4�ǋb�7 YD
���.bjSB@{rp��l2�r�=�ߛ�W��^c�U��s��]0�t��ߌ�J��j ��O=8�j�v�lvv�x;`� �$��(�zi�IG��#K/4σ?8������} E�����$ރ˦A6�Y�5@�������!��~�`[�L��B�(T=D=b��풄&>z���:���`��z�ul£�7����.-#%\���,��k���n7s���Ԥ�Ii��͚�~�0������i�Fm>��q�d-��UVޟ/2W>J$cA!�a��K��ҋ!�Hu���=Ĳ!���2^IU���Q*,��F\4�?V��7�g�Ď��ް�����I0B�x�`	\^�z>�Nw���c��Ќ���f����9n_�PUGum�m�K�i����WM���8ƜZ���K��΋���&��?��t��A�t�SIC:%�8��$Q���x(L�7�����DW{�^:<�!���]ƫ�L�[V��]b�@��L��W��¨�x�̍�� �� ��BT�����NKA��)?�78�p�����>2+��:�$!�W�0dNɽb?v\��c�2y�L�檩�nV.��d}Y�����4>�����FT�+�	}W�H����k�������`�G�e+�۲?!����"I�l#�S��9:C�CU�Eo��y�\Hq���9�eM���g��`!
�q�&��ݎC�b�h֭��[���#�"s��a����@O8�ĸHC�R��q-./�x1$�O��G���6���3ؑB��b�`#��T�I �Sr^�M�
d�gG�>8	DۭR}��ԣ_��M�O�e�RY�r�:yu͸A>�%>*.��KT�e�>l@N�r
��M�zb?{�Tg2�L�f-�p�FK�NHx���ݡ��nk�C���Yz)��y4}')��樤�Ҩ��K�%Fя�(��J��5�����SqUd�����#��.�i
��P�R�r�qK���Q8�z;�gЊ��#y��r��im)���*������L[B?� �ɿ��)���Rk�õ'}�Oμ\� ��3�e���A��r�6�� 浘���7��r�b�D9�@s��G
��Jk�xU��~x���ڡ<Nvd��-J9��j�m��D�'nC�m]C͇i�*�����Rd���"	'š��6#�O^�
�6Ns<($�n*�����2#$��o���wI���r�����0����nwcN7�ʧjǎ�1���WD��]���mu�$Ջ����Ix|�+��m}i�\ɕ3���FV��[z�?E����<Z4�����U��l�)T= ����ǁRo3),�/J2���叼?�{=�"?v��Pf���`1>�o�C �[��&;T}��K��'	����UoB�e������r*�#+"�W*ͻ�'su᜝ �U;���ϗN�]	�%� �0Hj]! �NAb�ԴUC=�Os���m"<k����<ގ���~���N�����7ե^�J���?��O#X�& ��6��:�\xV���.l��9��į(��4�ȳ�F�S���M8�ы��zI1Խ|j��0AJ�Si�d�A�u�k�Kr��U�����B�N��x�ץ[m�� <K
�Y�x׷+ظ{�<������R�$��T_�%~R�z�q������RT�t;�,�&(�X��]��Xޭ��6�m���k�	���'�%�'�Q݅n����%*ow� ���^J$�g;j��>�-L�/hA.W���55�j9+���3Z�>X��d/N"S���r n$�T��K��f�2�b� ���z;u��*0mP�+�#�G&���0���N@���iHf��1��� ��?1;�.�f��S�UQ�⻡�G�̅#�Gs�Q)+�J[4�N��m~G���'�Դ^=:x�Vi�������ř�޾4Z!w�.��;�鹭��M��V�E��c婵lF�.�o��[&T������H�O���@׀��7�?�����ʽC�?�YLnY,�R�cpz����z�Gt�ז���o����ax��^� ,�D'��f]S.���QrZ �3���'Эs������`'>�Ʀ�7d@�eC�����koH��N����
�`[�H���i�o��[���~�0�g�O�����XҤJ��l���\��,�]�o7��$���N)���xH+~ȵ���.�t�۶���f4���&��E���9�����y���v
h�2�v8_�������[f�;�����S;�u��.�ݧ�IFe(����������d�������֓�վ�^�Vf>�^�w��q {�I>,����\f����JG?�\^�O�ɲ#oэ���V���	)B�خ��Xc�}��i&�Iw�x�S
���N���oQY9Ǐ M�r��P�&+GpJ;��)`�c�>҉����k� ��^��a� \,λr�F�J���t���q��z�4���w��Ƞ]r#��C@�<�J@7��TN��b��s �%Tԅ�aC(8h���֛��kܽ+|c� @����ۢ�tؔ��>�k\"t4���*�_.�3��A4�*4wH��,a>{����e�ЊҌ�c�>W{�;.�nCɜu�Ij+�����a����:�h��5"t2͊I\"�5�̮:���V��j��M�OyDa�(l`�uG��b�J��Wo}�S�u7z9ͩ����A7����@�ɀn��|W�7:Nʢ��CT5zһ�B+�d�����`q����1�c��/g��c��`#2/�-,L:(�[�s��Ǹ�&�{��P"y.(�%P	l Un3+�Ix�dF#aA�	�!��7}���D���.��M��J�)�����b�kLǠoT���0��س��ޗ�h��47E*�Cł�h�YC*IbCjCBʛ�X��A���[7.ω��#�K��T=�522�UX�祖!���Qn��Ffj�u��i��lI��J��Q|,7�dTB4��"T���a���m��C<�c�����;t�����S�+�ۚ3�Qw1��\��9��t����Kj���2􊣗X�{~�g� T�!��Eo�Mgg�9G���qq����h���`b� k��L?�^\�<�nF��ٜh���^c�~�B#��+Q�����WoxgO�0zƷF�eHn���r�i��I��f���m��Ƶ>�BRHΞ�E�86�����N��#	���R%f�BT��.�����I��0=q��2R��A(��L�G9�� 2�m�W�J�0(dk=�=F��
��1v��8�]7�LK��r�{��6c��u�H^u���;�?�?��CS����B���W0��W�����J��@"9�_�ɐ�b(&��po�M�em���=���hՆߔ%�oo������-P�o��j�ѻ��R-�:����d-]���.^�d�έf�.��9X�#����遨�Fge������c ^rA)J�&�8B�:�g?�㨇���A�����u��K�W�u�4��r�-HI��C�?�z���`�$_�N�s�|I���]+~�q�9T����@])��{�|*S5&9L#���4w C�m`\��A��Ӛ׍�r�����iP}�����Ɣ�s8���������1��b��=?&�͟i�n���B�r���3��v�/�0��Nz�'�c�X��L�i}��1va���g]�ku�	��a$ő�8p��U%�Ek*B� ?jB�V�4ٯ���YF��:�8�]X��~��|�
�J�x*:�F���[8�bX�q*��d��n����R8� W:�k6@�{���++�Y�udm0P:Mr-��V��$w�#i��řŭ�[��?@� ���v1�e��@3(�6iρ��B���������c���枹~BA��2���H��+/c��I|��Vx��R#��Uَ_b�g�H�T�!�ge����sw�[�����Y����ND�SH'?��P.}'�}Ʊq�����~��p�g�g�P�/�3<U�Q`��4�p����h�A��]���3�կ��1��ɜ;C�#�c��?\0�y����l��+fA{��Ig�����xu�ؓ��)��ǓZk��Ӂ�z��R�Z�4`��ʳ��s5�' ��T8#����쩞9�zn%Lx�{�)�Θ�d����ܭ����tj�;o7�/���� �Ĭ�Tϱs¹݇9����J�}-���<+c�{$L)��_�X���^Jz͗��x�X�q�4&��E��E�dy2Á��D��D5��&=��H`�8M�m3���5w\"���u MӔ��0�fU@��Q��ZX�5Y��"���ǳ�ɏ6|�#2�N1�BC�hX;��vx[�X�\�h ���Æ����	;""�~f/8��ؒ��w�N�fE'��#�OH�to�.�N�zB00�u���+����[-tP�w{��lL>-�Dڲ��gx�'	�>���Lo���}&�����(j�=���JƾA���5N��$��X��p>�jX6}���B�Ijp��f���0~Ȍ�هb��:Tay\}g�Tι�Z�y�F�ڢ
ϳ��y��6�_%�K�S,��;v���<���<�[�
�k����*�/�~	̷"-�)b@��*)l��!M1�!B7���).A��FT��|�r�dER����=~*8�3#_���`�Dި�-ިj�U���w%��@�_�_K=���%�
�����b.\��⌂�5lG�(��_�f�G��m�-��� ����x��.�-2̓�ĝ(�tml��g��5�B54_?��߅��ޠ�_�j�$��b�wwfk:��[~5�%�!a�K�U��%I�'�7�ҎX�+p�p"��ꎷO���H����O����ۯ�7�JibC �*u��IoZw67������I��6�A5��BѼ���Rޮ&!E���u���)���^5��uv���N�i�.�*C�"S����'Y���S��2i1W���ӽQ�1�f�d��0��}��G���){=N3ڎ8A�L_#r�c -�]����"`B� �����C���$�|D���=���E�6�T�2�ö �
V���yd�=��7��"t%�oQ��S�j����tJD��H���-���	�j��!q���n��b��i�����5�S�.g�+80����{���a�.��b2��K�C{�?�{#:��"[JÑ�x��aI�<�\-�m$�!��B?`�X�&�g�.�z�`N��+�������������6RJ��.���U���2|�P��m�q���H��|�&�f�8��A��������Z�d�Tt�*�f��a@Ѫ'��۫����7���얏-��i�م)�x?�D `��/+�W��t)~Il