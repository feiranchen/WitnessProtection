��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�5��3���}��8'�G�㠚�S�L�C�L��I*�5�4�>ڎc�����I�$���*�N#[jlg���e�gv?Ɠb"��/��c4�}���=f0��@����*p�i���:!�.�;������������Xo�Z�>�[a�����b��_�H%M8��d|�54��^7s�"�tV2z2��C1�7p�jH���������O��\|x�]�K�A��ψ%�p��������c�r9��z�1�����ff�Yy}v��m��n]�ǩ��Q��B�\��l^Q�l+oj����/����*iM���z�h"��A)t���l�[����Q�%b����,���R\d���Ҁq����~ׁ'p����>� �\��`��ă:���5e=K:yRR��+e^���^=3�ܤf�}�>��1Q()5t���S���#|�@!�k�?�8�2���ȟ��k7�ԈY��jV�4\[&��}�|7k�]ƚ��\P>�u;�7��o�D�6�JdeE&
K��YB(�����{�A
'#�4�іvƌ%Z���3B�&B�װC�zɯ �S:�rY�>?bo�kދ��yuGɬcy��ɺ�cҚv{^-�AF!Xk��Onq!iQA�xσ�n�$S�zL�A��JO��a&��.
0{7�\GY*h�j��x�#�#����-�~��E��y=B�Y��u���F��-?��[`�ӳ��_]���} =T� �ςNfj��j����\�X��m��|�X�텎UH~�H2�g.��E��&c�L.GGy�H�l:�M�)"A�j~W�(P^�l��3�F�z����!Qg�mVN�\0<J��4K�����_J���IS� ����V����	������K��C���P�@��Ϻ�=��A]*	�� i�i9�07P��|UͮcB�v�>1x���9��T��Ʌ}����sC5,�8��ϦU��q���ʂ�e0)ksiГNk� 5P���Z+J�"�,�M�73��0�N�a���Ћ����ޞ�
 N��nl�� �b�QƁr��z�
,�:*�P>2�U��RN8��!6��䕴\�E�?g�+��$�p��(�*j�$���T�>�F�$��9r�S���"!�bg�{�����|�.��+�-�^`�7=��W����܈EL��u���x��3��^,�F%G��4�9��m��[O��cݫxV�@	l��J����|�{PmZ�@txf�o�G��{���1՛1t���R��{75�n[������9h��N	TO/�-�2X,�͈�?�L�`��2:I\�ba �m��a3�2��yHs�O\��\l/�97w�`/�)`�|�Z�G�:��JjIa�cSJ���-�֐�	��кS)S�:IIp�tl�sm��OKI��(G�S%T�5��N���}�M. Z�=1�L
I�(����S�dR��$v�����qp7����|2,Z۴ �4aW��!�����ѽ�u��7�(彡"�!�d�d��S���y� 
b_���+@�>0��9b�uU���eS$�)1�@u�Vp��u��S���>tm��HG�ӱ/Aოm��Q'}ՇTu �A�W�G?���T��0c���l�I�A_�=[�v�����'@�mhOG�Q|X��?�p�{���L�W=�f��z?���fu�D�;�偏���yqj�3��Apԡ��;�����M2S�$#'���k����mE��>��Z�M:8L?�I�a�nu��|"L�����S�I9}4L:c�U0~i�,��xI&pg�@qx�Y�+��6� IA�ù��VBs6��\k����N�^��P�����������C/G?�%O���%��#������#����b`��먿�^���Z"
ÿ݇狼%F8*��r�`Ox��?�z��к�k؉Ж;���ۿ���w�4vr~����ԛV^�Yik�K��ʎ���Ϙ�?\DGJa7�9#ƽn�蛝 �>|kGA}�bۺ$px&4_�ظ́�̅��ξ�bf�5��V��8�(!LL݂�@Dc��4�uC{v�H\l ��=�L�&�>�l_��!����H�ӹ���y��=J�}t��,.�&*���@�bZ0A����hu���I�F ���S���1$4> ^��F>TDFڲw�@>�ALjѵ\���1!ő�������gZT��Tn��3V�!�d�C��l"Q6*6��ʞ�v�)̓�PW��h��<ٗg���1�è�1����VM��1���o� �u�!o��ɥc3Ғn���fm*�pΧ��`�e�%�e5�3O����.�-M������i�;���o�(ee�G�_�O��'�W��x��`ݱ�0���;D1�pJ��x�l����z0�i��	ԜR��ퟫ�����j������J^[Tu��X� ?�8�_�"A��
�Sv�e�eo%�ǡU���(�'�s���%
#T�\4gA<�]����s�1�����e���!�ʓ�g��ZFv�G��2
Z�ʥO�7�J4�/�r�1<�%GFO[��UC��|�vH"ǹ�`#�wͷER
�C%kH$FR;&�"���H')C�ץ�r��Gv *��Sz[>	��?��8��!�=SÍ<�I� �L���d�2� ��Jv�5r��ђ3%�Gj���`��5����j;��ɼv͡�>�y˨_��mJE�F�8�dL{��K(��-l�!bs
��������$����R=ՠ�F��k#۴�t@��	`���Gñ�G�d::B��hIw˳BT�������T�K%��M]�u�B�b�-f���ȷ����̊>s����L���̴1I�z�`⇭���&�7�q@���t?)���1���F5g�%�47'�&����N��K�Q�m;�3�A �>���e����0��s��~d*w�5�c��
g=�c� @x�Ic���|�1ϳ	w�5�1����b�-�n�� t&��-;�c��vVѶ�~/��`H�D�����𼾦�&�͹�l��TVQ9k4�^��6|><�9��e��GU�|�8�/Nr*�mݪ�t犿Ł�R9{`ǴI�bş�jx��|!Fp���Z�X�b2Oa�Hn���owAA�٢��3�$�k[�q�	��.��"<%w֤�pMDȧ���J�a+�+k����t����xY�U�������R�PB{'���R�n�e�"�IQ�٪)l�uW���')����;��n��ɥh�	B{�Vѕf0�S�pe�-�ꂔ�b{]��2�V�HKޥ?�f�c��q�ζI� ;�W!��t|���{��b��HH�p�%�� �h�<�y�U��b+���Z_�e邝ل���U��q?E,&[�aI�↢�E�Rق�5�/\4�up��n��<���x����p����90Q8�@#�����Bu࿶�KZ�b���aHTb��B��G�� �8`ev9Y[����׊�{e�^���G�����lS��L���q���/n����,_�|��ZU��wz�tPNd���t��8�_��v��l��M8�gv��;p�}��`҄���21��%�d��^TA��%ј4)�,����£c��,�w6�R-n����l&�~�KO;T����n@��opJle�OΧ1 ���[񎦘�s� ��"��z�3&����j)�i�MZ�gP�y�b4�;M����28��6�(�%;�U�ta��5y�]$�G���E����/r~��q���I�HT$�5�Y���o�-���ٖL�� �����+a�>��`�8I�R�!�'� ��uN�E^��U2e~>oŵƪtL~���_���Y�3�_ڒ�r�E8��ݔ[�V�
����R�|\6ǯ%
���G�H�l[���OY���3|gf�}ux������]Y8Γ�\B:��gU��Ź��JU+I٠&v��Y+a>���t���MN���M�b�&�3��t[�F��:��KPx!:�^������rm\S� ��+Q��d-��?5	֢>���I�0�b�a�fn7*	_���K�`�x��\K����c|�i�q��N)2�z� ���ć�\o^���0C�R�@�9�=d�
�2�e���G��?��}��P/6w��I����!Eu�<�r�s������,���!�_�U{�������8�P1D��v!��'�߹.�m�������~�>t�/��NO��g.jJu�q�h�|�o����}��M[q4K� M�n��K&�Ɣ�[�7i�^2O\��:m��\�����*u6��2�i\]Xp~e^�M&�)��i�4��'��5ZHh�N:����+Փ__�\h�8���g$�2�P�x��Y�?��ic����W	���H��d��ƨ��.=N{����v�z��]΅ҫ�T�Ҿ�0t�?��gm�#���j�~��3�Dˌ'mmsN��8�6(��/��� ���T0���6'�sڳ���e�rZ#i&�������t�^��f�̹�U�Y��rۥd�e����}M\*Z}jҼ�tF@O�%"%�2׍�Z�E��^��c �"�[����*�ܹ�ہ�J��WH�~�4����ǼQc3��@��Y���$�.�G��*E7���\5���ЎӋ1�U�f�Z\����-@_����]/!P)�I�Q�{H��#����jЁ�z�;��S&�8��o�Hy��hf���}�¸5�����sV�ML;�͎9r0�6=뎇O����=R�|��%?GI]<�����Gf�}�O�n�9�����2v;S)0�ǁ��X�;C���ہ4E��m]j�.qA;�S�-�$�y�E����i�Ř��OH���e������>�,��I�c;�N�[��
���'���������/p�b葼5�G��$C&��8��q2���ebo{	���V5���s�E%�9���U��fݹ8��[�@L��x.�Q2?Y���`�+I���9J�GJ۫ʱ�J����}V�](i�u���(m}נ�ߐ��02�9I��VO���SE�3��n�������ә�^�P��&��de>@���9�����G׼�K�=��3-L�
�(��E�` ��O���?�t�o�.썘q}�*�Q���߿-�3R@a7v�X�%]���o�v��f���嚿t�����S�� ���E��hn�SmFU��#Z7I��$%��[�_�����H����JHm8mK�O�L۟������1NXw�z`��[���3��a��۴]8��]=#��%��1A?v�U��~&�IL�����L~6S��>���M���K=x��K ̡�V������cRfI���\�/̟�7 %��)�؞
aC�Nl���C~�1�=���7F+�qۢ��?����
߆g�D~�UBG�� }[+\��s��5�F�}<0mJ��ە��Pb֊��|ڹ�4�!����F��#�IB�������J�i��Ő;z��	�mZ�# �������q�Kk��L$��+��H�DQ8����V����E����ws��a7H�6#��[Y ,���>�sv�r�T��}G����Pw�,+V�"��P���-#�~(�s����3��oa��%��͇����x?�mRdO��X�?e�A���x���r�|�w�Qƺ��Z��u�� pi48�T���n�TT%�}���o撐�A�f�j�M��	h$��I��E����lC��"�09�%Ż5�S���B��z�o�ٲ�y����{��m!cÖ�I��c���D���:�G�Y�k���%.h8?z�����M����_��C�1��^!�H��EF��ح���6��L?�:m��\�(�5�Ic8�H������qSQ@>D1TPog�j����&W���L�,���]�u����ޗ멈܆_���S�@��s���G�G	���Ԃ�~̓�6�
���%60�R�~��m
���vsl;�`߅5M�7�^���5�V�s?��r�gAc<���?���<kM`�8��G���+�qD�1�LEN����l�v)��A��~�՘D�y�ST:|z����X�G[V_�c��Ʈa��0_����[������`�]��I���@)�neD[ٓ��{�>{�^o�S5į��.,2�(@��?^�Κ���en^5�\��q��S$������Ѱa�?0�Ϻ�y%��K|8��uzs-t�c�/`�Sʯ*�{#�bX�p��Z�2Ē�����.�r}
'��H��"w����e�L��l+�'_7��H��xqդc�SĄz7�?-�q�T��i2;.e�E
��1<x3&���R+%WZ`4q���,]~p����?^m���o�����y����y�R[�EU%�1ngb�e�S�(B��<�\�'~�mC����|p5�7�}����ˈdb�!��ؔ5�g�}�)�9n� _s�<\�w�:o;��;�j�QOh���͂ �= 9������$!Z�.���R<�kY��8��������Xv��.�=����>7y'{_�q(��ߡ�2U{�s �7�,�����	ٯK�=��H��韗7����d�slt�
z �:P5c#j�g�띱r�^JZA>��?�D!��")�a>A�
l�����^�>�:?�:���'hf�&�DT��7��1@M^-2��ݪ5���eA4?��,�-$.���$:�c�p��S��
�_߷\ϻ����)��
:���n��+������w��+~��-+_dG��@�,�wã>�v_�`���H`}���*8F$=�K0��ND]I���\.*��20�UD|�~��'§�V�z�F�zdLp}Pp��H�4���V�F�O�X����v�Z�塴�LMf�M�IB>��M�Ʀƿ��>Z�bPd�Z�����t>�H"�W:W~�����_YBr3u>Y�b��k�,	J�75��z�U0[��,�Q���F&o���,a����*�߸�f�2�ɞ�_��Wy�_�I2T����^�7=\����Gz���4�TD�r���3��[#*S��"���vcr�^�\�iEp���g��A!�
�o����u'��!9��w���A�v�eߓ�i��0�0Z�a+�>�Ŋ�j�v�n$�Zfz��k�Y�=u��?��俸%�D{�(��j �{M
��Z�	��l>�8�6� �#�Q0x�X�B;���u�9V�g^�I�h��q�NGw����}���s��������sś�=L1¶.�l�Ӳ�4[�gf��:/�z�m�DԿ��Ȭ殛#�5��-�_�T���y���\f��q���+��CM}+t�r��0�~�D��{A�z��8R��~k����n/"{f�J�Q}�&�~�5$W�oa(2��Lj��R��ۋ����7�}���RS��Xp&�Nߢ�	9��������5qG�2�2MÈ�SǙ�g�f1��cxÄu��0����N�0V@�19>�5>����,�����m����2�4J�q<Oԍ��Z���k�!�`.I~�7��YsH�5�a�`�.�����*��2T���^R[�/���^��=;#�7bN4���%޷�2��ʘ�" _��ⴐp���8��x��{�B_"������X:RB��V �{�j�@� 5�����ى#�Db&���>��	?0�9�p��=��Q�����Y%r������ڇ�QE�R�����(��W��V��v����5xj{J2��ÿ� f��� ����9��z�+�,v1��	�-��[59�}��o}Vd.\�HӸ���U�w��s�V�'��A��%�8Ŏ`�e������K�|�סr\�[�E=W�3��j�)i����r⦙��
�ȶ�L�#S�i*)|x�k��'	X GU��W�n���N�y��S�(&2����98w�=i��'�K ��*"57����5'�Գ�7��0�j´"m��S�n�E�~?�c��^�V�kL�@�T�v���l� 8��0]ѫ�3�ǀ(=>�g�Á��d��e{�m�*��¼��@:�7�0��Kc*��@�;��ť@��5 IВ�mp��4$t�s����{W��&���� 
Q���>���&��E�݇=Ž�O�9da�S>O�T`�JW}��YwAY�P�9~.��X*e��8Һ>LI�0d[����$�c�Fz�B��}��Ҭ�)�-r�j�}yᖳ���QW��l�+�n�%N�m��gH���`m/"Ju�n,WKL-�W>�e�rU�Nn��t�b���VLZ���Ȩ����-��9Z�u�+u?��Ư5�![�������jD�j7�
u9Z��uGy�u���1p5h<)Q��,�"�u�Y�E/��&����-����/W���4�g����p������Z�^�W�=r,����p�3��$��"�{3G)�=u���%����y�V{�����cǯ""���L����]�������t2u. En>�PХ��� 9�zKxO���~�b �O��JM��?Q#&C[(��{T�h<Ū�P���k���ۈy��1����|��6Kۗ�'2Zgus����h&�A��9���+���ߍ7YX<	�(0I��i��Ԅ���%�0�kp�L	�&���"ŉ��5Id/�W��L	���������k�X�Pբ�׭�ݰy��"�n8P*�����MV�*��l̅�����(�~k��亙�!�J��V��y���ڔ)�,.jP�O3�E�ݻϨ>Ҙ�a-- U�**^J�Kzy�����Z	�D�0��*��͋F*�&��9��:v�m$i)�)�#rs�E7�]A���E:��u��&
A�M"'l�_-Zh?r�7��d߈�z9�3��Ӟ�J�)-_)@��$�|���#Sgp�!�<��I�2ȱ�)͗4AQ�%���^	��y�ZJ����mY,��l2JoB�b/���f�Q��F#����+��84}��Ѹ��y�wи㢎� �5�}ܚw�;�~�4#
2*���[tŠ΅�!GBe�5h6�O���m���XO��Z�®�a��\ܜ��Z�U.�Ejq���Wh�ҽgm�2�s~�\��[�ԑ���כV.����*6VE~r�n����|���GҦ��7�o�x���R��~S��[���6m<񃺫���W�v{��òd~eHpx�k�J	j� Fq[�+�;q�(WFr#r�VU���)ʢ����Z&��<�gC]Dֶ�'x���9��b�X̝�Nk��s-���G�.^V�Ҩ8��>�@�{{!������FV�;�&PH��tʉ��=���@�R=� ��!\2E���R�=��|��(�ks�)����j/y���L�$�V�U���{�v�<�b�����g��%~��2���x�uS�BMM�y�x����򆍴��x����(b謣����;��B[��O��𜍺�r�����E˸��Ѿ�MD��:�laɸ��R�,�;�6
$�pK�Bᚬ�z�ðݵF�ɛ�b2�-R�
����\%������q�����j=��
�i!
n���/��Lɛ����4Ӧ�*����O�A��$ӈ��l��� �t�,	9�"]�c�����H��`��y's�W�*I&��g(�F�?1�7|��:��0���)KƲ�*�=锆��s�s�Z����Pc�N�pY�j�̨1��-��JO��5t@3���g�t�(�&���Q:��FG���Rpg�6A��\�|t����![��0}�� ��V:NNϚ�p�&n�ˡ�ӝ�	�����=�`o���s�hb?H}�e��e�'[r����:�)����.CDr�ڍ\���wR���l�{���<j�t5��`饹%�������Z��L�'.Sd�Ӓ���o��.�x.�x�9_k�k���~ǒU�7
D���(�����*�J48�fP�[O�f���*j�m����"�(XC^�y��n>2��y��<%��� ��0���g�sp�r�_N��KO~�� a���4�j�ЗZz~��!�k���=��7W\�O���	7?�'j6�/��Elٓ9�1OdQ�f�.��Q)6#)�k�*�*5f�)��W@JD1LG��~j/�ﲞ���xC���O�n��qB�����^X�K+�)�IvH?aE����'����+�+�_���6�0z&$�:h_a����\En���@� �����P5�p�_��t��Vc/ܔ��.�Ĝ��As�w��T�����k��+pO�jo��MX�SD<�#�?i���*mS���WY:.�`��Ҁ]��9_���:�N����	B]��,R��UcDv��^F�k�5)z8��H�?[� �~r�9��fb����{���7Q�~�-�^����װ�]Ud:eH#&��,\�T6��~�E��%�@5��>��G��Q�ȩ虆p<Kg$Р ��gE�gܭ{��.����?��8�26O0`թ�?�9�n�N�35-����m"�)������F�Т�7��N��c��G��<Y���lƛHKD�˃~�ZMhK�>�3S�faɮwT�d�g3o9=j5�`a��?�V�
�ӕ�"�b��g���{F܅ٶ]��Đ;���I�b��Rޓ� �di���=���b����[(�`vU�����h|%5ꚱ̽]r�Ej�*��;�e�呍W0�X�TՄ�R��5�6��%��"9�nd���e�?���ӵ��~xCF`�و���	���΋�?�
%ldF{P�(��!`�D+{���X�A~���[ݥ���We���i�GS=�.�Wg��Ã��=��F
_`A���X&Ә��εH�q�Q�՚�	$$�y*�y��h ���"g��x�/Y�����Ư��;����Q����.}>�S)�0���F^]��XMYi��xX�)�Qs�.�Wp��Q�(����2޲\i3W���m���Q�}KHM�r�-���
���\R_%�}��/$�r��N{��GI��e�L|�و@$��`�RTo;c�?�s((��=�2��J3��pE�j4w����� Μ��#�~�Yt�?��|�o�����o^�/�9g�3�n>׾���0*�>$����8Y'����uW�ȴb^@ 	�a�q0ǰ8q2��$���n��K���BߑW�Π3a!���u�s��"`N���ǔ?t�-����*!V	�J�M�:��Q�I�CD�p���J��&q]HX�!<�A�v�&T+��Ԥ'z�K�.���eL���:IE�ȴ�o�y܀�����
WS�=�L�ɛ�%ʵ���߶��ދ���c�7B�Y@��BB��𹓭@���
`o§�fg�Q�����|m/����m���n��=���u�����c�t�Q��@O��	5/fw]�<�|\����Z�����g���BD� %L�2�n��Am�]j&4e���B$�0a��y� #��#6)Aɶ�=n���f'�PU���Q�e�_m@͎���OQ ��ɧ	>�a-�E2r��v��� �Ƨ����.p�D{��5�4+�����V�ʬ�b�o|����^r-A:ӆ
#�$�%���`z�`�ڞV�@��@��-I�C�vp�s\���bN͢���<�:��Q�z$ǹI�-��!⯽��S�G��d�����rP?�2�h+�,;%��]Et��_�^4H��\��0x��ђ>6S�z��˟�A�q�����lƬy5~�<.��$b;}�t��
~��7��$v��c�۞����i�og&���-��g�k��.�[m�o	Hl7ӕ�w����>�֚���R5�`���vj%]-�=� ;,���_`�1O/�A�n����@�����F��\���]`��$©{��-:���>�PBO�Ǟ�kFD��^G��P!�cP@9F�?��v�r�mTߖ,-�����3�>ݘ)e+t��	C>7&s&�ZE��/B���4����σ�륽�������]�}"�d��1k���Y�>�6ӊqH��g�yM��<��S�Y}(pZ6r-|��g�M˗�C���|��}ܽ���9�<D(���4���\Ū�瑓q2��
�¯��ZybS������@�JD �j�D�����M+�b؋�TΔ&u�*#����@J�B���o8�o�o�Q��|0�� �5�Dr���=a�:W{�����F/H&ӓ#1�[��c�6P��j� s;�4��45�/�'[��0ʦ��Rz^ �>��K�[+0E wg9M�״�O�~���d'���fRns�=-�w��"�o�ظi���X.HX�V-.J�ԯ��m��w�BS:S8��}\�!#�͘蠦�����w���uIe˳�|�z����,b��'[��9���pf� bi���?��o+uuS�n3�ޡ�B$7Be��_��46b���!��n>���ń��Aq��D8���z^У��`�Q���UĚ��7����a���M�f� k�~Dw���^<^��m1ٙ����dع'x
؝�Jgz��s��l4 /�P��r��E����Wo�.�kP�����F����33�n"�kjK�u8�WA�x/Yq8���T�u�SUfL��^����g<���Ӊ��a���^��u!>,�#����Z���4��˝u͡sHĕ�	���П��.�$2���;��.�����]~/�`���}I�b�Z�F�y�hOr�r��)"�#�*-:NAp��?�ꖤd:�Y������J��v�=Q(�;�~�]�P0-� ���ѩS��1�"�؝�-������<z��=�braٓ���@���֍�g���s+eR�fd�f�3L���(�s�8��hC{�W?5����63��:�Z�jGj��6��n�����;}P��K�sM� �bA�ڔ4P!/��\Ҙ�]���Et=��҆f�A`5���7�6��w��1)N�X$�ق�Y
�Ӈa�|��.��,J{Z���CE�6�g��87����-��r�i�%�U��g�
����P%~)�"P̔6�2*��J��m��*��9=��S�!�z�V8�J;�)}u�О`R�_Qe�uR*`��MNs�h��i��rH��C�>�goCF��V�=v�7﹖. �]l=q8ft���:o vO9�ς�X��-�-5 W�'n/���/�A#eX�K-S�� ��+WP���(��(��s�=L��T]��-pW`P�j9IG�B6oQL���D,���g��v�z�k�X)p`"7Tʽ�.w{���<����0oU���u:w��/j?��)�t��3@Nj6��I������oLj�9��x`q�D���:cl�tB����Y1"Hs�4��� �ڠ�},�Y�E��EPY�X���dM��C�JU�M����B1�����g�e+��C�V���늚$����'�+œv��ycd9Ez?�ޝ��Lg��A�!L��j"��Xq�cբ�ҷ�	����a6��ǂRa�<���h�^+|D�ѭ�N���>�*��˱o�g�������W�;/��B��<���v9p�R-�8E�`T�z���!�}/�^��;
Ӓ9߂c�}�s��Q�����dU��ʘ���V}=.e��p����mm���� ����l��8]�����sSh�nR�s���],�R,hyf�B�h�v��0�[]�j�'��Sնtg�͟��J�Qp��-��!̇�%߀�
I�ɤ���^��Ё�p����Q������B�D��o�h:Z_�0w��jE0p�N>Jڇ��k��>�Xe��Ak��O�1�+�x��h�2'iD.�F�q�}�r|�x\>�˚z���ſ�s;v�G��w��O��l_?�}��\u�)rEJ�7T�����%<�,��ۏ�.`�-���Z��s(�Y�L�]�4�hM�Z:�(�u��
#=$�#��ԍ���7OQ�7�B��r$掘IQO$y̎��.u��R��B�+.�G�
���\��|��v{آ�D��J��KQ�2٬#ǋ-�8�����Y�yOk�q[N�j��G)6�ȸ6'#��l��0қې�i�6��%.�h� �ъ\x=��;܋l3 ����j�H��x%�J�#�X�� �����7�8o�W�t�U��V,�<�&E���N�@�O�!J��f��9���#��fsgRW[è�$H��BaX���
�x�f`		8��j�C��Ǣ��4��{�L�76yPE�Ѓ����n����8y�lFI�P���߳��u �/g�J����X+�����	q��s|zX��~� K�@�]N�-��	�}'�kY��k���#� Y��D(����?�u���C�,e`�z<{�cY���e�z��?�^7���`�.��Q`��DO�R\7L	$L�u7 ��y{7�C�d���R�vȝ���7G��绐�$�_�x��f����,A��\eޗ��\���S����7甊>�c|�!u�ά&��s>���x�M"�I#NOI�̕{;�"��._��7X�F�\#�BT� 9��qj�|���lm�|�[%棉���J�=e�y��'�|YW�(��MF�����˅��,���;!�?L*�[t���#��$*n�/�M�	[ع�6yD�͍�{n�U�B������NE:� �˱�+�MGݥ�����ǃe��<��b����/������,A�w��!-ڦ�'�m0��u�w(�/d <�[�+���(����=-�c%!��������s��_� ov�yEI2*~g��3e	��sW���2`u�kz�,D��ӺB0O������ "�-{!d�B�����i�qc{)���Aқ��#�Ku�b��A�}�%6�쫲��:'�C�\�8/c�!�$	mg��Y}Cι�W�܉��pd�M���<�^�"��������`lՙO��߳�(��3��������;���x��bK�ÙF��oK�X�}� �ܭ|B��%SAEٚ�^�{i��x�JVX��I֯-��'\tZ	�y'��
��	y�DE�^��%Wǩ�%�c,[vz(��$ǔ��_�t<��]�X/��tb�i��d`�r�]��Kv����8�?/�.��%�{�v�2�3�{�1�4�! -<*q '���P�\f��	�E���*�\��^l���e$����W� bj����Y�R^gPH�Aq��YB��j�cZy�c�A�<�Ө>7!��ms|��HѦ�s���i��':��y��y7�V뫣��)���>� n� �b3|�4���g$Wye������I��H���&�����VB�����b@n垡p�N��vl�u	�q�����DLݶ�s�C�����6��O˰4��K�_qʽ���� � Z��΍݉�P��{И}mD�x�Y��m�
��"�۔7D��> ���s�(k֣޽�ڎ�$B�*�H�[�!���t_�)�&�t���*F�ʤ?d5$o���{c�~a>�Ic%pL���:�Zx�uJzA�{<>1j�D��]��3���0�1�'��~cL�/��gN����b=W&���!D�\�"�!�b�<FU��biD@ߔ�6��s�JBОGb�r�
��R;o�R7�����4���8=��#�f���q؏�U�F��/�3�T����$)�^�i����9��K�a%���_�jA�37]Ab-��N���d�e�i��Q7�D�k}�a��=zo{7���c�QϬ%D��N\��`\7� �mL��9��H��,P��d��u�}OK%z�..| \�(/?�(��9xS�����;<E��M��=��`��K.<S/�\ۂCUecS��a�%���D�C�^��!��ʪ���I�g���X�1����@7F󺘛���|���)dg��m �\��O�;J�:�cU����^���mN�v�Հ5_��}�6��3 + o�����m������t����[��+��v[c�	����N^��Q���J��|�f��؛0&:l�'y�]{�YLi�:��qΘ_\�����<Wҁ�N���qY��/9(�B{]��3J�x��n$�&&ȴ��I�RT�2���Z|x)m)Ch������t�t��.l��1	=X�d|�(�����z0<�>���qs�V�~��w��,��d�Ջ��7u���ޏדٲ"�v$ͺO��F9~�����o���0���Gsx�u��K��e��u~��|aJ�i�5*ؐ'nW��W"��"��P���:�O����,D��r�h�,$-^VOj-��,��S�l���ԕ�]�9T�\)�s�1n�u�Dґᖭ��\ЏΉ|�\
$M%5w�SL�𛙄��K_O�|tl�x�E���.�Rبn4n!p���5�XSLt�l�r���F���ٓ-�z��%>�4��cM�z[d�8�x��F�Qw�Z#��U�+�@�ڬ%KK'��#o��h0���$,V0"����'�k}��ǈ���'E��Χ�=,��K��G�kR#��1���ܒ�jp����+^d!Ip;(/�~�H�XD����#��ʟ���;��Oò�m!� ��go��]���0@=R|7��h��ء"[�t�gc�J�!�m�_c�eo+*�	n�[P��pN+w#��i��v=v�v���ښ22Ͳ;��h:���L���@�N�w-�3�pה��������_�R�<��(�Y��jK�L����)1��D��Ǻ*x�S�(���6�|^��#�$#Ҁ4�۾�=���#.�ʻ��Rˈ�B:Q�_�)h)rVr��>;Z1T~��t�sD]+�
�����3n�>��zd�)JV�_6�TZZm�k�f���I�S�Y���%)��
�����P�n��Ry���*�4�i�T��fw��_/�qe��8�G�*/W3Elj+����-
;P��.mv�� ��+�����H�vaZ�Eu(H�оn�omxx2�0�y1D�nm ��7^q�<e��:)*2N�|Ra�IIGKn�oj#��A��c���>�a<8/��.Yq�_�e��z.����F�3!���A|^ȶ�a���̤Jxh�6<Q�z������l��������<��W-�k#��8
w:t�\����;����3�3�#�n.�v�3�õD�qdP2:Ko����Ji��w�e���-��1���_�"�~����9	�!�`�%b�a���t4�42[��_�2��xJ	�	�bc��:�f`Ǽ��庮�����:K�bC"����EL��qk�o��E��d �ӑ������k��z
����P07�9����&���7d��V��ʧn��fb�Hh��*�C;�������E+lbq������?�a5a���P��:�����Aw�<�p���u��ա�(}ˁX����b�LDlҮb4��}^�P
����#5���SM��T���[�2e)%�E �G�$�/%Ѭc�ށ�f�$y3s:YU�F�±����,��L���C�i��}NU]#4��%�S�d��O�O���8.�_Y*0U�a�t9�����.I�16������B��%pM&Z��� \���T<��j��ũ|h������\��@$b�(U��g��36���N������,BT��T�1��eo^Peۡ�2{f3v������qR�J�v�R�𚧝�wH ��3��TFoSP�G�6O�>�%�ѭ����hR#���^�
�o��p!w�.����{2����bFv��cQFQ�O��Q�>S�|��il���rJ������r�Ԟwa,K2��BbP� �$���HY�� ��̜Ո�=n�G�����he�Cl.�UL�z���e��,�'�N��v�t��(�B|
̯*��|�W�۞����p��=�Q�E����M��G�I��^�S����!�nġ�׸hk�
�@���I�4|�'����x9��iVn:��HL���˻o�6\�� oϠ�D�����7��;��G �7��Hv���
P�����P�����z8�7ڈr8KI/A9�0����[RviF4:\��~ρ��ކ@�*��cYBf�_�����1��\�ӝ��>%j�KYj^���/�	��"A������Dk�d���!�yO?m���@�f`��~���,j�1v,��lj�׿��gt���%�K��0Ԩ{���AFt���'�dZ(b�ߙ[�l���3�Z�
'���ڨ��ס P���N���StF���Z�5>��"4�k��	qn�2|��`�Q����K����1����,U�^�U"�5�|d@�~�$��4�eQ��͙>���w#���RC� -���ٚIV&�������z�ᱷcg���)��[V�z���\���he�A��+�GE �_t�=L��� xZ5���h�[�8�Ğq�7�8Ҭi�kSSﺺ�b�,�EI�p �4���v��e�N�I����'WYؔ\),|D��:@W��: <t2^ ��ZR��Q%��R��Ɠ�@zo�8��Zπ�{Vy�䰾Z)3�AG��m�`�v�[i������,� ��K�=�4ţ���X�~)�F����Q�=C�<c_ho���i$B�:�&*G,3�ğU����Ӎ��d�c���G���/cJg.W�u�m�;s�%�QRP�'��>y�p>6��Uk��y�$^������Ky,��&Jp@c��]m-�S��5{��rOC�	A��R�,��A[(B�O�tA$���_���d��S��%g��?�n�(*ӄ#���6M��:����[�=��D/b��,�V	�f�!͗lLьb�-�jFB��!�]ڑ�<yM=W���/��j�i��T�*�@,�	���u�Aa8�]n�s���!)���n��,?��'`¡��`��fVOwL½��e@�Ũ������J�����PzP���\ڗc�/�V3H~�R����$K%�g���I>ɚ��K����xpxǻ@�lMJG�.��r�u�D-�?͗��0a�:"�(�l�/�q'��}��#EUS���O��PIZ�gA!�<t��X�9���&��Z�'�&}6Ϡg�<Oy^�	�0�6�*H\ʀ�,,N������N�&�MM(��`���x83���"b96<�w�+���1'��Xr�R�I���8�k�,q,	2�	}����1��s=��~�,��UR����0찶���#�$e�6ʀ�O�:V��`��� ��W�Y������%>:!R��Kӡ	l��"Fr�]�Y��ɂ���R�k�x$G���[,�����8w��ݔ��A4M�t��rk:I�`5��j^���8�A�n�u��"2�RjXu���
v���=V�/�/dx�����>"� �8Q�0�����R�V��r���K�n�,��7#OM�@ӌ�qdQ=�Do��	��/��Z���EJ<2,ax��h�ҵ����{i�}��%��O:����fL
��s�l���u[m/�d>d9��}���P��(��Gw�@�W��;ؘ�dF�/ԌJ/7��k9D݀��W* �_X�Ʃ�L���?	W�uc۴�1�v���0S,�� ���Y ���g�l�tn�5��5țj\�����Eg�pcI�-"CWgo��^<:��*��e�x�� jׄ�y�}r�Q�u�춤��^����0�]��d��q��:3��r�20��1A�5�_9�B���1�z0 j�+~�t����g����ˋ�
���va����%�zL��P��!c~1��>��t?�PYi��Mʁ_%;���/"Sb��q���F�F	�I�o��G��
@ȯ����Z�1kpGi�;�ܨc����%cd\6=��d��h��
.�S�a��� k�A �a�$]SP�*襅-��*q��/� ^�"�7�*	�+�L.���f�lsY��`�mn3UQ)�5Hk�SQ%���i;}�����S;,PR�m���''��ƎFd��e��0l���F�@��Ȣ�@|���h��u<D������a����eE[�@Ii�ﰥK%Ú0��-�����e�s�̸昑~F���u-����0m܇71��+�n2ۯ�����C�#Z7�wW߱����׀�K/'b�~�GC�o���C4�y�,QVb�F�i
E�^ɳ��JC��"��j���9�Ʃ�0��d�2xW��S���W���05O�8�x�q�ܫ�e�_�[��,�O<	�|��Y��+���K��9��%'��8#��L��S��.�w�Um�!l"���]P8�5���:��YUޅZ���r�T_{��MI��8C�I�������Q�@�Ϭ{������ G�^}y(���ն��P�6F�)6�m�Xh����
�Q�RY�9{� �D��{i�+�]_v?M΃�4�ptw��H�~���p����/�qjl�GȩA-�M���gz{9}���1�$��Uͬ��n�Z5Z�����������S�`jӮ��>�+�l�~u��,�%�;q�^QZ �m�t���KQ��A�k�"7�ܣ�!r�#..��L>ӚFC��yf�&���V.��iɢ�ϼ�x��.U� �ވ��Q����p�ˤ^�Z�O���#��	��\K�-*o������;�/Q�l��@M�����צ� �af�Q��bJ
Ss_
a#���ߴlOTS��UW�<������8�%���Kh��tؚ���&�b�>��{%��/�D�G�*fH:Փ3�#V ���w"���ʅ�tQ��}�����c�{4c��0����<ј�0�r[��0g�]jaĥ�k�P<������~��y�9;�3�]
ĄRG(��O�T?����ݶZ��1�)I�L[ �PX�w�]DL�gxt�Y�/���n`�����6���|��U��O��=���s8��bU�;U��Am<�L�~Y_N�$k�j��d��������6�Y���7E��L9���5�ZeW�X�<n��=�DxyiGKčkт��g��ΉЬ�.��=[����K1�/`�E���#��ĩ:���76r�,�P�G��J�Μ�rYuC:~�� ד�bJ9��+s��x�5��T��;ۻ�Ԁۈ�`�`���U[����N�ng"� �Shb���dL��@3�������2�~�6�(�9R6X�|�a"���JI��n>7m=EoՍ�`eE�^��+�@f	woKJ~�V��@��v4Țُ�"�Dp�`� ��<���Vnp�8=Q�WοlvR#C4�a*\e3�����oMx�4�hx)���۽�"R{Yϥ:eu3B�d�=W��`��I��Ν�_�]}B�ۈSLt}��w�_|�)�6��w���>�ƥ�����[�b#ϑ�lĢq�9��R�?����@ӴĂ���+p���U1�,ҁh�Q�����w��'��X�8�t���v}$�R�%���D����3
7������G�I�ڋ�h����}���dH�n���=���YL
�*�_�Z�Ao���g�l#�v��JN-[HC�����C:M<-�� އ�#���^��V��A!=ݕ�]�z!�]��e����Q���ӄv@�_R؅����:D�B`��n~�gh���iq�EXO|w^`e���̻,z�1�q�-� 䆉K�N���br�u����p)>@쨒j�p@�8�n����/��b��t �PU�G�mN�!���$��JT<m�UK�h�����L�1��Jt/���x�����kP-��^�C	{��"�f!S�����Bu��|�� P�|e\��\�AT"���zj�,���I5ڠ�����'��2x�PF��*�&�N�� ��
au�cD�H�gO&�c<{$.�v�pw�e��z���&�{���o@�e�ldύ�!��dn��c7}��}Vrw���sk�a�ٞ�a�Kꤍh��#۳�$M�țr����1�+�}�ى����=E&1L�g�gŶG�.;}�2p���>t�=������X��rI�N�\���Ҟ*���"�W��o�W���-�	�x���_���`>�IwX�I 2��*���/<XſTWv�R?�^��B�?�m�kM��5!�xr�z���k�慼Ҋ�����I�Y�1a�'}k#�7��*aP�p1����d��7�qeǖ�Bo$�(4��-�=w��: �̕ @ �������]�cK�>�}R�u~^����M�n�\{
(6��q�P8P{��N���;�]��1ɍT��ַU@}\G&/�v�8�3t叮9"�h��@7M��3!<�~���ڽ�C�8	_弐$����g���c��(	�	�ĠY���C,4����M�4��4��|'��w3��F��=Q�yL®:�[miRSJi�1��+�i�z��+�:G8��u�x��AF�@��*2ª��ǌs���Sm��3����4h�Ў����3j��m�m�j"U'��xJ�8w&V��Y;�s� J�����Wm�����àʑV��q��<�C>�%ҳ3r�H����x��=�i�����J0��*)��Q��{����5m�,e �0r�{��"���H��SQ�H�Ӝxl:�[���B�$׆�`w�ߪkz�c7x�qS�o�gA���y�V��L��o�O�6�Cl}���s��v�;�No����%A��t,`���6jk��������~	y}*���1"Xrʣ#�^��rx~��5m��	U����B����6l�������0?��ٴ�#sESy?㝢j���������O��	�e�Q�rZt�����Qu�<�l]�š��f���a�6��Ԯ�8�ʨcb�����s�PY]����
��l=ybc��L��R*����ߞ�+8%ܻ�>�e��O#�%6�!C��Zߗ����4X��P?��פ��U������Ϡ;��m��}��Zg�8$���E�8п�=�0l����>}q<�w���!>S�6R%	ӷ�u�]=%\����	���Ņ�:�rٷ�-�݂o�&�T��!B����;(T�ㆥ����F�<�g�ұ�h	v�Ы��r�*�����o��l�	��.��c>��S���3����_��*��y�j�(#]��,�[��;��y}	�j���/::�P>Y;.Ҧ�8���~ �Em��4Mrn��2���`���>ihUY3��8�B"Q�	h�P^U09��J���>�y�˷�=Elp��OW��`^e1�;���`&�:�o_���9�ڹ��!��(�:�W�Sq��
�=,k+�t5��u*�1f�J�H���u��!e�����d��%�{��\Yh`�!q,D�I���-�l��r� �s�w��/��6�&����Fe��L''�Q'g�ń�ʿR!9i�67�	��]��N�#��l�y���ݝ�c��P�	sdP��~Ş)\�@��q3�*u�=��3z��F|�ڊ࣋sH�$Ɛ/�d)����N,�i��\�͟U%'��4�� �K�z�髅�Nn��()=���_�� ƭv��ö)�w\t:��,�ٿV������A���C��7x*�uc�nf�GH?i-�?�!������0{˨~���aQ��5���u���G��� _@?��H�~P��x���?��=Ba�̞��?bʢJʖְ]��DV��nM|`Nf8���V7n��nP�#��)�i��ևW���{�g|iM%
4s�W/V�X��8@��ӿ���ǔ�k<@��I7ksE���§�Ξ)��T��/ӿI��];�iuM��}bXX���VU K�q�mxW ���M �}���*�>�nJ��C�9��o�A�L$R�p��+�<�ޣthb�l�Mk~��tb���8�=Z�j2ƅJx�b
t0�~�Ճ�(3���
%4��V0E,�Ɵ�E�u�5.���o�HU��X�I��`�
�iv�\��=�Q�i�ʋ��g��f{�Η�/|թA����rL���-�>,!D��֠pi�E9�I� �m�HV6q&�~B���FF�c.�g5�s
tr!���f��J�{/m�wu�7W��%3B�O,&��G�+��E���0	l��g�?Y�w��X/�_����nZ���"T�.�FMg�zfo&**Ik��b�4\���
�{���^������ү����|F���gk:�ʳM)�ON��<]X5�%��
�'nk�7��v	H}����ǘ�O��1#h�X�BЦ�{r�LTʍ�81*�?l[����K�G8��B������d4�5�h楸c�Dj�ưf�f#s���͍Ʋ)�����w��G��<d�V�b�� "�\�R�3�ʁ��-X���Z�gX+&�	a%#Ȏ��Mb�ψ��K ���	K�-=@��Ag��Wz����W�����D��~�)����Ґϟٹ��qU���4el�e��y����恁��0�V,��3-P��M
� 	��t '�C2�I���L��e �T��vs�z���mY���_,�$�	��HS�a@��O��3�,�߫]Gm��b�������ߧ�"I �E�˥�}(B�>����nV���d�'!]R��bMg݌��f	�|F8��.(�����Y_�t���%.Hr�R^����'���B=����7�ċnʧ�E�<B���A�ǫN�����D���(��vU���jli�1) !p2��6P�_�h������wp/��$v���=�Q�j,T�,�-�ww'J����]I'T��w��wŲ�u'���dGW���y_QDe� t8��~!��}V��
l����j�Y�R���@c=ϛ�E_Abwh#�'��kk]��]��ֺ�cgҮ����c����0@�Ɯ��~�/�\t�M*�5*Gy�Lt]�.���<`�9�va�~t4�&�C�|��u��\���NP=	��/��O��^�׵�p�b\g�_�\�!t��{z�BW�U����28|�Tu�r<����{�����x8,�q���i::���&EU��Ab�G�$� j@�gl>ρt2퀦���r��o,�N3À:�V=������vq\	9�E�ԋ������?�X��f��ny���K4O@���Ǎ<�rK��uʫ9�ԩ�M7��qm5ݛ�\����g��\DE�����\��*I�)Kǥ�JCEYB��:�ɩn�$��.h�@� �\���%�QJ!�Oy��&v���c!Y��!�r���������݁�����x̗hb^�]�A�m�ࠖ�F��Hx�l�O� �,��d9LΖ�K��wd����}�Z�D#�R����3!��a�~��!���G���E���Ԃ1�5'a���x��%"?�L��2oBB?���D�i� |+f�1�ݳ��z��$�h�p�ZZ�C�f�u)�&�L6d�ّ%���[��|n�ʟ�����.��V�UBHʑ��꾐�q�����-�~j*�)t5��#T�ϔ� ԭJ�������+ ���s����n��x��a��v!ؔƃ�b˛H=��l�M���n,�uu���^�ĩX�-��LbQ��f��Ω�9#c#z������AVצ��a���M���ؼ�MÛ�� w?�V�����z��b��T�-ǍL\��0''@{�	cm��<S��6�w�\[��7"o���hz���hvJJ���_݆�Xp�`�݃O9�v9 g���j2�!V' ����{�A{�֚���.��SV�+�s��+i$�K�Q'氧8^EU ���yw(�*o���&L>!��6{����f-��G�0=%�Ͷs�A��g���Q�E���Ŋ� �p��`ׇ���)^}!$d�
�7�nlF٧l\WP��P��a�����ES���||�²��Y�N�]���.ؕ5�[�˻�p�&}�!�M �N��P���kaI�j;~��q7��K�<3!���a��'�	v�d�{���:< ����aW�mZ�R�Z��9 ���.��V��t*0�����s�jo��:�<&�ӱu��4� {��Ֆ��A�x��2�
��$mJ[N�)?~�*�aɳ��ُ�!���拡���Ofg����|KE�Q�L�qd�F�m�^�l)6}��q��+���DCQC�d�����j&{�o���'���p��w�x�KN������e�*�|�h���N��>�L1�0%�. .�m	�\��u��>$��;���R�<�4)����焍;+�x�pjp�a�gKC\o7�-؋o����"��h-?`��{�ʁ`1�~F#�g�
�ɟW]u�'mUVH ű�^1s�R���+RF���j��^�:$*�Q9�; L�1���Ȧ�V����C9eH<y;��dN_�(%�)��P�}���N}�~(H	,�`4!7I�Xg�[g� �0�P(UQP�z��ڂ^����$-9�*���?�xA�m�`f�Z��17{���n���0������D���z�~��4�K-3m��vZ��n��$��~<��-l@��CP,$8n��8c��05M��˃�����4��b��Hm ,�S���E,��75~��M�~*�hO��b�A3�iQ]���Ws����`���@�~�����m/x��ˊ �.��<4+��s��0F"ָ��u�p	�9\_�;^�,/�$*�����,D�肷�%j�;#D~a�M�i:�-��]�k���_��(���A_0D��h�Ғ�#�}�C�E���$w�T]%��=���o�]W?:||�A��@9U�����&O�m���Wp�JYK����*f���G��ə����?|���;����!Y�t�l���'�shά���.���d������c�����I�0��h��Ӏ=��:����o�d+Q&rs�dFfl<�����ߢj�R%Mߝ�9���7C�b������0�ƾY�X�et�eUL��ٴ�Ml�f���w�#��A�r_[d���o`�a/����ڛ +���e�K�dOW�wB���e���Gկ��7�`A����pP�w(2ڕ����Y�~S ~T69(����v8l��Lٰ~C�!�70����S�2�;9f������N��P��Q�����?BЊL��l�7��?^������E����$�t���|E�4����?��3.�uIW�`���ף8�]U�αڧ�i�`�)�Z��Aa2m�;q�lE��A��K��L#CI�	�?���_c�4^�ײ@�`��!�@o��@�N����+�)�SG���p��j6�T�1�J>�vV�����a� uL^_�i<���Nj[p�c�S���K=?�>�۹����Bf��t�����?_�CI�t���=t�k��6��^�uc��P�#'��qv�c���gK"�^�2��L��
ٻ�Í�;���	2��F�X$�{�c1c���b��f����^7E�&+�R/-PQD�����^��~$T��U,�	��'F�gC�߇��{h�"��
�@��,����S&�K��pv`۶-�MJ���U���T��I��܋eW�uF����6x�!�=ѝy)H�:��t����P� ���%y9�����!�&{�����=��ƕN?��d��~�n�01#dq{�:~wO ��I�v��f+G'iõ�K�8����J���\��uy���OH��*�)8�3��Ǻ%~(��&Jy�L�$��0�� �C .�#��z���������@�14p
�#C�/�n����gl7��v��N$���r���+��9�d���V�����%��,�ӂ>�HW(����J��f�qm_�p�x�+0�����vOXU{��o`R�$�(m��c�~or��W>�-�N*���)8���}�m�!P3pT���.���Hy��f�B��t ^��cjN�:��p
i"�|t���f�z[�FL�@��s��$?:�S?/�&��x*Y�E�� "`�J���,���u>�R*s����P
$n���7m����%Lm�����z]�l�3��<䷰��Z�i��Xri�i�{m﾿�'?�����������Z4Ix���X��;%�N��u���j�|��=�T�P|���d�V/��
/8k��/2���la���[䨥T��&	�ӛ��������Sg�3�&ɹ\�(��.�V,�J.�[�`S2%�y�^���db��/��D2��0+_�V�cu�Ћ�%J���.����@/��>G��7��1���PB�L�8�A�[T[A�J�A[�����ᮝ��&d��n����W)Z]i�ZF
}U�a�9}}x�g �V���z9쬣��E �5������S�^X2˅<3��[n���,r#AL�5��l�=�|�0�W~*\ʎ�����̗��2��r��ƈ0�X3<����op����m����3�N��d�/�4�]ԫ9%E����/,ׯ\M�IX���$��Ǧ���0�n��,S��i�D�{��U�p���!�js�d��譭�jǭ�~S�̤��j�%���G0�E~��yAo�b]�&�g4��� u+����-���l�ȳ���3E63�=��v����H୘&h�h����Px�b:�~M�$R5"���Z����K	�����G���M`��Sv�bG�(��5P8i����?���VY��a�|{���?"����+%��k<�Nk�ڄ��� X�/x�^]q�:�F_�"&��Cr
#�9�.)��D��2B1�u�l�Q��/���޿�$�a��mڿ���(g�4|:W�n�]ʩ@7��)���͑�Ț��E.�0K��>��s"&p���˅h�]|k���
�~-�ћF���+�u���Vw��	,�:���5������%��G����ρ��86��fί
Qǋ��9�s߉��\�X�,��eî]�rZ�D���}�T��t�K���Y�Jk�*sZT-"8�~e-�!K3���-�_=�P"n��\�����g��-� 5�l�7Yށ��5�V�f�$�[���;�Z�Q{�=wl��n�;
���1���wHn��Џ��L��&'��`�(�K��;r�����LTtX��.�_S�~\�[��q�gFCII>a�ݟ�71/R
_���sG�Fu-b������C
>��	;�x���d��BS�
���t��y2#H"���!����q#�w�ԩ�b��T�R!��O�_sc�	�{��9�M�Q-�z��O8t
��K��(�h]�1۴�6m�"t9U�����d����He�E��z�Zf�'��L�P|��C�gf��\}@�uz�1D���YBW��Yf�&[}骠�=z���8�o���c��N���I��Z��Jw�t+J��9C`��E�����>�K�\��Ԗ<�R�2R����: �}l�y$f�C}�-�����^��[�HL#Ѣ��T>|�u�-0t�@F�﵆��=P� ͈s��;�ٝ6��S���b��[��W(�攱�NE|�s2��C��$&Y �
�,�.��W��"��	�3 ?H�{�4ζᨋ�@&�<��O��C�k����:q�W%��VpR���>*��X���{����k٪&�B7h?��	����,�Ot�!��.[?"2D.I��nxr��Q���a�0��\Jq1�	��ʏio�	}V�mn����%��
SaV�*���v�s�9&aF��S�:{��ɋ�o��#߾�@���N���(���$�_�cw�P��蒙@ߴ�?������|�S����Ză�^�Se��l�����|K9���H�j(U�y_L�H��S�+!pg���qV�"#���u�F��#��3����o�e�����*�UP��Nlأ��:
���]6��)�<�>�8���X�ݮ�җ�|o&�k2���-vګE��dCXC��m��o�|�ålL����S����by�!�#�d�K�OE��{�qcџ;�Zմ,����i�Z-�#MsEή؂����|�z���M�3��w?2��[�^�ȷ�`u���F2�H2L��=�?X�H�>�.�����ї|�� ���W&V'MW+	�t �g�3�Kd�Ǽ+���S9d5�sŇӂS��s������Զ������8�{g�%A㠫��t��W��h��{,��z=�Iӊ�ޯ0�mL��2^����r1J$~��h�@;��\<��#.g��x�~��Mr\���PϞǝ�8�MjOs���=Է1���m�M5����-��wE.��t23j8t����.I�%p<���*����T�)�O;4^�Dd�2	��{�#1���@d�T$�C�[�E���G��v��aF��\�q���76��Z��\뺩�a�8��d���h��r$��k(�_���cl�lT�X[
�,:���ƥZm5�lyϓ�������c)@^���;Ă�D�\B}Wݵ���O��=}�O���!@���dp<��%>�i=Δؐ#�EB`v��:@H�^�\���MP�'���+VB}�g�Dz(�9��e{�0�e��͆�3�:(N��JG���y�S�|����>��"1i, i�A�(2p[8���L{\�P�UF�wE���ޒ��F\���A
��>�Ϋ���O�G�� �P�w����T��%�x�s�{�S"	טp>d���h�ia�P���v�A��&����t>���Z�/D��h��a"�����-�l�*v��K�J;����,{[,m�x��҃ð]�k �����"�os�#�`&����HI~x��``���n$�)m�2y4�I�n�.�U�:>;,Rv
��|���Ѷ�+�8��Lް��t��Z����c�����Xn��-��ߪ�qU���\�(�������A�E+��7�h;��8�u�L�����ɰt9s��G�sLM��R�j����S��H���a�Ь�O$3vw�ݹ��E-��]�#c�z$},9AOM:_3�ꉽ���t�5� 򧠦��&w�|=�LE'ww�d\���B�k� �y|c�����8vk7U����m���(�amW�h���QV���4-1�?����Bn4�B<V�C
�G�:����ڍ�L������]�ǉRR�Yg�+��h��cOk��c��~��ͭ5C&���a�S��/�@G�92�)<��ј��9�Q\m�)C|��+�#�R>����m���4�s4�C���q�M�Jh�P�{A ���V���aL�˓w�e���-5���B�1��R�e^�F��uh�('��Yi����u�X�~�6d�ʥ��Q��a�����X���%����Kק�v��`��B�4�':� ����
S;W5ň�IOA���O�&�n	��;��_OO%E*�S���Ӣ/���sEOr�m�d����@�lh��1�N[h-��;ڀ�3���>����^W�}¯4�8�(i�h�5A&c�P#w���рRu��������x�|!�b�HT\�\{��8dt�;E�P�����Uͣ�re���.l?k�c�F�*��_��F@��t�}Gg��4�� p�����I_��V��|����$�Ѳ9?"��x!�d��5����Pw6L���@E�p_t�Nu��zUN!��N����I6�2���+�_3>������>�F�Ӡ�W��T���6A��[_��XB���ص�Q���WDƀ�,�\�p�M~��3�
0s���#���~ܥ�XF��Y��Q攛��S0=i�>t��iB�n�����Q�S\�8E��KdG�.C�-��|��d�YW�V���� �5}F�_ �jj!����s��3�L~���5��S[�i>zu��qqJP�gN�h÷��!~ ��'-��r|����np��gA.:P�*���_/j��E��~�	 �����G����:�"Z�,�-j5h��n���ŮP`�u�����)��[�2�W��ֹ$8j�K�-�[%� #�u�ǵ�,��3�"�׽u��E���c�U�����-aU�mL�R�ce�L��Oւ�����-ֿ�􏹑];/�.n���ME��UíNX�;^���{���/��W8r����[���{���ɿVU)�|��Еr?LR��Q�	L/_2���M�yT�L����D����$�K�9K�{�9��M�sO?��S`�-h���R�U3D�&�k��zI����YSG<�>���@�9|+*>���-M�i��B�m�$�N��*B�o>��V�_*+�����@ F-I��s�V�P@8��r���
�w;�J��"�f���j'I�<I駟ֺ9�O�:��JL�t��&�S�g���T�̿��`!@Hz�ד�u��*Y]�%�1����h|>}�6%�W��H%O�DJ��b{~ejnI���5�Eo�}Ԁr\Y�d�_��nIe)3��C�՞�3���g*���S9�'
��o9]��nZ�I��r��︓��Y�i��O==���0r������	tC먴����v�#��׉g����`&3=�A�����1̩0���T��7���e�تk�u`"�6
�(�zg�$��g
�z�nARap����%��JM#��[j4�ֳq��c��?�Ae���N|�աG�U��ד�?�a"l+�~�8&�V� �� �Q1"��#�,�D����X��L��ίwنy\�ށ ���>�m�=�wh���²Ǽ�~�e'�Gu��9��ݟ��wUa����ة��\�Vp���Q����/�Q�찼��(�� �Ρ�+�#X�~���|,���Ss����Qϸ�<	�1�
�G����z��e1��	���=���fq�\���&�^�.7��Zf\jo僗���������2��%M���:��+ŏ �r�,���IӬ�%k=�}I�z�&fyhg�{<�Q��#��W�$�[��[���F���U����N?V,�˾qd�p�=-`F�i Z)�f_�ﲔ�\�?�\gl��ǝ������Gyg�L��VƜQ��:�Kl��i|��v{�]�B��.��\g��y9������!XƳ#��#�A������<���O
-�1��עh
��6D�|({$9@�B�<]�.���+�.1PU�nX��3v�%�����
|��4\T�P,}VS��C����[b]���[I���1İ�<A�ʸ=�PFn9<���}b�6�:$�-pvC!`���d����cТ�nκ��1q'�f���r���|C��z�;��9��-y�F�����E��bN荺ؽ|���>o�'��s�h�`�E�8�����	p<����5���TD;�S঩�����Gu&�m8���i'�>�C�#�z��wg8���|[����I�y�J��]#nTW��2�H];�9��s;mT�����N�Z�T�ɟ��𰭱�g����W�/�m� ��D5�*,��jdw��~�����d����'��v���G�m��^Kr�3����/ ѐO��i�3pF�+n��������W���[�/���p}��������\v�.b�ǌ�R1./P�wn�x�@3G������剅$8t�q�UUW�;�،���ER&�4P!�������7�]�6C&�h6�u�Ѡ�,Xw��/�?>h��&��8��hzK�;ݸ�����|��������OMg��3�a��rL����qJ��u��3�/M2�縵��br�EM�UϺ�:O�'��v�5��%|e�/(�kO&�9�G6���Z�Q�jER��в����t�t0F��~��b�(�ҝۄ�;!YSg�]C�۳J0ܞ�3h�B����;�@���i�:�}����C�:�r�hxM~�L ��4����z��/���TRvd3
�2���H�6���>7�Z��݀�s�����{�#;��,�N��[$�׃#�#Xb����Y�Q��C��	!� +J�p�M���iN�s�rW3��:��� f�|4�u����9����E��*��`���
��+>t&��|ԗ .�e�z��4���h�:�C'J��dޡ~:�ydٶ|Z��㠃\��m<��H���^BI�u$`�M���^U%���o$MJh�{�U�D��Sɽ��2�#PVG�z�¹����#C����ȷ]w�A#`�}E���4�b{�>�d�e�F`�=��wS8����0L��_�T[��"����Y�q_1J�0]��*��o���RҜ�_'�#�hc=�m��( �VD@yi��F����.�����{_f���?��?���<Sn��M)���ٓ���\=DF���*E����۝V|Q�K��K	��4��x6���M�+{I��T�� u��d=A�VS;^,�:p��d��a�h=�Ϝ-).���b
E=�ew��;��ۯ�B�B�}�C*pﱯ��G���kS����r ��3^svn���xI�/���C(iC�75*�)�\�?ӾE��[�ɵ ك�¥��yz.�y��lq��ϒ��8��|`9��m�ͬ��� ��
�1�Ð��q񝥣��v��տ�/��ʦ�<�_~_J�,�`����}������о�+��RA�K�=�����e��k/�8Bv�2����cL֠�6A-;�.�Ց� i�����(��Qp�1��2jX֣��Pc���-{ة
i����a,~�?���e�xe���=O�z�jm��O���8t�Z����8K)"SC��2*��O�Ii��F�a.�b�v��Ώ���x|� zd