��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�o��ȃ|s4�;�u�B �+=s��@��M����,0��@���%�H2��a�}�DD?~�%��n���q:�Y*��\�� Y.�lU�0-s�2$�g:M*)�<@H݃���V��ٕ(���ơFHxK��	kq.R���[%�/��%�|=�M�ŝ�
q�>�E*v��(R@���>���M�*��'��oҚ�Hf�,ݝ�ܚ]�������W�e���a�S����Y���=�5f%孰s��;�r���S��;ä.�u1��ԯ�C��XCI�:�ih�&St��t���1WC�������DFnaW�`�s�)]6�F{�g�{�=V:p�
3����@����	����ߠ��`��>����주�얗��D�@O�1`��E���ܱE�K;�JO�v�R(�fo=QP����0N^9�o��7�{�h`YWR}��rφ������\�F����m0�]��
&�R`p�6������]��	 ~��X�-���w8�@�:?<��$������*���X�PU��ZZ�U�������EaQ�Cg�5 �@��u/�%X�pcB,b��梍� sw���X?�yU���Y�_=N�,��`��'��J't��Sv��� F�.���^ AM3!�0S��%G�c��� ��n�n�Q�_9�$�.|�Z⇈k����3�V����&����=�
;-�(�ݪ�.��ԄP�_S4"�����sv�����\u�&��fD>�T�m�g��G��Wy��CفQ"k/M�l#av��^F?� |R9�L������5�Y6A3oJ�����N�땀��9�kln�8[��4���;_ɑ=����.�`GK�ݕ��W�/�,	^L[b��£Z)oP�qW�jR�SC(.���-l}��Dm�[g��
&�A�A��Py Ԑ�@]�-Ҫ�=)%Gi��t��▂�w������<o���!tp8�=�N,#!+�f�}�,��jٔ�q$��iə�Pb�qdB�͘��u�p�<s�pFR aՕk�l-[m� QL��}�mf
��]�fuo��&#!�?8����0z���ȰC
3�f!���F���f�<�&þ7^$�wɦ):X�B��hGB�-|g�^2�X~��[������Ty��\�3�{����߈]�U�S;�Jԩ�v0�O0���?�xR�9޻
�ϐHsk��^̚>��-�LG�9try*z>��,�X<�|i�]�9MvF��Zu�<zn�Hjz Ĺ\��y�@�9*o�~^�],���B���˨����)�����x��Ct�w���j�(�賉���?�gDu���Pwep<C�6V��Y��w`RtI� e���{�O(�NF�ȧף�f=�֡GdTB����M*��]�0zS'fm�X9ֿ>����>��ߎkh����6U�p���4�q
���!?q_{�%���4 wcP�1�Nh�������'#]����ѵ�L�v��.��}��'ݻ�-��1����P4i�_� }^�%�p
;�J��IQ�~6L�M&�6a���J�.�+�vh��U��d�sD���&�7[M��yD����o���3�s��p'G��(��i�I���!{�Mp֕t�]��k�quv�W����X��k�r����ψ5I�s(�A�k7��>5k�gb��wf��t"�F����d��x�S� �%.��OO�
�L�u��}%�s'��Q0������<�NBu�����M)^�UUUؔ�KL׵�њ]�ŵ�����Z�8WJ����s��B�B���24[��̩���P����3U0=mj�ѠP�o�DͯR�w0�|�>B"�v�iK+V�e%�}G)�:��O�dm�6hN��y?�T��Ɓ��"3���w&�jnL���>m:͑�������t�y)���8�Y�"��~|����=���t�s�C�=�/	�(�mF0����!`�c�o�5����g$�˜H�Ѽ���#EfP�}+�f�h�J�M����;����j����G��:R����^P��+�}-�m�ç0�*�u�d�K��J�ś`�#�L[7��͙?�e�kdn˕�lC�WoJ�+�pSd2(�⻨4��;HGP�Q�m�o~g�	������Y��8�`�S�dx�.�/]	ƎP�46�6�8�����
IY��m�?U7��bގ�R/��� �i]׬�!PTeJ�]r���Ц��h�֘��p}V6!}F�f�|��X�����p.7\���d8��a�C���ڄ p`3�`�4�m��J�aH/�.�� I�\�����nv������78bF%B�R�֐#7<�F���I�U�g���Vӱ\�or1�CT���<\����������.sőw�_�jN�4����C�|��R���5�|�6�F�X���M����#�f�:l���&�ZD�R4��!W�u�b2��6.jPxP:o��"uOz/�*���39_�e��+t��3�f��f����S{��A �v��?Ю����h�/7��45���1T�_�-��k&�$�R�Jc̶U���h{A�U��N����y7��I[���,��d�
#=�K����vD���]�LI�2)��`�l�l.A����kT�MC�D������"Et\�{�*R�����u{�/�v������O9.�̇(J��K����}�2LY����,��Vs;�U�Ďg�n�=�ivnx����ц�����-a�s�m5l�����D��Ăc���:�߀>qh�<��%�#��x���2��0��Q>-�{���9L�9�
��)�.�#~`�o0Ō���>H��6���r����8Q�f�RY�	�KU�Q)y�O�K���??UD���<�`��
2N7#-/3f�P�n|(]��W?x��������M�­N���ڃc��/�j{�t��v��%�$��B���j���j�w��1t�ʀ�ϭ�5�0?œ�ׯe\E���Y؝��U�|w�h��������V�k��]��_Y0�eZ�Z?sO߉��fn�${�S�p��5�}e�j����Em�)�e�'y���&t!��%)�Y�%B�) Z�ȹ6'lsQO��#%�a��Is�z|���by��k#�����1qWtSCM8�	w��T2k�v��6lU�8_��E* /t����j%�n5+ �iy�ɔ�Cj��w9��/�ڦ�� �L�3��p�KܤS�2�����E�x��<���P����:>( ��,�>�s�u@dI�N��zf��Mq�=�Q����A��S��4O��rK�q�\)N�i���#;�a� �7W��٩�)��p{e�cg������#����C��\�å�w�3�NVuEP�a�Rֽ|��S���|14gS{���H�є�?��&Cּ�(jgw�d���܏�5:	h�$K�����]�>�!+����:�b�O��,FzM�"����L�L��b��uܿ0�"V_�o��˧x`U��@���*�w�YS�Co-���Li����,Kb����������`g�јT�\4X|�z!��4R�BoV��C�u�)�Ziy���[��ų_˭N� -<tƞ0X9�󻕌���̤�d䷥잝�ƕ� Q�B��kA�@_�6����Qx�����U��l\�`γ} ��x�YP͋=�)���ko�+�/}�&o�-x~���W�r�V�|%|҆s��x��
�����iJ��K��(���ە��()�鏢=f#���˵����҈Zf?	���μ��j�( O̾�6�Cڢn�H�>��y}�$�3��A�^�!�[
���'C�͢��T%�b�0�<	{>�\���*���ǩ�U<t7a�k>
�ٞ���~|���$gԄU��ڪ�M'N�S�f#[��)=nR���3\��t��gq՜-��"�I�m_�l�#1��8W��`�> ��E��0�����ٞ����pU��w�G���4��.���*.�`F�-�>S�?�ζt<���
��)�;8Û�_qe�(��� 4r���	ܭB�s"H]j��w'�Ga>�6û9�pj���Y���)�L��z�ozm����I�*O�
|`t[�	���o/yy�+�^L+��f�����N�J4a+�wq�)��`�/v�F�8��m�D�yt���y�yu���?���'z��������X�g]eY-^�9�'}�rT�ڼ={���/�S~���U���4���(�N�<�͍��:��kB��Mw��b,��{ �E�4�a vseM���J���3����i���:۱���ژ��ۧ�jNp#��в���:�9�Q���|��pd�0�P�`���1�D��*��s�ԁ�^�uឡC�@�biRTώ/F�{��v֓!�w;m{ՈcM<c�l�g�r��3�	;؎*<u�ii�q����f ���@��p����2���5��	���lm -��L*7�G��"]gy����c��.�"#��2�n��sۋL��s7����˵&��:>V��1Jd�u�a[K
��H�f�~Ā��D�0>����u����+릥��������E�1y(�������6-�y�4��ˣ��L|0�P@��(/���hf��Z� ����c�{U!�ib4˺�bj��Ưĩ�#O�!���g��IY�*4��g�TB���L%���H�/�z\�٘�~})��3;�S����s�%8^��z�#m�0?�g�^bs��엔+��>Ĉe7~\ޥ�l�#,�/d��R�~�i	�}c�WŖ�Z'���$ MDB��0~��z�s!M���A	��S9L�^d�����Ba
7�Y��.px�+��kkJV*1��׶)y�VK������Қ~�[�c��[������������� nȒ�k����^��'fX��'�M����mr���H:c�$ gz�%��NFUoi���v)��Ȝ�Iڧ��V.f���prp�j�����LS��f3��q���e�~p7�[�� 	����2d	��[��� n;�dQ�q���Sϖ+�:aV�Hī�(��9�nڜ*�k�y b>q�dܢF{[,&��|���Zg�TB����\��~�����<�(�W�h?�j���W����L�q�J 棷��W�ڜ�X�5)����83��>�x��l��n�QHV�I a�F*e�{:.fWǓ�`$���=����XO_~s�i�1�9��!��-]!f=��&��=��a'�����Q!� �>���������~Ь?���zS>���� ���om�O�l�g�!�ރ�Zz>�U�";^�4S��Ґ���=��&���,O�u�
�-�wC�u��x���;�2R����!�$p��b��S��Ǌ��B�Br*\�ʨ�\k��8C���DXOF!~�<�1L]�/t����o��ed�D���,.�-�UA�DvdC�5��S���B�Mƹ���t����l��e�wY`��E"�@�F�f<c���PL�i1���~��M����g\#ZIk�B��%�h��ͬLso�ڸs�����͟��;�I�\�A�M�۞}�
�����j��6��b(���V��A���I��_��F��<?!5�x�㬺�y�/�m$����Hx�Ϣ�?tdb3NW�}�� 0Ex^תx���J�jO&k�҉�+?-C��H�t@}��@����1��$��i�փ��q�_����D<�����`Z(����N%V�<��ىꥩ�5�g�r���;�-��ƭ�1��.�Ϣ#��s�V�`��
�1�����´q��(ȸ�h��#�v�7��8�~C.��H��b��x���A�{�?��Ə���)��`ʄ��Q�kzҊȨqm5�Q��m���A�:�'~�Et��R�(�vQ�1��%�V+��ҽ�d�i�^����<���;�z�]��'�q�j��#J���1�VBa4�&� �I��������i��;p�X/�dMH��>ϖs�A��6e+�@*�]����d�R���(�,g�ld�f�6��rNF��[��z�Ɨ\~�̆�j�?��p0(PL��7���!�ϸVV���\%|�����2H�b��x�R�#�<�&�Q'���;�5K��Y��m+�V�����8(�s�[5E�	�V�34���2�g V W�N��t*O����8���*klɻЭ�&ZS�����=�_�L�]�#<��2^�-��o��t���.i�a��^��uO,�S��a���T�����������IS���!�A1��F��~��
��ɛμ��- e�� �3��h4�V�W�MP�(ώ)"c�r��e����"a�WK���?S������Y�� a3q3$&��^��g�}(����q0���������<�P�m������L��=��G��"5bSXF���N[��u����sZ��<I�`����25��!�Z��@0�����u���;�X�:kO	�%̆:����R����"�	���sJh��&V���Ω��oH��+��6�Z��2A�^F��o���{B��L�F��K�M|p�t7�K�%���P��ϋ�cM��v�:k�b<�>���ʚ��k��;�R%8�����y���{�y���"2+>nz]~a������?3�h��/Z_/��!�1-�iɈ���O�J3��H���)<�?�{?w)��������J�Q���.�֭/'�f���Gg�L<����$& 8OX8�0:�ф�# �Y۫�ni� !/��1?�����/z�lgl���
{G|�$�+����Ɇ�M�hn�A\0Fɱ�I�3���Ӑ�����J�{^
������.7�+��?�Tu���������	��B���T�9/���%���r�ՄTe\��mWԱ���� ��L:���ur��-g��b�δ� �yX�.��=%�	���+�#h�}�וdو͚�E'נ�<?�@��ka$��$ �F�C�c��L6�~��	����a�8,�G=�dމlkD�g��q& 	�rs �ʅ�ք4�;���j��J_L�~]O��b*>��f��P����A6am�Y�a�d���CaL�.F����n"�=�j?n�jҔ� �����Ɵ"�dR�fR&��#�i}ѽ�%�R�[�<�"��@��`C���8�u$�ԹLj�	���Wq�HI�<�q��2Q�e<R��?�$�<�)(&��.��L\����ֈ��_���$xtZ3T�9d]�a�O]+�&1V�:;���� �0��\��ϖ�"���+�b//)������2�L�MhT\;���
Ć�Ǯئ"y�������rͦ�h��T�lD��H��X������B�2l�s1P�Ё:�1��OC*�$%~`�����ἧp})�e��Ü���<�m+�-�4o�,��J� ����XQ+�u��8|�c�����Ng��)M6��S� Q��w��u~��8�gj�nk���M÷�{P��
0�>�dC@��A���Y<&-̩2��;DQ\�厓�d�k�e�F�W �{@��F���>]�QO��nu"��Q�Χ�PsM�����,����ѡ=L�d��������9l�Q,������C�>��;�7�j7���
�Ȧ�c䁇=��.�A��0�$~΢s�\��{�����W�$W�x��S�<rYUD&���������Ľ��t�����+�1֡2���yJ4s�n�J��RN�5�@L	r"7L7(�dfP����<���8sw_ºl�<���M�ptސ-��U�^ȂpzT%%� E�B�|�3|�z�z�o�W��\�څN�&�TM�ŭ���->����=�]��%mq�'3D���}���)!���k$�U@&��|�;��Ҷm;T~�䩜�m�H�*�L�k�Qe���0��K��0kny;.e�8�U���� ��g�0r��D�X�i=�pxĿ<�� ����j�ZHY��l1�;*7�\ �u[ӭ�f�҈��'[���:�����n�B����!���F�[	.a�:ϙ����������v�.<�(��J�RO�-(j�iK�W�V5�U�px��W�X�m�e��|	4�̮����1�E�������3��_�h��%C\<ס1�S��t!w[�&J��wO$��)��%<���M�հ��m��(B�����C�/3�~���pgeUC|�
K�����g�����D