��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟx�ɅT2n�x��p����Xh	H���9�Ҿ�z�1�� dT�h6��[I�����B�?Oq�_2�9Ӑ@�p���G:26�[�6T%,&'�#JeR�+񸊎2�Դ��E�Jc�������5N�{�����Jz����+�:��G˦�<�_�	�'��k�Ov-��5l��|~+��,�Z��r(?�! WD_����J���K���םcE4��%2���qb�B^���p�G�A�t�D�&<�aC�`$��v��&�W>J�4��q��r}�Rx����_����?��	2��@����K�P'a�g�LT2?��~�_��x&�'�>$"�&Ϫ���GǢ(�݆?Y��B�(�'��#��ֽd��~�U,�j��@�I�mY���^���� G��0׳�Z|�4�J�����y�c�f�����]�Ʀs@7�J�� G��MaV�����zv��N���ٮ�������=@$ F��qi���G��4䀞�+W'm�O�����_��b۹%�x�{�1
��Lφ�K,U�G).�4%��Y
nFr����� w�,.���5�U�aK�A�F����m��n���\�4O�.�������
��&-�l7�h	��]�o �2Þ���́d=�A�#u2o���hn2"/p���O��W�g�l3���دL�F=�s��!fˮ�r�C9d �n��%5�!b�RU�� �?O-$|�����9R~��_G4߷�k�I�ިiC�߄9D�"�E}L9NL�8߯�t��lf@�{���`��M�ہo(+`���(�؜Iz4k÷�'$�M#jGQb.~킺LY~�����B[Л����>�"����U��&_ύA�x�����|��<���T�5�7� �� �,��a����ȼ���Y>��&�a��������S%-oE��������iR�X"�Q��&J���m73�����-0ݝ@�.ʹi#c�ǀ��L�Ë`N`s���]��J��w�����/�˵���������6O�E��*�3�.ö$�g� KO��U�O��{V.�pY��Z�nÓ�OaB'l���G7,iD�\����SDd�\�-�I$d[�d.�h{�ڰ�a�;�xO�ݺ�������P�Ū��Sٷ �,�'!�eӻ��_�٬U�),'�)NL����F�tȵ��4���ꉪ��d��; ������ڡA��v���Rhɒ�4���X��v�i���Lk&Ӂ�a��ZVH	;jH��`=8UJ*���Gd޵�3��Sѵ]��[���P�y*~(��Bt�ւ"R\%�g!�ֺLJ����׌�� ۨ��鈭��o'a���Ck�u����˘��[�Vi��U��k�@�Xg!�G�!G�6 �lKdC�U����~�FTm���I���6�)}������"�Ҵݰ�N94�f�;I�vF�
���O��Y�U�xZ��{��d=��k�s�I�D�	*�8�nWW�F`�nSR�f�g\`�_ޓ����P:*�+�0bz'��N��uس�����!��X?I���0� ��}/��Wf�7e�31��up}��(m~�"��9�(���駤�Ae�inSp2�����j���"-y�׵�7J7���V���{"�gg���9e��t�V�
�j�|ms�)���)+����1�l7Ε�����X�dpz+���O>nHA�F��6��	���'���&2Jk�
&����3'�Ӎ>d37�1{��ah�7,�M�N���n�b�9`�V�����]\ht{���~S�^l/ "����%�A�@�,c�t{�.-ݺ%O�2�&"A<��S\5�\�<���6�~)pg����{/�x{���Ǘ���o|l�����z�-�98ĺ<w&��ÀV���N%7��Op�tE�B�~�h��N���dk��:���M����{Ug%��,E77�+��*�����>�7H�B`��TBh�@��������]����B�#��Z�⑓��|���o�>o�*-�H�ߢ�˱>3���!R�L�qJ{k{F=E�-���A-Sϔ�
n�8�����o���)���]3͕[3�3odwa��a
�� z "��+�w���14 -[�,�t!Bo�����<���"��1���oc�T�o7�D�x9�M�ih*\�����d�|�ȹ�x�����K�f����$)�p����) r�T���v�y��{�k���"Ei�	a_u�X��FI��ѵz%��N������Mz�MM=ml������R?��v����~���~�r]�Jj9���l4�+��$3�s���hu��Β���n'��B����X&���N�ӷ���M�