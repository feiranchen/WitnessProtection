��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]�������B%��;��ʽ��M	i"�7ݡH�jn�$
WYB�7B���](����HX#�X7&?2%���p���T�(1.�tp®'�/��?�yX�7�>z�LX�TT�L����̛���y�"eǩ�^b��[ (Dp4!;%�p~j�,2���͞U-r����+>�a֐C\���J����Yrjs�֛��#�){��VP}{b&Y(��Ov�ɨ�S�pL�k�*��5b��{fV}��
rv��#�)���\dM3A]�a�aON�c�E�����hV�����r� �uQ�Wc�H�>'*wtL�Q�_]���~`��,σϳ�?��`�!|P��@�J�lK���ے}�$>Is\3:�W��6a���F}	L����iK|��N�b��A��\��z �@mi�83iL�2-6�,��sT�tt���u��1�ﺘh=0M(���'7>�T��*"�M���Y�*��o�z^0Ҏ�w�_	��~*���^/_�,@2��eC�82ˮ���������:3�;��f��z斃�h8c	��J�����"�M�>xm�{��y�z�0��%�{�%s%)�h:�'hl��})����S���.Y�6 nO����s�����"nM(����D��J���&����Y,�,�7g��M��r-J����a�$��Qi29d�.p�?�@�ϯ�JW��*2v���+0������ȯZ����G�`���ӚB���YK]pn(�wX&��2e" *���~{�NJ�t�ߤ���y�ƈ��.�&y���r�e�EV��(Y˞9|�Uި���{|c�~�6N��﹋͚~�W�0�}����g�����uQ8i\Sf$ζ�
chb�栓u$�q�5R��R�Ϧ(�&��ϒvB�@����C�7;Қ���J�P�z��כF[V������Ѭ�+�#��yᖘ�,"|I�1�LC
rES�X��}�6�☪��O�q�郌U�ݴ�EEV��@(� �Gb�86���C;0�L&�Pf]�L?`*�2���^�Qx&�-�����J EgM9F� ��ƺwgǸA[Ͻ	R��.3��˛�k�h+~@kz����E&p���
��F!4��Ƙ��?����8Z�]�em����Ѕ��wK�lC���j/��4��a a�j/��
F4��tm���:�=�ʒ �dX�������K&� ��k�h�!�g���k`'�I�mb/�$�I�yR���)������*� ����O�ב�&�r��݈t��
PgM� �I�[�oK-X�MYMfT��c�x=�G�mt�x�4��A`
��o҉D	� �,u%�=����ӌ�4�����ǘ����0���3}W���g|�����UM*�ymM�kQ4}|��u�/O�.����AAHJ�c�6��"�PԒ�0�B%��ùS�3�V!���YP�>��A�޷[�+��nC���Å`�}ɽa�H�����6��B���$��!��u7��HCmy�V$&̓D��j����њ�ɺ�Tg��i���zzm^1���E�4��yg���~���;��5�A�.��ŀ���������6��d���^m'c?�$�<�z��I�5�l���(�x���KQNW4���<*�ޗ|[7'z(��xZa��	#N[
mBKHŧ�g/<�H�o�8����g�&�U[�4��])2^�&��N��P#�;3|i�:U���"5���&�{M��AL/��4ۤ<q���^���ʆB���r/^%�_�x���"9�_�L���N��S���|W��Rlam�n�S�`1��H�Dc-y&TuF��D��DG���T|�g`/$]���zf�4^����E�Q6���(-v�&#!6�	b��6%�:n���N�$����q����zE����/E����)�O~�k�����T5�ЩGN#9�����q�6���({�/5x�)О��2��)���x��
@}�O�* <���E��	-g��,@�}w�,��K����탰l���4V�]�-p��糍I�<�u�#�'B>�?r����*_] +�{��iĿ�lW�d&�� :w������-e�ϔ_����˚5�h�ˇ]��C���u��)I��ˎ��9T9&n��C$aƧ�"� c�v����P�-�5ݒ$&�p���P�+NT�^�>�̊�9w����s׊����?-���rS�:#2�~���ZQ��Ƞ��_Һ舐����0�w�Ç��X��)	n�^D�
-Z]����[n|n�o`�]��H��D�-��Ŷ�I��TuwK���/��^���Ю�&��2�diW�����ę���~N�4�/��m�U����L;.`�X%G0B:��C	��'a�60[Ṥ#�Ix�w)��@
��v8�	i�[��T�%�!��I���������ɂ7�(-��ࡓ
wu������K��)t��[�bV�D?ϊ�>�g�R6h��ӹ�I?m����7``W�.W8�&;�>5�u��|oCA��&��\�����|�¤��k�1��r�B�/�|�eu�U����&����u�j6@ �*�
rf��v�};'x�W���Js�bג�䝳S4hIޫ�\��&z�:�5���ͼtyUK�bx�Gc��O�s���3�¤<�����}��\w-SzC��]��g��+c���bԔ��P*i�1A��SE�U���KM����[��fݢ$��'���Q���:Wx�$��p�2L�Y�	-& ���`��J�C� d��%��T+�1��;��ɱ��h�ۇ5�Bm���G
]R�R0n�3�l�:�&����l�2�{&jX�}�j9����J��*�M�Ҿ�Bd���yy�GoS]{ۏ������ba�I��������I\��ޔ�+|�piXc#�1��� D����nv5[ǀ,�ًyC���ȫ�%�`G\&>C�ؤ���qs�n���0��7����߹پK�t���/_��nwF�J '��ؖ����[�����g{�X��E��#`mC���c�X�kp��JWI/�ʃd9n%w��א%�;�K�wP�0����r����4YPO㫞!����'�ק��7�p,Sm�.��@�)�]R����9].�����.� ��@�=�8�x��p�����YC�����u�/w�`��|��d+�#��z�RHNG�� )dʆ�h;�`���^4x�7��� ]"����;PM<��Z-�Iғ0�}�c�C(h8��d|����QXI����؏W���) ��@�\���dp
Ns�xZvF0��BF�{��Z;���u��0�I6O�'��nm�Oކnk�7N�Q�O(J;���� 'I�c��H�Tk������BOQ�3M���<'��J��
�r��eԚ�J���1���*�O�|���Le9B�J~�R��W���"��y�ڻ`�m"�'���=wxHd����K��9�癧7�FlA�d���E���N�7��h�,f[�\�D�J�o[�[��ڔ�+J���w�`�F�Xy�8��4�:m�}~4{��}����'h3��EjKF�n�6w	1팈�=