��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք�tb�R;i����	Q4��{�6�!�Y�x�p�)$��5��o&͐	�+����CCE���� �؝�ɒ垒���R2&w���B�w���ق�5�ʓt
�kqY�m��Iq�d�Rh,���AD�,Py��AA�Q��ƪn�^̘�� g��d�Yu&;{d׌��G���ortc����R�Gi������y��'0���S-V����Y�B��L�i�FF���ͳv
mE�����EFCW�)�Ս�1�y��4M�%�{Uk�0���p�ؾX�6��6��|��W�y�X:Wi��O�Q�����X/�����c�Nwͱ��%�c'=̆-����H�;<�<u`�K���̏�r��h���mֺ�]�V�/�ɰ`���/i@80��d�K�=-lү�8��~V	8�������3�|�N#�Vn���׿zK'q�[�*=�Eu�8]���tN�\��	����T\�M��>[Q����_�_Im+�=|#�ͷ�C��V�i����S�	��ş$(U�/H趙B�,Z����x#y�U���������	����=��K��_��FeFO���ͭ�¡H����֦C�b��b`bFf�9$yu�ӐM	E
�a�c{u��q��POzH���;ȲW��
+��#G:"�_����q�n�ZO{�fC݄��F�
���M��[��Y�R�5��L�d�&% �W#��9�(Q	��W^�e�#�<仾�<̷�]��P�ň��W�����P�a��� ��RM�w'���ǋ=��tx��c��/޴+�@��\�-?��M��o�RFD1|C"�c����@�C=*d 𭄿J���+&��M�Y���Z�z`�ji�X�s�_�N����������(|�R��` �=��0-d^*��K�]#@��+i��<���dvґ�K��D:�B.��<px�0B��\�[���v�0����8iR�{y�ȅ�9H�׃�W��^�M��� |��d�|F�J<ҟ���d5_�ى�7۬2�Iټ5{z\�ֺh.YY.��h]OG��R���u��+d�\�����H�A�&�Z���0P�ν{�ܫuQ������y��}�= ����k�T��D�^[�9���EBkУ��3N�jx�����1:�D��_��	 �4�QU�S��-	��;��,���
�8��&�����S���}R�('OLG���H�XޕFO��EB�j��ư~��Ưf��'RS�gw����.|�
o�iz�w�����u�~i��'�l�D��L���.���)}�/�]�m��Q;�����~��׍of��d���pC�CTY�_�d��he��t�I@-_T�%�ȿ�F�iSקF���O)g+����m��(W�/B�C[�f2���z2
����SA�{��a�0 !��S;� ���D�VC�<ͮ���n��iq_E�������I�M*�N/�8N֤�<��l��j+0B��70i�=]-��x`ӋLA����P����2�~ڊ9�D��7~�+��V\\m�=��QFgՀ��F+�`�����ϸ����uj1��,��Oc�̬�Ԑ� �c)��{7�l�[�d�?��N��ʰ�TN0�j(��N��#WW0q�����g��^j�D������7�Z�X}���N�O����b�6e��@�AȧJӝmz��*�зXj�3p�kgH,�l.����vIA�u+o4j`v�3�*M�q��	����Q��P��fq��W�II����VP����Jgj�|�2�O���e	��>E>F�`j1�͢^�8ܖlV�,LC���ޠ?��FUX� �c�������(Or��h3�^j�r�ꐿ�c�|Szd�j3-Ôl}K?\�����p�z/7G�_���j{ 6 q�gH}�֔.�ڜ}7��O���_���`�N��Gn�L����>N��D����	�8󧑫kG�����W-�*�G���n�L<e�,�
�����2��_��qū��r���V���b�;��t�9��d�����1b_Zu�ݮ#�4�4<�6��p��џ��Ά̞}�y��Jn�.v���Ѧ	v2�R��hX0*s�+!���z�E��U>#�0"��k\��b4��P9��I���s�p��q��*����%Ќ��� ���A =x�l-U�_�M~���>��<ѡ���t)F��^�7?�em�;�/H-Ԏ�۬9�Y!%[S�O>.���
������-�c�ə%,�f��2w��n�I�**�B�|��%��)ZN$C�� `��c�n��HM���up�Wɥ0���|�fl�]AڷuI�ȯ�z���Y�e�'a��GK8?.�t��)��8��~�j�����5�zK,��hԤ�]����������3F����!�e�����3g���K�K���Du�-���P�&v~�wD�Aj0�7����%�!�f���>}.� &L�����빢2�r�C�A.p��f��/���r�N�$յ�,7�#Rn��뻬�Qҷ���c#b�2e��l�[�E��(�U��؅���-�P��3^���|�R�[�ɕz	۸���T�JÔ����*߇�K�`����������'S|�_ꌩ�ʚ}4�0�k��^Q��8�pBt0�=X���X���n�`51}Uh���f�е�r��Ѳ<�^��b"�ri��rӈ�g��Y�f<�,�JM�A�P�s���B}��?�`eGUOI�c϶�V���n���c�F#N��yp#agNӨF2Y�Rܹ���bix��bX>`�q��y< ����X0�Y�!w��C�8�6 �ķ�U`���W�������Ub��ߞG͛�`�krV�ԗl)��j�Ơ�d���KJ1�;l��!&�K�ڒ��
3Vb��ۀ�e��4�Z/W�Z�!�q2#Dr΍�m:!�F��l�.��<�l��!���8O�v/�1J�i�5m�h��ɼ��ř������Ysu#oץ et�wm���r&����t<FƉ#�*u�
M	M��"m~\!:Zy��^p=�]Ê��(�-�.��6dT��	_0/��� b+�2E
�x���w�s���\���U@�95�I�'�X&]݅�B�cL���5����)L�C�g�B��C(G �w�i[-{xs,*��KJ`Qdv�Ԛ/�J�ޫd�"�@z�2�Zϕ`PWS?V����WPK���~�M��#����f��� 쯩b��뉶���#:N�Je��d΁�#�����T�=KRkP� 뼵����LB�b�'��"5��IYePu�̞Dm�w���t�&�1Mxƥ�)Cm��%�~W��ݘ�Φ1��3߮C�տ���$�7Vh/�׈n���E�s������ 򶲙��#fE �����3�.��uEO��X&�ԩ���Y�lTU����4�\�~��_ͥm�S�O$o�lS;��F�I�:���8��!x��6�_�A�����A�jZZ;�<h
����-w��ω=y�M3x�٥*����{$ژw�?&4U����qw/�t���s��*��@�����zO�%Y���t�H�E<ܪ`T�F|c��dj*�d��|���Rc4qO�Z�{I�6r"�8�w�Za3F��?��t4;dU�1��-���P����� �Y��,Y�|*�r��Y�6�؈7n���-� �&��,��Ff�PU�,���&���W�R[:	tS����6���<U�Ҽ��_����-���:TC|����:�\�o�)P�p��Zp���$]B ���9}c�^>[�7i9��f�2�H�s�:'�} 㒗:-��a���u�����sq>�����R'86g�iA��A�R�ˏ���D�\��>	�n�]��U�V� ��ko=33Z3�-�˺+:6Xe��w�^�.�=�1�����ko��4����3�lfm�~#��,�Z]�����~��!#�
�bc­#-�X�"|Om �o{q�?lⓜ���]&�U�Ө.y�����K0C"o�����S_�{����X5�-{�<E�˕r"ß���G�ps��v����2����\�o�9���-�/�3�����^��~W �}<�u>3%قXA����4��`d���s|E��XX��&z
5��jT��\�{�9r��6}�r�X��;ך�^(��'JXU��Q��F���g�7Xa6�4Yԟ�i�xW��s��V�fvo��p���K�X

��w�*�(���n������t*
Pwm~�����LE�9��/k�9�����K�T{�z����م���[���4<O8\Y�sN��$�ԩ��l8&KC�t#S�D��5�Iw��ɍ��K��C�p�͑��!����/�'g�8��U�}� I���S�Z�@a�jp�wnUIr�˗�p��8�?e�x��ӻ#��D�q`R�֟���v���ꐪ~T2��!��蓰*V���k7?��^Ȋ��~�P��E��X&}��?�@�Cح��bH�������o���m�uy���R��`�~�3F����tb���	cN>|ʲ��1s!|I��Q��ɫ<w��V�w��.���&:�)\ax[1�~J�t13����F��o�X3'*�0*2=��7O�nW~�a򏒥;$���4G��kJ�o5�Ӧ�\zV��N4L��]����<'_4��%!�#�ҨD��Y�E�2	�U�o��h_�x�U��f'9k�og���@[�Y�꠬��?�yD�Tbx��L�$�W-6t`�c ~oa��Z���#}+�7���h�\}��g*��@uNv��Z�gݶx���%D�W���\X�w�����b%UBC�	_���8�Ź$^��cٓ�X(.|�{�$��i��4� �����2�+�$P�]���9��J�%��A���ˍ�n@X+J$b�т5Ӆ�>OL�����g@�Cd|�����[ZA�F��QGM�!���H%�Rhd�b�@���KIqқ���r���T�wkĒ�0��趽�_=)E�yW��Wa�>���V{���	�M$�cs��P(a���%_�c�*�~)N ���F6֤_�!5�\��1z�߭IU�*w�oub�q3x��?��
����od���>w�J���ks�k�x~/��V��C�-e�sVGBO&�����F�*z	<"�����`td~��z�J�x�@���Xo{�L��$�
r�e��^"�2󗊿���+�iȜV��ʩ#-�IQI8\��oT �.m ݣ�',w��ߏ�y�m����T��<�^*�ES�O�\�;�Ee��˱qNX���	Io�nn�����p	.Bpnn�"_<}lY#uT�s0�c�v��W���+"-��� ��:_�iU�N^5���6�$���}�� ����*�t�r*�J�X�ij�F�H}ಫ����X����vp�Y����@sң�y�<9�%h��N�.� ���"�38��^���Ji��a�N�[&���:���40�u�6�ڎA�h�I��/+T�uQ���=P����Ӵſ׻Rh�l`�gWf�kX`~��n��rb�O�����_��9�T�}��z�^t�B��0�K~*1,���a�0�W dޒs����54���X����b��;:��
5�)2�BOIb�+ c������:c�V1礻�l]�"ݚ��-ʵ}�F&
���eE#5�1��n;�nO�M)��Y�����7�O=��77�@a�sM-�{�U� �n��������w��� Q�ڐ�?-���L�p2a�F�^7[Y`�#8NSulA{t=q<�Cǆ~�4X�v�>��rX
W��F�M� ବ3��V���=��P���G�˫Bk�o�i����<΍�x��3�|u	+�GPMR�"�� ��z9o������{;����[��D!����w43�j�~�
%��k���)����.��*���t�'�h�'�6�d��:�p����KY�i,��ҜW5�GM�ۙk��%S�6c�Һx"G���I�K��Tb����?� �.��4�,���tǊ'zHA������44��$��Y�F[�Fɕ_��v��-h�x���	qT�r���d�)��J��fD����LA�&M�f~�*�8�Gt��)��5T��S�s�6m<�|��:g��ېKWJc�l}n��ybS��]���ޭ��LT�+uH������|q�uOF�ӭC�	��#���^�4"�0]��V�:ծ�3|��G\+�}<"L�d�j��|G�OKA�}��`�(�$ߖZF�o����IS��� ����{Ƿ:�"z��?
����0Xv�f�!�rp,B�]w�5�v�_J�R��es�4ܥK �Ĳ��f�=�`T�A�
-�#y���A�@ZsS[������5���f0rG��C�6m��$�ڶ'^U����H���<�6���Kq5�.��o'GͷJ��V���A�
�󏶡��J�h�-�m���z����a���!��@�]���0�ѩ�����#W�,��=�Eh*8$��k���/Æ��X�Z�1���GG�7p&¼���u0_��H���b�a����B"<|R0g��Hy�b��Za0O�����U�'��F ��;�z�=���\[�� _$>@A[�~��H_l����0�K��@a�]� �в�������.:N��-�I\d���	��^���R��@a~x�[3���%��e&�.l���e�[��-�.�L>��@c߸3��r4K�b�U��&���U�ዩ߿V�f�'~���M�ďDܹ�0~���Ɩ����Sɿ���@$��gX��;�
�P��~3O��
�L��P��a �:�{�n�*6��6b�3-��^��{R����O
�M]1$�u�� E�w�|7�����k��ٯG9��k�ġX$�#�ykC���9V��޽�~I���_��%��V�U��`�%�Am��<t�?�&T`|��yN<���	~�����i�X�D�`뀓)����, �X>�))�x@?bbl�����B�sY�����-��1�Y���N�
�k�3�E�Rƫ������,������V�8a\�����qT�ke�/ג�<ͲO�V� ��+`����&~�?�k�S��ѝK*��g&�"�꬗��@�a�@�����b,�w�۲!�ߋ~�b���9��e�����'u�h �A��1`�i���-6AP��|���+�I��S�z�m7���mq��5�c����Ҷ?�i��jO�J���~Z;�
@t?nqR�S����}������S[�YR�����m�Y%��V��R��l�u&T���S�����:$׶�q�O�9ڮ��PjJ�00��	��ul���F�Ű�������]��t�+�z��+B���<Sa�
!ô[*ω��8\D�h��''%��aP����?���ސ=ˌZ2��y<��)�K��3)"d�1�ku��+��-��7�y����?�MR�����]gw�P�3~ʫ5G�	m��?��>�J�c%�v�	�}���'���NH���T:?3�.��sw�˖�ih�]�̈�+{R��<Hs���!����8#�|F&Zd��� C�)^�K��鏻�\s��r��bC���	6T�����(.s����ƩG����T�Wr�N�:,ޒ��6��^X�{x��P�ze���YG��b�t9/l���3�K=(�%��f�a1>�;�
��uƀ�K��%�3vv����9�K���UA�8���3��Gl$a�4�U��w�/T��Cx�'L�_ |)��ī�Ep���H}�B��`�7c�q`"v9a(�І�=Q���:��������%賖͔*���	��z�0�'Z>�/�z�2�����#��1��u�]���h#TcJ��6�q�0~��؉ـU�ĭ�+�^S��!�-���O�J��_�W�u�!��K����D�ɖ*q&l�>U���E��l��p�eV0��%���������r�LqO��ו��8��_7.n^����ٛ����i�d������.	�Y얥��^��J0��x�f�FMo�	���]�x����k�V���5d��bx����F�J�u���I�����}U���נ:uNI�gC���bK�K�����.��i��	&�)m��P��*�[ށ��2�U�L?���������w�{��� &�A��$���W��_�a����Ѷh1[z�w1��k�� ��z�7H�cO: ��i�~�+���ε+NUF��� ���֬�/(���-�/<#��PI2����菾��E#ʽI�2q֒7�N���)j�z�ü��\�l�	�O"׉D?�e�6O{��x����~����!�1^�1�>�'��t��^(ܲNh��o�F��Z}h"���c<���&ˋI��*��ג티�a9��9m(i|Vq63���g��阞s��F������0F?Bd[�A4"'>V���*};e��6"�v}���b�q)�3*/4g�|��,�����J�D{OlޛI)�C�j3�ed��/��uzn�̢h@���K،TĀ�/��i���?�2^"�`�~~�:���7?�P����屐�s�+��rz�,���4W$@}��E�X�_Q�7	�0k-$�D����4&Id@y ��*V>�Q��Ḳ�����1� -)��j:S��?\C��a
S����`8TZL��i=���q�bE�:�qң,�	)�#��e���z"3@Kz�=g���5�A)E�j�Ht�R7�*%>Ӈ��]�_�L�t&%�O?n�JQ3N:����ή��N	��/�j���9Y��pD)�>����
���m�>~�	>�њd3�ۺ�)	,^]�E(0G*Ø���ԁ�+�OG�lĜG��.[���/c��j	g|i"Η��At��܎=YI�uM{��(% �m�m�����t����e�+��(JfE+����3Bi3/w*���̓6�w��@�@�Ԅm@�χͤ��=�jJ@6�������N���k��C�Q��U�=��iʁ�5���5n��?0�>Kݎo.�(�W2M���rA��j����v��S=�Z���5.㍯��d�y-KG��Bl��!�Ȁ�_a�3�H�W�I`y��u0u22��،�/~|����t����e�%>d��=uzU&'1X�� efڍ��Dbg����<�6�,���	�7gxy�z�����*M�x��b�~�ەXn�\���|Ӌ�f��^ZyK0��E���<(~��%h�Hl�F��Yǻ���X !>�5�X���"�l�<O��F�5S;�~Wt����}g E��X��"�~�����>�4.� ���>>�8�ߓ���pdzJY��#�XraqX#�G�:�!}��F߉��gY�;�`�>�B 9�G�g��ٓm�oM�,�M��1�S�x%!�P��|��ETҫ��U�^k_J�*y��>\0Y�1�U3L��YE�E�����U���q������U#t���h��?š��`6�����  �Q�x/y*����[l]-\	c〃^~:�̎��	�,2�[\���~ ��
����[�X
O&ĉ�̴�����y~��e�;8h?:��!uU
�p�8Z�dݮ�����"T�q/�On�@�X���ۧ]�V��ĩ\:9�l��oR�ݍ��:F�^G�Z>�Z�J�Y�?#��>$�D��@|�<�-���K`�L�����C�_����ˢ�&$��l4۸�/��S�GY�/�5��Y!���M"?q;`�T�;u�0|z"H�!p���	��,��;���nnz���n�{�S�T�~K	�@�L�DSX�G�$k�oݶ�^��+�X�4�o�0�z�8kx�gMr���R����Gc�������ߋ�FW��fD)m;���;IF����uZ3��}v!�۰R�[��i�=�q'��:�"N.�~�������o���`*j�F�H���[݌O��g{�X��:/5cY;5YFG��l9����3#�Wmf��ЙGQ1|�����1��y6��xq��E���_�1B\8q�Z|t]W��2�dC��r�D��������v�$ZJB��aU0r��G����N��JZ)d�
����]�$�D_���zD�fN�Z���N c�䄙��Cޣl�'�1�2��|�{+�%DÙ6��Xx��\2��|�!m��Lu���^m�y���Z���zo�f�``����x�qhR�d��*������Se}�k�u���;�ZIHs�N;�����ฑ�"x̉���%Z��rH�p����J��N���^����9;b�#������k�%y'�0����tm�++n��� ��Ot�m�|y'���|�?����8�u|����7fe0V�_���I�t���T�G�W�=Î#+gwD$j0q���<`��n"�pB���Q��D(/��D�b�
o1!ey]�i�$���C%%?�H9]���yO��E�뢭��L�dH����B��{}i���ьȀ(��t@��0����s"��I�=e�B�8�h�Ʒ�a0p��D��.'�/�X�h��b9�!RC���h.ء��(����>�������ku��9F����}HcZ;�:���%�m� &�c�ߑ�70������]40�G��ה1����X��a�%	D�� Q�LXA��;�~�-�,�}����yя"��MUE�r<Fv�@�}2d�������-u
��O�LT
̺W�����r���ҹ۴B��@�t�S�4Mq���oh0�o���d3#C?*�e�9���1p�a�'X�֊Ӌ�A��#�^j��/������>��L�]-\�|�T�woI��LT�������I��ZO��̓]&H ؆�.�{�'�@G��:X�b��Jn�8%�aEf�A����)��HJ��:�|P��8-(. 0o8�A�u�ʪ�g�7����3	{��;�E	�E�`���%�tt���mRi��t���m� [��ݟ��Dm�@
�6O�=�Aѭ�15�	T7�[�m�>;4��c���i=a)c�i�Q0uL�$r��eQ�KyH��0�ڸ�!wpK�ߺ��N�Ptbw�l���;gh��5��w�p�z��S;�vx�;�)�)���^�)��"���跗H!<�b����Yb�~��$7mDН#�]nI�"{T"OD����#.�O����^�'����b
+&��l)��X �5p�4>+��BxH)sp��2'�ƸFF���^#�AՂ�`mя���Ҳ����F�EA]o��F�a�8��w�=a���{P�E>���� �2Ke�U�����7��$�������+'K�	W��]�J6\�Q�yM�,wjL�am�V(np^a5VRs�0	�����ћ�мo��@Y��;��ې��2�Q h�v��3A�)��9踠ؤ׺�}2��k=^&���<�� ��E�9�F}���'ʶ���'iI)�{�s�4E	�;�o���ؘ�L:x����F�mK�~��H��Pm��8���B�t��Q�3Q='>AK�d�_�͖��o���Q0q�s���� �����P�V�����w *ܱ�2�A��1�b����r֊��ͬ*����1 �6F��*��-u8�?���ꭳpJv�f�W�@��X
,��zZ�kS})���"���s�eͷ%����W	+H��ID�<��{Sp%����MӀ~�M廋M��Q� �I9�m��+�F���A��+3b�{�Ű�g~`���O)��@���k��f>�3:�k�-�~x[�������G~	Zq?�EW@M��
��& |H�X���uaJCȽB6q�O xYYdD�}�o%!��LUel�^�Z�7Q$v�"Z���^a���y�]^�C&�f)\x�h���'`�D��`����Ċ;�Ń��d}����2^�lp`	�jKPH��]�nwA�B�tZr�� 1�����>a}�x�Jl�r&�+!�0�dϖ3r�)~"�fX�{�4����#������7�� ���]�w�>4�8����..���/�ryQ��k5�"�G��X� s�̛�O\�7������ی�pa�������F��2���~}9#�*�ߌ4�s�3�P!�E���S�F���{a��狻��c_0LF�x��/���j<�t� ��ݓ��A/V�xpi*��i��B��v�B�gf�U�Z���Uн�� ��g{��{{U�1�E��U;���߉�S��É�a�ۓ��!6waͥ�}�׻׉Z��0y5��a�zC�w
i_�h��ڸw�~ �m��)��u��Z �`p,I��;{�5��������f-5�0KՇ��'(�������T}ge�~�9���ۥ�35�B�S��#j��t=�		��&�P�ۊ�a�X�g;&���� �@��߲A|X�d$���ۦ����������L�!,��;kتkR�'!EoF��H]�H�;oԀ/�B&>�x��X��k080� rS����+qV�g泒�&���)��01v����\aP��o�Ǟ9����$�Q����LHi��1�hp�-�n�'�~vG�G��m�#&�^�y�i�S�q��	�֓r���.��G�ʩ��&I�^�h��:�-�gVp���:�=�H��Q��.M}������W��u���/�1�é\�=�(9�P�њ�)�46�)�ɠ�+�T]R�M����3?�H�P/!��x\��gr@�����t��O�͊���p�˃�#�C�Z�E���ǫ�>�%�Ub��#k�R����Z�ә��
���u�-�h��k,��ѽۼ��G��H���~��evn����o+S2˷�Loe�.Rz��d o|�� Iڌ�����2���
�Tm�b�I��Ui?�1x��v���Q�.�Zd-�x,u�w}h)b��,%�.���ؓ� 0�l���!���o8�jQ�]ݓd:E�e��7�����W'd��kJJo)>ɣZ+����"���W�C��]���g�g��(��z��5�p��( d-��U*<���O��]y[�\����q�LeO�x��v�z���q-5��g�2��A�RĒe��i�1_EZY*�L4���� �1.��R�Vo���WV�LX��NQ ��ݩL�rL.NZC�'VV�O 1�ܷ����-a9v�MoɈ�u��\��3�D�2��H��W=��B�n>�j<:�K�;�/`dl��q�c�Z��@u�����.�ި~�o�pyL�Uln	���ɋ����v(Ծ/�����-zH+��Ҿ�U��9��N%ۧU��zE�9b�i����'�5�0�~z��p��|t7�.��"��N���W=������ s`�#q<6��\"K��n�#�(�w����gc�<��D�[H�)�4$�ɤU��[�{QrK� �	���mij��Y�����'ZrKnTĥK�,g�
W�,.H朞���0�YЛ�S��u��A�w����O��5��o�˪9U��ߛqd��\�<����^�B�'@�%�g~4si�m��p���^p!��o�
a��?�1@��Ӄ�v?u�=�O�w�_*p�.5�ָF F��:�s�ȟ��i1Gx&����VD�FE�Ų��a��6���v�.���z�$���ʍR�pMAɞ�UM;0��n,gb�{E[�?�l$�}M~������֊[���N�nEYw�K��9�#����{�'��7���w�p�{>�,�V���M铍V�#![K��QI���G�����dE���h�s�/4�*M'^��&���/��S-��G>H����O�fJ���6._���5V&T7#Y���|� �q0�r&��̱H����;r�b���*��4G�nU�]�i�'�����
#0ö%r��IV���4Z+"Z��qO*��p\��Qm�� �E1m~�!�c�T��+p%�̏��|����CRJ��vd?thO��?�yM�1�cF�F�f���2�	�DS�
���1��W|�'m����*��3_Ф���g���.:�b&\i�4:Z��A[�"�:��v�
)��M6O�-6�Z<6�5�
x�́� �z.�����r�Eu�3^1D�S���}
�'����9U����	%�3+��
�6��A�@�.���6`�dE�pס˞]�F:%|��.�M}��׬�^++H�l#��������:Ɲ�;_(�n��X5R>��������3bH9��+�V�+����?���I�2��0u�fC
]�&�;�# r��s/�����~&��(�5�X<+�E}��x���o�=>�����S*��I���F:��;�ͮbό�<�����^�u����V,,���_�$Z������)ZR��s�Jh劔����݃�(2��Q�be�)k?�0�PMHr��Q�dHD��P@D�ϰ9����c@e��h��k�Y 6$G�H���	4P���4�Od샖�H�lL1c��*���'#`=�__�B���
ы[��N\���Q���Bd�7��i�09����8(@i��94���	�X�(� N��|e��F}iA.�.���OJ6��^��D��)s�y������?��f'e�I��ke���>���'�"*�����&���%
:�I��#��d��E�ֺ�"�K�$'hC]�嚫�������i5�&T/�yv%�s�d:�����O�@�e=�(�ϗr��P�	��$-�q��+nѣdQN>�[8��*Z�C��yQl�w˺�(%kxH�7��A����腣,t(͔ʾ�㍊�,���;k:��!�^)�8�ixп���j�x!7�sŭLYL�IC(�����ݓh��9ܼFI�P�U�u_�k>a{+(~ ��&c�&Jh����P�	;�s[E]�`�s� ��"Oǘ�]�_e-4Z�\M���_�>�Ŧ��'�3 �PG1D4�٪� ������1Bō[���G�p&ث ^�����Zk���`���*lL��g�3P�����+̕4	����T~5jlP`k7�愋�仫n��\����¬�č��
�# O���ç�o�+��~�5ՎȈzgA)��&`����u�7b���`����6ָiHgp��kl0��a,��$4�ʄ�|�!.�̟�݅V��r��=l����1U�5>R���Pg��%qJ�yW������=@)_��M�E(#�ݲ�N �����9��02>�E����X�-��Yb�cI�~� �2�:߶*�`��dP���������\ǡ��/� q9���$.O�z'K`���٩n4�=�`A��ZO�1������$�.�(\{��P�h��&�I��R�V�v�1�k{o)	p�D3�ҭ��B���<��.6���MK�gq�!�"9�K,ˏ�_!��pOY���)����Q�u�a�"NZ���./���C5笸3kr���L �2kız}�n�sX6W4v�L��p��nX�t�PT��۟��"�lQ[��;~�րQ'�Ԟ����X�0�3�3l�D��Ŭ������QV�jvB�b�H/̸۳�X��������ʴ�{R�ٙD��a^��s����{b�J)+�6p(��@����m�	!F�>g�|2��a��r����L�S�"k�~��8�2��[�Y5QTi\��h��V�ھ&�`;�y�����k�����1`h��A�A{6ws&K7����:��*�a��X��{o ��v��u˥i�k���j�}�1�k����o��U���<�E��%�?3A�� ��kS�9U�W�83Pq(au�=�l�,䛂�囎���M�6����\��J��M�{�]��#c��m��4�AP��죆Z2��"]���L��Y�l[�U�m�ѭ�Uv�GA,Mz4|�A�o8Xh�\[X٪Ʀ����u���J|���h�AH���i�)�#�r�j�WT�F_DB��#ӊX�~^�6q7�/�}�򎊻��Nzl��f��q�����?�t4��8WMi�(rNAr�����2����w�ԣ&b���a���s}n(�y�	˝U�ߨr<��|���������9̲�?Rk B5h���O��0����A3�z��b^J���M�]O��"趇\�K1d��IN���1__zy�H���o�f*�\'��Rg�38�k��/Uk'۴f������Ǔm��6�¸N�~�7�����a낙�k�`H����YY�?�� w�.ꈉ���<۝��0�;f�X��w��#3'�\��v�5u�'����U��	]�N� ��}�otb�������2+�0#�4LK�y� ��rA����v�@?-�-�)d�����7����@�!���Pp��d�:��o�X�F�Q��2d���ڐ7�+B]�4�bV1�G�$��v�累4�]�;l��W�^fX��?�"�˟���\)�{/:}�����?9B7�s�3����E���n*�ةI��#�8M4V�����&*c$@ƻ�~oŇ�E����i/��+8��T���a �M��t���(�c#�� �Y3ŝHʃ�`�x�ܽe��u \��0�ÉS���S���e��U�sT��p�-.q�B�W��9^>��MT ��y������>��?�!U���-��U�{m��pb��N�lsS��`H2�}�C}O5�x���o�[�����q�h�y�9���U�`���W&�ʺS�sv���vYWH19.zc!;j��Oʦ�*4ӷdrb�jSr�ޟ���\�E�.T6��.3�L�	:qծAq2�Cl���9��x���'��qx�~���"���9�z��np�Dݳ���~����/ WTn!OD��x�ۭ��:�bY�Ŝ`������Qf�.x.5���eKO��1�p��o�:$r"�#���2(WW҃���`4�1>����X]J6��zU�2%�����Iuda����q���R{�1R�QH�h��L�[�����RMXkz1��{����[ ��m�T�7�� �(k�/���X�� �X��gfT9��8��$��p[��t!����W�m��}#EU�*��޴.X��b;hEg��P��W�,����АoG	^:ˉc��%t{a�J�VZ�� �B�'��eZ*!g�����v�l ������uқ��9K�#�_iϫ��L��Kq޳�꛻��n�k���c�>\<'-i�l�,�^º�ĥ<���Y`37���
CA @v�7�[����P�L�+!=����-\:�n}�/v�,k�{}؏�����v�����4i��YV�6��!2k�0C�f��L[>s���&uu=<�� j���M��\WG��[��U�R͙Р������c���D����Hկ�FMY4W��f^pk⊵5�M{D�k��a@�p،��� ��tR�x���8|��Uk�_�]d<`�����CE$�9�l���E��tS���f�ߵ��9Q�S�#���ɬ��/1f �9k�hJ(�*o �Q��&E5Z߲�ӭ�J'�"X� :`���%ˌb�/g�,�#�w�{������^�����2۟'��g���
hqxN&�����w�(G��1�[H�������?�
�;�k�ޝc�IP@MOw�Y$��9����4X�/븈b���L6��S�[H���������~S�%L���Ò$��R����x���i��M�v��~��c��%A��Z�fICj�Ͻm	ܨx��5�Qi�sP͵��٣�n�Y ���5d�YP�R���zx	E���h�� ф7�L��G͓�� ۜ0��ɰTІ�(i�5ᠼ�������(��9D����|uA��Vx���a���F�T�c�Ayq�����#Lzg��:u�>3J�����́wń+���Ga����_zσ�`y�ʷ`b��l���Y�"��7���N�iV�G��0a	r�M^t��kȘ [ޡ2�.a��Hv^)��2�M��.?g�C��Pj��@o�(�m
�UN�^4�@���sz|a3���ϰ�fKKy��4)���0[�4�K�� U<X�������m d�a��Z�N�"�­q��Z�И�_�O��j�V��(,��䄆/�"+�ȟ6�p^�̮gu�Dl�k�[����8�i��Dz넚ld�[��.L����~k��������lC���7�ܩ!��U>�,E��9I�2��Y�LϜ`����>ݵ;�2�o���֒!���������p�P>���WE��;^	�d��Wc� !�E"�K���ӣ]:������__4��s|d�����F���(�Ԉ*�{��R��;�Z@�{�Xj�%P�U�c�X�;e��q[l��]��=���ԑ8&���-�H���;A��)�R��䷠>/ň��ȵ�����1��?!��+�e�ԋQ�&���F�:_�m+�!r�Y�2��D��ծS���QTFl��,�v�r��s29:.1�b�:�;fw�/T��|���� KT�����D�J6V꠪�rGJ9�ǝ(B���\:p���#dҶ�,���ÚD���c�N�[3�J'*U_��[�'�qt�0fo�´�(����u9��Zo\��Rg�(Uv��[.�mGTʻ5C���i�`�b�F�y�͖1�����0�(���Y�HПڇ����5�`'o�����"���I�b�zj��3�eU��氈<[�dM�n����Sv=��	�Bg=
+����)J���=��b��b�m�.�wP�0����D�ܠ���7*Xq\:�L��vى�'�iI�v��0ѫh��m*�n�5}1	��{?�s��T�u��Y�ˣm,,#�;�"iI��݅�(S�\rYMޮ0.Z�ɴ�Hl�/AH��ΘcB{6ц���cO,FJ�"�;:���A�]�iR� (�����	3�����W����*X�,~����X����@<E�x�0LY��cզb�\���c�%\ ")����Ǻ�n;�`vڶ�%:PD?MYM1��G�j�����!�t\j�P��G}|�篴�l�.���˅ۧڵѲ
���#���X�gaU��C�i��Jep.�F+K���͛�1"N�J� �P�!,�k9�
��7j\i�g��"9s��+�Ȅ��gd>�w(�#�G������'N��m2}���+�'�۹%��d���?���gђM���q췔�z3�˛�������
�A�3�~��O+�"K�� aau.�u|T���C�rYU�d��1&�f�2wu�tm�c%)���}/�V�!zM��YppT���&`�M���/�$�J���wJ�z���,��1�jw�`���mZ厵3w���+-��X��٤�ʸY.�������74��>�h�r�n���R)��^�V�)F�F�4��<I���"��K��:�UӖ����ͱ~m�sb_��Г���b�pȖ"�Ό%x�k����iU�Ia�5���ӧo;湿���D0g#��:�'�y��ݐ��U�"�uO�k��FXzL#:�q��1��@Z����`1@�52Ob�#�D�i���;��6|4���V/�Q�ۂB3s|;����b=�F������=O�ɶ��-�]1X�r� ��8�B�W�R�bI�7�T�5mA���,=���X	��c�ǹ�3$e�W�`�
���*WWQ���Z�D@{�����̈́��=�~�/[x�=���;K	�5=Y��o_����HI���V��y�&����2j�+ �gb��E٫Os��?��"����luo���$�߉g$�	�	���[r$�:��ZF�8�A�$�^�����Xx��7��z�0�P�(!$�}�.*�T�86�\��<;F�(���xS�|{�h9I􆞞���j"�v����:�p_E����m(,]Z�W����z3����-��C�6b��v�F��)�&��m��	ð�i����^T`����edP�֣���U��fy7���T��R��f�Ӥ8��	����ڕ݀M%p��^|}]�5*�X�pm��BG�����|[gZ���,�yd�5��~��׳�8��k��\�j�h��}������p�Ég~�v"�÷Y�-��V�%%|���K�Y;��Ҟ,���K�[b�v?['��q�ă�F�I�5�`g�x��<���pI#��?����f��E�<���p���ycL�WŒ#�t½�	�>�1w���3���V��h�s�y�}�ٵ�:��P|�	�{y��{���\V��?6��}B�R>���e��?�C+Hi����]J����4�� ��/��Ɏx����G�T�IR�Z	�o�L�����B��^�����e��_&)�4!��i� d�e_�O *6G�k˩I���U+6I�4z�q�8p %�ɓ=��ŭ�շ����q �i�#Y���yd[���͑�ɭ0YD�5����XU��s��[9�<�y�m�L2��R�:����d�hC�f�L��l�g������d��c D�I���kd�T�r�����owwA21��,N*-A�(gx�(��W5�0m��&m��D��W!HA���A]��c��vC����:�l}��1��_ʱ6�|Z���/j��ه�;������&�T������P9��/�_�g��P�+�NV�bsg(�B�BL��?|�8��7�ye�&��x�ʙ�?���#Ҝ���d��$\ as�`�J�h�u%
Wc��i��3�M
�$�q���D��JA�H�'Α�!2�m8���迼l�a$D�`L�4;_#ۻ�P
&���de��8�5�UF�E��Z7J�{��kPc:�p`�u�Y0�.�wkA׻�6O����d��ĩ䞴��s]xn!ߜ��X:�[�	 b�h^�{F�p�Gr�;/�.E;�ۥ5$1��Xc e9NaM�.�Iz�&܏Õk�V�ZpZ�'���(8fu!��o�#��ٳ�����V,ؘ��YB1��K?2�p�����Y�:QD�TeN\�t���5`�������C�n��N��bIIIK�'0v�.�\�?7U��b���g��ww���8�˘�es�����Q���M&�QxW�j4k�w�����!��5�`�.��������h� L%S{�j�O�Z��B;\(��P�wH�U�l�,<A�3�7ae��ӿ8���z"~�T��Y#����:���b9��C����ky�L2���#/|-����»TB���GIw$�[+�I��6�$�̆@�� q��EU�Bo�Fc;�o4�IH���0]5�b"u&�^�~Yg���X� �RK�_��_ �>���:�}2`�3MB�ܖ_�/c�DT��F�Ƌ4kD 0��f*����+����U=/�Y5<&����?;U�>��ڮe^�˓�x�Q@����-���W2�n�ʏ��$B�>��}NZ�D�M���h�����j�}Ż�����°B	�oap7D"�>j;W	�ހ���,�,�C��~��r�:T����V���������$	R��T��й�:�z tc�[�~ jN:�����v` <�d\������ɦ�sݠ��̜�'G�b�/������������=L#��3}C�	��;>L̀1eԹ;�žh�1QLZ
}���p�WIW���jblfz�����4˾+����>���$�j@q�w �?�Y|0��{m��{Q{yCR=�_�Cg?D�l5��OQaU<�X<�g*�!�� ���$�'�g��*��=o��uy��M*�c�5j��F�*������Ϙ�n���0�/?��s[ܐ���Oұ6��JK��P	X^'��闖tH?.�Y�_��:y�"(4�S��<��*
ȗfm�����Czp����"a�E�L@���q|a�h>a�4} t�8X�ѹV%e�I�#�;�[X�X��{�՚Z�H.XZ����l̦"�ݼ�+�/Z����c-���#f��p�Þ"x�R&M�+Ag1�4����_Ǆ丧gO�yЬ��8$����A�Nb��S��o��<I�;2Y��ȣ��`�k:0CC$�F)�f���(�:����%�M�T�W�wi�ذK �?�~[���m!$H�l��O�n}=�nz�e�c��K��Մ��d{4AS���ï[���Uav��W�p��Z2�x#O�af�k�롿�q��_�;NB�H�xw���T�]w�@�����2c"6Q� R�#R���' ���z�k�V�H�H�&m�D!���y�_���w�Tֺ�����!E����[?Rc�rP���.�BJ�c~�]݋�i��4��)�����ο{b1Gi-G�*�>.x�y����DKeL��Q�
ey	g��6�1|#�>�~����J��'p���˛bt�_�0�H���w���טe��������+�7�	`��T�Fo�AcgS��؂I�x��o��L�+������Nu��:ۦ/0���
��$$U�u�w����)������JUL�UYCU��*��v�`>3�Lx�3�g_�R>}��Xsߡv���L�ex�'���P�;ꆉ�'`q���ڃ��7�(�!CF�_��*�R�1�Ϳ�(zJ��0qģ�RtgV ���g"?�Y�kC?ٴ0e����j�{�t��]��w��v�ck6(cU9���"�+�"[�'��o��(���w#F��u8�wF�W���E��˩��5}��o�*)�M6rC����g��A�cJ>t81�Ba]�	��$�DռKB����΅��TzZ�C��d�1��&t�,�dVݘ'Msr�G�`&���/<���HK���ƒ�ƻp����)�9߆��<�:�t1�c]�<@C��E�+��o�u�:�R��r	ѭ�D-�L� r�$�`��`V����"��'��25�Ḿ' s���;��X�=ȫ�!��=H�}j�]&0�?��~��.ࡲ���e<&1��L�:�H�1|��.�K�ۯ�5�rߩc��"�@����5�%�F������J&p9��JXQ��S�8�>�-�p��]-��`w�5��ޟ�Ku����4v7G1��	G�5I��oQ�N��y�aq�Cv2{c�����������|1�z��|8ӕ3���_��(~,�qO�-�J�К[5�I���%8%����_�$	ß�����D��4S���:L��]?��̰A�X%���>�@�̷�OL_a�@L�V���*4�Ű���W��e8F�f�
v"u�keXsk�c"g6 ғ.!���]�2
�D�\�zh+����׏b�V��+�O���z�W~��3��̱Ə�B��s��e�?Qsv\cn�қ2%�)f�P��\�"^�~eF�H۩)E\J��b}�/�g(�D~�ē�5�G���=��
�Y��G�D`R-"dm�Q�n��>uK2���o�Nn�l�a�7�ܙ�|(�@�d98j�Xd���r�<�����bQ~
�a���!^��#�
�d�r�f>ϖ+��͆��*5<�|�7��&qsVo)���:	��LD���1��U�`�yZ�Ƥ|�����\u-�J����� )��~�۫�6'C���t�����k�d�C�Oi� ���-5aO�\�#�H	p�J��S�k逺�XnL��-w�]�{iO�ơb������q"�ڤ�.���فif����<9�kq�*V��T�ȩY�͸Pf<��<���b�6�W��s�u'r�!EU���|P"���?��c�i�.��9�����z;c\[��\�F7����,Ko���a{!BlluS0�r��q��7�W���%Ln�V�%��MY1t��)�9���9$�C��F!�8O[ȣ�k�<Gݗɣ��@�\���Ⱥ�5��� ~�C�P[8�#���7�kb�� [ӌor���V��׻��3/3��W?��[���ﭽƳ!,Ad'3�$s��T�A�H6��N�(?D�	�Q������& Ǘ!�߻�OSL�5�$��?M���ΪKxbV7�[�~��vO��@d5�� x4/U��x��|j��@�klG�X2��ap���#3T p�<�>{U(�@� �A��惸 ̌�V	�!��	�[B�+��t�a���Y[d<\����ˇ�x��v���>��x�:&{HK��N]�I�vP�Օ�bM��/�=-��߸��̝B+�$[�� W8�&I����Ø�����t�Ox�k�r*��Oh�^��Y��Lyp���xf�]f����E�§���j��Z�+���w�h��*�N�z*�n{4�l�- �t��2�EZ��7�ZO��_$ �P�=��Ws�
w$�(�Hٜ?Vrcy�x��Ar1N#T�B����j�oR�"�ų���ޔ��1�����NY��P��������Ap��7�ը*�oA펷�n/���x�%QW��&*V��5fv"ȳ�����]��1`#�'��spj'
z�ݡ%����kH����?��!{��U��zRL�Oj��0����0�,�f�Oi�kOvs\�a7`�h��5��D�2+�L�t��b�d%�� ��.�:'���ϣ��z�o珶U[��\�6�z���n _?�C94�Tu���d�􋙺a�n^{�(= �?�n����^����r%��*n�wO���ǆDs���M �N���ΞZG�ݭoXe�=��C(qN�B�=H1Fvi�������)�>uoI]�<�,�j�mж?հ�W�����lgm����Ψ� �=߷^�n��2���DM��J�7?{�"�b:���,����Ѓǩ�eK���"�-�0 ��MER|-�uJ���Ne��aL�n�K˭!�s�ވf �W���������,�c���}}��W�Cv*�ޡ��w:C�muY�U���>��ԍ���(��`5K�q3US����j��VT�V?L�-�K�e�$_�0���Ԓƌ ѥ���^G��˒ q.B�F��Z���t~��A;�g��M6$�86�?3 �B�И���-�,Ľ��}�A􀟳���;�"�&�
L��C��&�>�U�څ�5����*V}�*
�4����B���
�yr3λ�3���`��ί���te��ҳ�o�����<� ��ф 	����Oʐ,�eN��b �|�j�) ��,ww���7���}�!�i�ail���u�o�	i<�t�"�}����#t/G'ң ]�J�,`eu =��?M���D�"ݦVy�!}=F-aNP�g(y��}L�t���p$���@�&��+��A��:5mzn�����7'7�~+�WtGņ��Ԇ^�xyo���.ܕ6%>�1��1*��y��)z����g�WF����T�T�q��=�Tc���^ ,��VBg�(�[�1�T�ڡNP����"C�@�;k�Ԋ���7� ��2 �F(�dS�MӨ�����;	����L�[C����A7k#�f%j+�-��f(��Ev�OV�H�	:y�&r����S���o�4�ӽ;,*�����"����g\i1���x��	��	5�$+d��p�5	�Hm���Z�|X�ϖV��m�i�)��@N{W�* B/�,t��A��6	���x-�>J��Y/�]~��"�6���i�xdo�:mP�vz�3�~�exQ���YW�$C�L�V�.�7���NI�d���{i�/�s�(W�ch
��f��M^h�?��$
Y��%ǣP;��Q�6׏VC�L �45D����rnY���� �bF�O�5�'�7��sq��I�b�ʕ0�ǈ^P&����4�ͰN���v���:�X����UȘ��~���>4i��0�ʞ�bs���\����Z��^RW��=���|�\D�M��o�[ɓכ��������y�����Ϊ�����j<Hx�[���n�a�s�J�V���iJ�����#��V����Ǆ���"?>�d{V�`��e�0[t�r�I!)#w�U���ڣ1~2�}	�y�r��s0���������S��%�ᦟ�v��cr8��UR�jiJ~W��P̍�"em�
n&�7��t���2��+�s%@m@�(U{�i�S���+l�g�^�I�N!��
��B��!�"�ԁJ�+�6��v�^�����y��L1�� ��;����|�|�Zp�"$��Z�d���#ƽ���%s��s�D,y����Z�tY �[����\woF7�y��_x��-��=-��S$N��6�>��p�E�R�=�谠�����*J6s|Cs}~�`꜑0���t��M�կHS�S��kK�"�ݖ�f�r��Ů�A �DZW��b�k.�i]��݁�x�q�aȾ�Xׅ>�x-�"��3z����������#�d��6�dZ�����젯������¾ԲB����m$���5	��|��q3�ho9uT��
�G>��˰�����O����ۓ�+����e�/��;[(�};��6��$���aG���&|� ��Cr13�R��b����a�2	�~�&G�7rȤ�^(�]�@�������o��4Ր|��;��sʨq"����&,�)\}j�o�L�O���R�!\a_4�h7����w&�N��s��LVx@���&��ɲ@7\Q�f�p�H�6�3].�K�+�����T>��$q�6>M��nK�G�y��U\���l�^�u��ެ0?�����RwlA�bЇ�:�p��������q/>q��Ⓧ�\��[���at�^2ҳ��轶(��u(��aAV�ɞ1�:�3���"?kWpj������<����"2��T;��q�:P�@��_}�ǳ̕x��zј�>
��=�6��Jc�#3�
�Iۑ{�{Oo4�Z��E����7�Q�P�Fi��n0�?u���dʥ����܇�p:*��E���gN��[x � ����e��S��/��^=t�N��s�2���g�)�.�/�	�2��w�C	'����N}GNU���  B��;���R���Vnv徯=��煖P�J� �/v%�0��0�,c�Se���G���ݮ�OW�>gs�v��ɰ�צ�z�[Xgj�Ä\E��7Ji��|���V��S��@f�1�s̈�֝`���+���3�;;�;ΊJ�14�ꀺˁK(��K��L��6�R�"�ol�JB�?מ ô�q��sq��5)�<Bf^�����xo��f#�/h�$�A��&�E'�Ut>�_�.������?G��є[j�oK����gI�^�菻�D���F����E�����eR����E�t�$H�5xB`���f��J�p)2m��B�@)���{�/�#*h�Y�:�]�۳%s)�~�"�T9s��:�H�N �r�$�����A]#�Ͳ)Z/��4~[!�!k��'�O�߱������Z4�q��y����<�V�_+�`�����
�q
���ѵ4cN�m1�[���MH@��^v[%�x�y�;��kF�u��:�<5��OK_N����3 (����W�C�9���;[��9>�H��BeRRG��8�:�']ݤ|r�P�n�g���I�:=+��sOJJ��
M�t��	��L���#*i\�e!r�-7�HVI)yaxh���_��?�CS� ⧋&D]� �5"��<~�'��w_X*Ѹ��[n�,)�#��(̖ɯe벱P>d:F�a������Jв]�����|����?l���$��J�G� \JчÓ�$���bq��ڬt���i`�������7�z1/��AL	[E!�Λ�K�7�s^}q ^b���(d����ܬ@�C�<�������J�h��N^j3a^���#��~3D�B��5f����Wԛ��Z;Y��_�<��{�#{J?���ܩ+K=���2��%�O�J|C�<��>ւ�e���x�� F �"�hMv��j���	<��U=�ڛ����Le/�Jn�J��ũn�򉸫�~O�0u�����m�ak>V[�)��<��"����Tc�:���>��'@�]�_���[��$�Iͪ� ��X�	.=��W�
t��n"/� ��q#��\T/��Qj� }��z��qpY���G��P�!�mg�P���|�S.����B�:,��y�ݥg��c�����Xa���w ���?\}֝~7��E�r����a��a�l�T]0FLW�����_���]͔Җ�T�=61%�h�B���w��,��(`Yɇxh�T���i��Q��*ɰ����d��?�{s-�/�$ݠw�4{�v�{�h���p�|���@v��^��M�2���*�cd��ް�T~�|�NWÛu��dD��_�:�W.����A�� �K50�*�C��'�D�4�
��0@dGT�"V�N{��ʶ~�H�X���h��?�ؤ��ut/�M	 ݔ�d��Rc"�B�ʅ���]�$Zx���r���T�	�i�5�vK��Z����H�7�Z��S�.ގ2���,ĉ�]�4��2q	H��C ��M�ݧ<puB�2qⶾ��T���mH)w|�v�����Ga�A.�-�%�������#\�!��[%� ��8~;�sH�e�r�⛻AEj^��d��yI��S�2��H�JV؊.�nc�65�K��
��tkEJ�h�@=1�O��s7V-t��tߗwt����I{��؁Ke�����C�����nG5��O!hA_���R���T���������^IN��7�s�l�aO� V$l"�1��	�$e��;�5q,ryD��4΄�e�������|�5Iv�+H�1��v�����dk��.�z�����o��Fe8{��&�6��d����u�q%Mzn�� �IE����d�J�-3�;������G�~�sP-O������˫��ӌ T���P< a�κs:3��J|�@���N�Թuȴz"W��Q3p�8�S����t;('n���aϊ?
�=������S[�u��	[wנ�chO]�X3�M�о�ԥ�4� �!�ܡ�%lJ���'O�mYl,;�Y�r �_oL������^օn�`�����S��� ���*<��t!�S~��nQ������٤��D�ͥ�a�1t�Eq�m�ʔ2	�h��o-�7���L�z���v���la��j���{"�0N6�7|��V���OH�X
����d�W��q�~����Ԑ�W֥���E�ŉ'Rȶ��站?��_/x����Ҕ�j([�29c-iB��6�%�UF�n.p�|���f���}[�8Xm}%m�~n��ٯ�S���O��"˭�b߆3�J���"��nے5�Ypꠊ�Ų >'E�V��쳎��w�!��*]�����\FX�+�ˮ��	]i����ڣh���^iOj?_���ń+�H3ђ� !���J�ȉ"�=��!�������bdkA(�e��M�E,o\��oW���o�����'�f�*�6���TZ��#�'!�W�xJ�0��H���F�7���.���.F"�i
�L�bk�S3ۭV��`7����Z��)�.Oә=�4��U>tg�g��^��-A,%T�_9Ǖg<��ږ�F^\�@2(`�%�*)-����~X��njM�`�i[v�S@�U��>� ��7B��م܇�>�[{?=bB��E���Uq���T�eT'C�G�D#�����Fߙ�O�bF^���� �\Fd�⛸�z���e�<YƈD��[�{���D1@�f�.p2��h�Za�_��Z>��j�_��| �*җBčB����2NK�u`iD����.�%_.w씺;�U�������A���KP����[�DE{�a��D�}E[d���ݥO�U��
�q��v�����u�AD�c)F�-Z*���Q��|в�o�����Z�����H�nR`�A��W�ǳ�[��,�B��!M�_�6�B/@�LGW�&��x�-b%�!�H�h�y�W��j8���tS���"&7�)߲дZ$�B̥$n�����JʂJU}��������A�F/������ӛuT����-Y~��o�g��^u*�i�@��)ъH\��Nb�����k8�A0����e)�S$oNi�������yo�X\���������D��d���Ě�m����`�0}����x�v��C�M/�z���[�{���o��1%�v��3�&w*��B�#�$��v��!�?=��m��ڟM'���D�a!S����=Q��obQʹ�^a��؂��e�svH�ɇ1����B�T�CwG��&�%�4&�˒��x����Z����q����צ�.�B��	@nE�so!�a�ZԬrҸ�M8�d�c�����=,z�-��|��ŅrC,)V�0O�Q������&��d�j9�]�A�)���P��Q���X�8y>�W�%��_���cs-���ш��\Q�͞��TՋڷ�1�3o��0C��m+��B䖒���=��b�8C�Y�r�{��~�'��$���."�QW;�kv}J[٘�]���U��G�At/|�����嗟�21���=�e�ȹ�E1��.7�q�4En�+������*ܱ��Է��f�,%&$�{�9@�A���.����`c(	���k�s���_�Yc�$Ѹ=N�)J��^���șE3��Q��W�
�\!�������|�!qH?ش%�$(,��G "!�G��!�P�%���'����3��Q4�p`�[����r?���>:J5���j{ ғA6��5�� ���1���С3�dX\�w�ͥy�Evv��tb���ɂ|D�|F��RpJ�;��uNDgI�޺*��vq��>;�|�q���("ݢ�w��<�p�P�s�S�m)�h��|��3��RMN�E}ET��7d�p�!�rO"'>������y�l1��ٍ��C��	F�u���ʳc��Zl����A��4�^���������]�0�g���ɕ�7mD�ĺ=L�����@>�~��8��N�m�"�����֘v�X�]3�[�G:�:�jm�Ռ�|�8A���b��9���w�3�:3�7��P��7>�5,��4'��R���&oW��B��9�V:��S�Ӽ�~��g,:�d82�}A?w��ă��8�}������ƥMm#�P��Wu��Q-��Sm:�(Bf,ia���:���_'k�Y�~�61�Ô�o���֋q�"I�_vs����e�ߒ�%u3^��\���!V��jѡ��L��Q����<R"f�ʺ�H�AҥBb�B3�i�>c���Χ��|o�4��bg�y�H�"�^6,���f�t��J��B�y� �Z�%Hl;��̢��rR!�G����ʇeR�� ������k~|:��e�t~lE��K$�m8��Jh�"��+�����+C��Q�[2L�1�Ę�4EF 4��%w��	���U>zKuO�|u;_q��6�#�v��D�����l��dÈ�W���L}`��9�ʷ	�!���r�e7=�]�2;�ك�-���8��{�/����+�13(�Yz�@}Z����G������ĨOM���þ�N��d��`����	�m]�&N�Btp��_;doZ��n���8f8�2x7�$�ư����FQ�!��d�#������?��{��}4v$��s��b���Ә�� ��_"�������a!Q���YJɣ�n�����v�PO�h�w�W�̆��ʟ�:S��w��4'3m!�?�<|1�T'��p�f�{�dՠXO^X��S�Wm�����엌1�A�c-�kWN��8�׭vd�Jq,&'5���yv7�)�i�,���V��'��aa(��qpX2�aY�	y��J�p��ocy y��?i��pr��?�����l�j�Io�)�N��6��8r{+��+2�E-��#<F���#�K�`��P�0˦�@|4�]?� x�B�� �H�܌�����PGQ+��Оy4��A�j��(��L߄ ��Q0a�@:B���A�<�bB���U��f���p(���EI6)�!. �g,����@�����Wz֐��V��g�9�G�G��۬Cܺ�v�E��giE���,��������Ci�E�±��5��'ɔT&�8IQ�C蔨�NtW��e�h��S*��������ɮ�u�m[�u��~��&N��8�%`k����G1�"�GP" ����|$Pe�ҹ����Ŀ|��~+V�e��~ɐ����6?��a��ص��(|�	?���L�gB8�dfɆ�;��.�Włt�az�b 'm?�:*%���]01��)�d��c3}���j�3����R�Ҡ��]�ge0F�p�>:u9��%�r��3�)`5�{��\b�,5$�yH�S�.Z���=d�*�lں�,G�xm!0��G�Q��Nh��ͱ������w�B�X]�g@���Ŷ�'����W�o �M*�;�s���Y�"�_�W�?_H�))��D#�2GLD���?Hc�+ָ
}�v̓EY�/��є�7�s���sn�2�4�|rH�y�M�{��=�p�	�Ta��|re�X/��&�6��^w���j��3�E��~�:� K9�/�=�!LM���K�(�ϵ,��
���֭l#��\L�;�.z@�(+�:�F�����1U��R��j�=E��u*4GՑ�%��"�=�%�����j��xL�0X��_G2h�d5\�7�ap-bG�)}���	;�l�mă�[�.�89/�6lzo��L[�8���p7G�f���ӫ�MUkD�f;��=��u&?S��D/2��O�%B ����ͥ~���ֿ��� �g~���}���߁�gz���G�MZL?�n�)�O��/�a�Q��B� ������Ù�O��Z&�e����S����W�!�ҥǴ�J�nM)�/u�̚(נ��nct���qr�i{��͍Q���޼���Q��+r�d(��j��8h�n�X���p�t���7�H�^m4��RI���Т^-ZW����2�i���G��H������#�����!+"Y@�D���f�R��f8��Z��YE�5=Q��iN���k�V�k���S�| �ۣ@m��k�x���Q�rx|��'Y�������t\����M��E�#,�r��i�VG�r���8���溕 1�?=�2�K~�V�ՙ�����̕�tƗ*�/�Ĺt.�`!��C��ɔ�Xڸ=9~��+�J@bB�Aĺ#bLɿwH�_@��phʢCr�� kObaJX�ͼ���c���(�mZS峐�4���^�Ak��i)��_��C ��?��/��"�I>H˞E���Dx�NU>�n)$���nOV*0@��Ц��j��I"�����sa�5�l|p�<��D~��yg�w����$p�m�����jw�~N��X�������n�Mf�f�Y5~��ޅ3�����>:���iaԥ�[J����3��w^�!KsL�ap�1�����B�"̸����5w1@�߰� �\9��0i'N�f7���1��*��I9P�)Bg�ЁY�|<��4W�x���S�H�y�{-�^}_~��n�NN�¬q!,��r��ŷݓ{d4^k%E-��^&����}��y	�~��/�����Ǆ�.���D��"��rU���.jP�}��0����+Z��T�nH�a�������钛�U��r�r̈́�kas�X�)���Y�й��wi�@)���+�3H��@��n$=��k�vW�:ubb�5���Oڄ��I���O�'o �T%�m���C���x�>)��_����M��-���o�qvJ�!�h�`{��Ԃ�����7~�NHv3룏� t��YH��0����%πJ)ظ%�n��h����e,�)��dj��E�Ns#~� 
~���:�>=!�ߍ��9�!w �'Ol� -"��V����LH��?�q��X<�1#�@�__t>�>� s;�֨V8��K��";Nd�I�>���)����l��!u�:��$u��j�0���8\�C�ڸL��1M�wW(�o�1
��+���[ w?uq=�.�'���i��9�I��L,h�%���98X����C�}w~K��A�A������L��C��,��x�O�e�U��H��`ӝɢ|�Y�T�3UbI���d�����Iil��������a��<��i׶�bj:���PS�m��+�1r8��ͻ�+�"P�������:�b�� ��L`�3���WR��˨Y+�(���K��Q| ���(J۠�f�Kz#���1��;��ߠ1�����F������4���wiP.S�k����s��C���J<;r3���>�VN��� ��[�f#�&�?f�H�n�W�����:��"��zo�����Hԇ��y"L��ʹqQ|�[ɴ���CV�#ɕ��(SM�k�860�kWF���V�(NB�Y->Tq�|�t�Y�Tuu�%�IG���Wi��A@ӅzdL����lF�&Z
ZqW�Z���8voM]5�}&sX�IC6���n6�ʑ�Xe�@T���}�������"}��Ď/J������ci!��G]��B\�^�6v4g�Խ#�[�'��7o�Nꋪ�C6� ������A���@��Ār�;�W
��wZ]{p����'��J�>��DZ�s�������f���-gJ�������n������X)�J՛����[���QR�5[�׶�u�4���d2V/����� �/H�g�͗]f�"��Q70��T;���&��f�9%7p�L��B����J��=ѫ�V��2�D�(���4)�2��MH��#�c%6̋`�{�&�]!2B�1�Q!�S���h<	�f_�xRT}o�α���X)�vi;���6k����{.���,�����t"�L�'���b<��W��d7=�~�D� =l3�z�uK���s�$�#�[��;��I�˽+�������>�OE�οq����T�[�4�ʝ`��5�|����)����*݉�F[�dUvW�ê��B�-e�Jޭ��g�dm�.5��0��X;�1�o�m���+��.5���Dۚ9����X��b1 ���s�H��#��uJ�D��sZ_	�
B9#�LTFmf�x�
$A,̏Z�P�r n��^=T�/��]ĥ?��=]�����'S�CS�
O��#���C()vD��@{o�lm�Q�!�7��C	C���g+�ZL|���^�hd�ٙIE|:����Bk��_����������#���@�%b�56M�A9Y]�(�ПbI�&H������o�ʌt���$�
`�T �d^O�tVӝ���AH�ՠ1��GG��,>ݪ�-TXA�G�?��ę���
���4���LnEL�}]�0����V?�Ç�M�X��>�3Yb.���[��ݚ��p}7&k��mc&�."��U ev��[L�CA��#��\$�i*�m�:�lN�����349n�W�-�9�JO)�S��'�RϲhVw�Bp�ۄ!,�.�D�I��]e�d����!)32=�G�n��*�C��!��Hig�x�� ;7�(�/n�G\:\���K�3`t>=���S'���������_��5���.MM�%ES�\K^�E.�o�ɼ�O$	[���2O�OmH*يZ�ܳ��y:g{O�ć1ѩ?�؀��Aj�9�\ú[g�q�W�Y7*#�7���I���@�c��y�c�0��Ԉ��*f% y45�#���@���Έ���3p��RE�b�p�W���S��l��F�y<_h6M�!���n��ٵ,��Qdi�=8 yu��ȿ���A��+nk�3��0��>[�z�D�+�����V�ӄ5v�CJ"nǙ�`ITt���^��ok�z����^��Ԃ����(���MU!$�A�z�O���m"Z4i�d7í�W��ԍ���3���g��ݍs�� �sWy�<,3�e�$�?ly�.�ށh�Š��zh��^G~X��Z*��9�vr&�e����%7Ջ�c$;�N������;�Q���l��ܯ+�*	)#�IF�zv}'��h&۶ʅv��La�~nJ��zV�c�=s�,8�P�W ��E,lk��/���%7 ��ǐ���(X	�+}C���*�It��bS��8�jp*IA+���1:y��A�0kcgyt-p*4�z�旤5ɱ�c��:)Į���J~��U-�.S�˛"]]�sk`�W��=!Ɗ[N*[k��l�"��k��0�*�Aq�3�<�3�K�Vzc�~E7k�4͛�V�A���O�ԃz��LX�^|4L��+r��#$�d��L�c̈́����Kh�C��O:⵻����2贈��, 4�4�K��2�<̞xY�X�x��vgZ�H�B�_��ٌ�w:�R|����xU1;I:��}�(����z'��M��Ј��x�L�c���FV|��Gt�@;�t9x+�ߒ[ǸY�]R�1�\6�����+	W^ı�Ǯvr�q�q��O2!U� �&�S�(�C�
&�Ş���&0z+м�
�����Y(��dm�.>��+��w��|6���xOز"�v����M�w�0fq�M�� �\��F�IH�"@����d��u�ͱ�����Ŗ�����V�J�Don�^ڛ���Ѕ�����\Hx����&��'��F`8�X/ԥ�� ���s2j��W�굖dc�~ې���a�Z��wS��n�i�β=3�G�L�ma�0ۣ_�qN��^	����g5�AnP����R��Q��������Q��J��l���L3+F�C���'O
�VdJ�L�l2��̭�Q'��:s7Y���}���Ɛ�]v��r��DP�����A��+��Enu(�eyx�$��gG��#�Dм�7�&f+���E�v��O}2��� ��>��&�GB����Ѹ���8�'����2�$YƔ!%?5U�ĺ/�v]��w��Ϻ6�X�kk����_�]��.HQ����J<|�^n�$Ȝ����Tw����n�_���G�Oތf04��	�;/l����cR��S|��#>s��qk��QI�P��{!
&���`�yby����M˖�i��I}ƇR �ۗG�+=�]l0��d���Py*�k�@�~��3�˷�0F��.���i�F�uw���ޞצ��i����hyK�����F&I���$�J���&M����a��J�7AǾ9��c��d���q�EFT��3�D���Y�G90��~�� �y��o�a�&�ǣפ�aW@�EU_9F�m��R��)M�s�y�a���UZ�����n:$����� �kW�G��@&}�]��ݾ�s5�R��m�^p����}nN�N�S?�4z+��R��	RN��Wǽ��lg��Ǳ�@��QC1��c��On���ì����E -o�r��;ji�0|O�M}pL�C��%�*u^�+�=:����֒ܞ������A*�(���7�W1��$HQ6_�l�2��C�w�Z�f4xC��էiGs��3%8�*9�#ւBs�	��sP���>��/$K9�*��'�f}9oփB"	��.�:��Q���ɥq�A�d��'�5�1���8F�͋t���
�ʲ�P���-zWyߟ�X"袽��л>ϐ(�~��;Gs����2��W�����0��x�H�sB\LKc%��d S���VĮ�ׇ�d%~��m�dn>��P�ȈE#��e� ي��]�#aR֑�?��Gc���8�"�H����V��+wB7�$�{�(�PZok!�F(��њ��b�,�Uq�v���������5�V�����`�����4r�?0��g報tA��0��7�R�g�Ӛ9L�5�,M��S�Ie��E;�[:�__Cf-Ĕ�v�"gQOg+C�W�؋N�Z���#��zg#<(�-P0um�	����1K�NA"{K����\)]�s��g\��RT���m�4��K�*T�b��V��5�Ĉ��z�L� �MeB�-fkx���J�C�'-ܒz1Z�i��Hؚ�PE¼�}�!����v�3�<Q<�$��Ri�h��(���k=����!�*�]dN�[�l?�
عJ��͏�0��6��O5����r֍"��{Q�9\����&T�:�3�pU��b�/�]�p��]珗�p6�����iG��^D�;�/����LK�����\���`��1Lp�L��.��#Y<�o*	�����>�_;��D8�߁9�]�vǝ4��j^�zN!#�x{��#�8ܙ���꜈rb1�M�3Bψ3&-Ч��D%��f�L��kN?�c�أ��^�3(-�ٔ�~y�9:=�"q���-a�:����!����D��r�Hs�m�CKx&�Kc��Hx@�z��q�X�D�*�9�]Y3!{P�i�8q���!�x����($�`@ G� r�[0�b�b(��<T�b� �[���֜�,?ͥg{a��Z#ߔ��`�J}��m�(}b��a�nNQ�plIi����8pԮͻ��9d�����F*A@�Y�I�U�'�-�$�|φ���2df�rϞh��8�<�T嬉�n���ˇ�8֫�P�hK)p�:7O��G�V!��������|3�{�(�����HKQӁ��$^���܇_�-�Tw����`��ED}�'c`�'���oM�\#1th�A�o�j��)1w��aXq�/El������1+���.����1�����9��$��/�E��fLn�n�[?Q%*%�����L��u��&�0Ns�b����^�A� I�ԃ��).���dۊ�Z�N,��'O�6�\�q��������`b�B�S.M����s$��Q��j��
D�!�ib��R�����DOPebUG�|	��!�6�Xs��cX�����tq������H��Js��q����Ƹ%]<W�-S's�-N�&��Y$*�CR����0��7s�C���mܺ�E�j��?�H}���}��b�U�YN�� �����s�ݦ���\��f��d������Ne���f�����ۢ�Ϭfߞ,�u10���ک�#��r�(L߉TU$�9���=���O1�E��7o���K�m�
��}����\��\��}/��`��
f�ʃ�<���5S
�S�^��H%mGl���rÙt�U3ךQ�h���`�N!�rjerkm'ژ�g�i�,��V��F:���#�i�b8;�[�&P�נ���Ծ����Rυ�s���5��I����U��¤qe
���m�m�ȓ~S���]�9sю�WY?w��UٌA��el�`�Ng�2�^��,�V�|��*c	V�{|��T%2��n�{�zE�YD��v�޾!�r�W��9�%�'B���~�����}���f�\n%����%>JY�G���o!��&�D\�2� �C�^4�~TXv���J��4�߿47��U����3*~8K5�˚ )cf?sc�_#�����ć���Bt�Q��yzș�D;��;u:�x��Y���:�wz
�S��!�n8н��̗@�<�z))��5B"�P���խ?�k�
���N��\}T�9�$�g��A����b�}�#�O�����6+�_���q���$x��g�,[w���S$R�OT��'C�_����7ųc�_�=>��:ңfO�^��7%7�Νym�|13.*r(�sj��DnA��_��v%��kt� Ы��_y��BQ:��^#>\ �g������pV-y�>����k�pc|��&��H:��f�Oz�n�E�|Ƅ���.V3-��a�3O��T+l��x��K���e���b揣��Ta�Lx
 zv�֧!���[��X�Xc�1�Av���:������`N����=��ۂ�Jc���5"�ʭW|4��˫2��ĩ%L�o�N�����Oxa��2�X��U_�u��!�#he���8�EQS�m*I�Ӆ�}�|a�l��Xi���z����n����ǟ��A;��+��%0^�R O.Xʥ{b0�T��[Ҧ|O�T��L��4�@�;�5u��m��llq5��6F���?{<�0D�L�
uuY�9������?T6��D݃�(H�5��:��R��׋uS������iwRUc��Ώ��D(!T�¾��ù5z����o�a�GA�t�f��9f�Y����[z��_r_O���n��1��77�Wo�ǏK���<��=:�������P�R�I�U�
z� ���n{j@�V)Z�#7���կ��[&
0�ҬX1~�lQ�8�@�����H����W'��Lz���iq.Q/�g�8D�}��o�PL�ߔz��1���+��kU�x`|��=_�O���H�8���u���#=��E���Ce�`�x��0�W���A9p2�\/xj^!��E�f�l�U��	��+w~�P_?_܎�e��u
Ǌ�s�_T���M>��LN��JL��6����d��vh���T���9�ůS}��0��A>>��832�x����E㶉�P;ZKs��n����@���@�[I��B�����S��^�auTf���G���s_�2a#��lZ2�l/�
h�6�ǲ󿇁c]�Mi�a{�G��)XSI�<qC�/%l���у������T���U�h.�A�x��1��] �����ds¥�ߞ�w�u��n�������̈���>�Z7�>�/)q��Z��!d\a0ڠ&�Nx�  5o!�\;�^�w~I��~
�x׆'��>֢��/���4>ν���?�"�*@
�:� c��/yQ�t �R\+�,R��(��k#(X� ������ڸ/S��1����w��j��j7�BУ��]nC��6�?�k��M1���2�Ɂ�s(<��KC,�rJ�z;�����i=��Y���
A6�S2K@1�hϓ��w�yf��@U"#��
<ۑe'��*y�-���h�X�Z~�蜊����3ƶ�k�Z��@K��n��jpt���~����'�\PT��Z��R�;��)���Z0OVgsv�@��D�h}*9�$)K��x]VO\�v�fv�ɬ�&U���O3FEA�I	W���2"��Kdu7���~"�z7P>@�+�qN{�5`�-	i�ݪT�ڣ3���aԳW�Kֳ��OD\�r����,*a���\��A��ddi(�_��\*;�쑐�/a�|^u�gW�a�s9�ߔ�����=PB*oU�QS�]Vz�m���O;`���=I3���_T(���H�� �)�:�#��O`�>�S�,�ԜǊ��Pz���Y���h�-�`yч�9������䌠���V�����=�K)���Y;+�0տKj�����̏����b��rV�0��
�JYhlc�*��6z��:�
��?T�t���xx��+����pe�;�b��6ί�3؎!���Kܹ�C�!�����&o�kص���UӎTHY��~�{���M���z磜#�'�03���5�~i:r�Z������CXE�K�9�K*�����L��ۈ�u�jkD�lR�r4�(�W��=�����d���~�`����{˞	����j�q8��qm���L�u���]�%ja��#A�������]ӟ~R��������Mi���*7��~H0��;H��wK�=����uN�r���V�4+��n ^�� :�U�����_l��1۞|-W�р� ��J*3m._~�L1._��/�$+����B3��՜�-*�"�r������p:�:�����=2%��h��	�%�2�4��F8���ڇ�R�Z�3(4��	�s��8!CͲ�6E�U��c�b��u�����y08����u��|y�s9�,�N���RZ�z����1�uh��Q�����4�Z�Fh�C�,�#�e���(�?�:���U�;Q&��U�y{�p��¹;uMc�J]�\f��&^�z\�*UAb!��f�E�j���������,v��E���a�`;��R��,��	)�ϼK�տ&m!������XM(5�:�=�l6����{uS��O��3��W�Z%i�9lv�/'��P���J&�2>.u<�b�Ɵ��Т�y��k%B�~C?(?-9.upm�� e������-���>~6�>��ˌ�c��&g�5�u�[��	d>�#b��j��*,p�~�w2�L����ӂLU�S dt�6bI����ӻ
� ;�}[��]g|���_���dY8`_"�B���ɴ��I����~)Ms�>�6����$��<E(s������.c�7f�� p+�K׺	�L��p���㽓�/��ss�q��$qGW�cr�_	.8WH[��D�t`�#Pͫp�;�v��F�~X��wĥ\π���ު�V��q��r)����L�IxR2�i�U��r����������v��1	��IG��]�c�.��F����u���7�\L.�,̊����o���(b���i��G�sw�#�'��Ӑ�O����Ϳ�݃CW���fp���S�Jp�I!��j���^+�1r=u�}?���XW�ܒ^l+K�}��f���\F�w����a9����g�4���qE�^��M{�f���>e�#��p��]���M��"�3Q�X�w�����\��������pZ�c\R=5����Վ1��`�N�qCU����=sI.	�l��f�L"�
���*��ar�<]r��wS4���6nJ�C�;�v������U�����}�k��k0�a��mO$�ZԄ^!b4ǭ'd�����bJ��.[�H��/�3�$>�7���G���Xt�����Ǎ@:�O�F����r�N8Q����cTߣv�ƿc\��Vb��ۮ����wx���-p��n��:�|�)�=Պ<����4�r��Op=i	�"��M��Ζ��8	�Vw+�Y�pK|��wx?)P���5<j�Sȗw2/Ϯ,ɶ�i����[���i?���k�kd��i���	� <[ed�XK�m�9/Ft~��.Cϐsp���\Kv�ُ�p�
����Dr�&�~�ZxR�6�H��с�̚�{)�~�� 4~3��I-�����n�Ǿ1�]���〆�YśS���E�t���4@����sϓϚ|���Zsi'��"Ġ�ݧ���PM�Ĥ�gP8�����@)����ۿ4�B�n�����n��]+�\�$���v�f�
�`g�[UY���T�<���yӿ����]Y�O�l�q����/���K�vT�S�T�CF��Ȋ���͊w4�;����ɴ��m���*�H���?�)�FX_N�Nѩ~SZ��l03�X�CjŚV�>�/i�p3���A�] }Ee��T}T��HV�Q3�����eH�1`q�I�p0"�'�wE%)���h�	~��E�歅�dk����4�h�@�4,��{=��,K%;�$�n���q�5Z�S��.9����-��Jĵ:�H����F��)c���MNU����sQ�:vc. -��i�p:�,��A�&!ʘx�!�Y�ئ��C<�3C�)踁!K5�֌��+m.�����o�}�b�o�!����X��ħd.
�i��@@����G:�Q���\$7�oU+4��1�
��a��M�glYx�6�]��K�-Y�`�/C$�x�����tQ�g����f�S_�!Z7�η�2���K*��pt>��/m��xa����^K`�(^T�W����}Q�k������U��:�=�1KL�%H�NFk�TFEg`@���8�F��¶�-�MV����'P�4:�Ra�\S�Y�@���4�h�w�?I[�+��J�}�V��>�9S�֍���ɜ��c����D�A?��`z	��g�8߂��vgOM�2�����8��΋G���V�l���B~��_O�WBٌ�>�VPCi���TM����L4�H�s��/���t�[�zYco����eV��?��O����T^8��N��Zl&VP���՝����?��ɂ��ma��ʁdM1��*}���/~�����a�NK�r�ؐtO����"m~/	���J�&a�륗�(��nGi�� R�G�MW%��<Ѫ�2;C�p7!�d�ꑐ��w�l8x�C�8����m����8��ZoJ�md$㭩��jJt��+����� Ow��;����2��C
����a�����,�� �{����x�Y�7
h����_Tc4��@\y�2X����@�-3U1�*�ߣ,�%nw�B��	��
�M7��k�k,`�c�.~˸rlׅP_?n)F6�(QG㿻�N)�+c���QK8�6��k�m�]k���I�Z/���R�"逵�?zJ��8�Vc�X�^q��-�sB?�=�7@$�@�`	��22�z�z�(�F~�A,W��h�3�O�k�}���o�����7�d�Z�tB��/;d��H�F���� ��^�祢@#bN��c��e�,(ƈ.�D8k��&��)���Җ�Ł>y�cȿ4���"B���D���05n��X1؝=��]��(%�3&Z��H.*0��Zj�I��K���}��t.X`��Í�yR��8�t���%qD0W�<}u͑��֡c?-�:e�s�(Z�%m �u�P"N���>���J�f�M>��x������mW�&ȭ�w�>n9?��@��G_B��S+6�P�,IM��dp5��6�]�րE�;������ q�޹�"����؉�We�tM!�V�yfa}I����j��H䙦S�Jt��Ey�&}e�顳1xsd�sXf(��W���+&��1$6~�.k�|�*}U��(䏟-)ΐ�,D��y8����Ƨ�<��k�zL��G]��v�҆O]�,�%=:���M�dE����xUd}���p�b��e�b���͙}O�Z��$ɒ}�����5d�=?a�_Q�$᠏
�چ�|6�7���a�$?�8Hଋi0�
t��^����y�D�f�1λNNܲV�i�>ޜpW�^�ֳ$J�p1М-"D
SS*D�!T�Zq$������uQo����=WH|+�QF�[��X.q�P����LS��:�4���/�	Go>  ����\����'s��Ȥ��<1%�_����� h�o�D�&�i4j�2%���۹ $6`8+@%#�"�hk4�̺�+�������$���&t��􏵘��P,4�	2��5q^L�ѝ�t��A�"�A:�%m"���/��=a�iS�Ɋ��e�bOEI�����*ʞ��Ү��=3n5}�=>�U���i�|ю�� ��͑���Nv�-��X��x�#�])p��E�����D��Wl/&C�ΙlېrV���8آ�Y�O]�k��+��� I��vE(�	�s�j2H�߾��������z��?F�C�`��i"���P0�&!j�uTl�'r�5*�R���4���6�[(���TEw>�(�=x����U�?M<[���d�L��t�$ܭ�uq�T\�W�p-��>�0I֝�n�q�[U������o_�#S��'��|����RՄ;��s��ՠ��({��K�	��PjV��n�"�l]Q0�R}D9Z��*�`�]�r~� ��R���{'�m�R�s�����6`aT"v���b[v�/ ˁ ��V�7(�{c�
��35����H:�i߲�H��iBr:�����:Ij%T�.d�]W?nCq�,=��3D�¡�(agz�7k��樅*:;�Nu��Յ�J6:сS�~��!ҵ���Ym[�c���h�c&>��JYQ_TA�6@�f�l�4[�(�ktѓ�V@�~��v�>�|���)�l;uZ�;��#UDi<Z5�mb��}�xB?�l��U��P���t�m��;7+%��]��`V[���B�"��ot��,f�A`��7��ܹ���wcA݇��8��5Ѹ�^Ș�(g��V�8�:�dvJ����!��<�ψ[d+͋`~=5:d;���,�sw�X���8,Q�N��xq9��#+�_ޞc}��UT�;m�͵���m�E0R���cK��8;۪Z���F��̛�h�o�)�9��Fo_�
Pc�CY��ivA�C�������ƣ����H�Y�Ɉ�崟Z����V��h�7��z;�DL��&���#Զ',91�C�3:��!�����.�`����/�[Bv�|��;U�����<��и�����i�c%�������=�Ć^s�B�%��>'���_"��(������c8��gl���yrJ.�0�ș��6�;�K��W>��3����~�ސu�p$gT���}���v	�G�pS����-{9Y�;���'��	�eU�t��$��͹0bCc�\�m���{#l|5ւ���#��`��p�oCbk�n{d�TS�XA�� �4{z�|�<W�n�z�fjE���F��H�y꥞�@ �l�m�K�$�I��
i��c6^�Gi�eT���ތ'~YZ	�z����祧�_���h�DV]�6�oiI����d��路���
~�R� 5�"o+ ��t�Y�h�M"ɡ_��3I�ɂ����P��G,&g���;q��p��>H���~��(M ���[�D���<��rۃ��:�U��Y�j��qC�{�[���>a�@[C���h�?�����E�C��!#{���X�I+6�6�����F����`2��ة��逰���T���6�� �}��*�q�1��r����W��8�YǏ�v^�]c�2- Ji>8F�%Y��Z*��rr�"�7��d]Tb~6i�L�d����H�>@7��	� �M/����X�_���e��VF��Ὢ�P�-L*��9k�[ѡ�m-���O��sA8]*ű*Qf�'T��~��)���G�j��;�+�����A�j�1Aw��@�ÖU�d�ż��6H�k߭���͹�Ű�D�JQ�خ��9��l���å�o���޻x)�	�.�0 ��* �-�����4����a�$tϟMڙr.E�q����]w��K$�d�.�e"�2��R	3��Uخg�<�>������8\���aR��3�S�z�#=�~��˱��3��Ėm�=/���B�����=L�2�$��K�-;������L�׬sw�s��`U�����{�����+�<��c7ߎ�d�bU�j�*+��J�x���no#c���݋�7K�UB�xj��QU__��Lm�U��keK��eX�/�!��kR*�}U}~�!����*熲�X�oڗ����O�l��ᕎ��_F�]���&pm�ᦃr����pb<�i1�`��B0�����Y�	���Ƀ.��>�M�c<�dX�"1�ZRj�d�nO��)FDa��+=|
eb<o8S��Aÿ���K�$1�dyy�%RR�-g��Z 0
XAuy?��r��)Po:�F��P���u�@��9.Ñ����ҿY
+	��pژ�-����gߙ���6���C��7��nIOJ
[P��lՎ�%9U�b,�'��)>�{�Hbq�#��Ȥ�EI�,�,)�{ ]�lU�bҠ�=�	�IQܔU_��rگ�Z	cNT[���$��*|c��	Cu��u�6��Y����v6��/��ۄb�	ZL�se���l�M�8��y0 ��i�Ҵ}���.r�����6iq�w�Ob6�kC%H�KL��%N1����/��f���J^h)
����3�C�x2gx�<+��Ё|�;��~4�1���n"φ��u�K�N��ϯ2�Z^R��%�.,I�K+�xt���<����͆�g�g�ʊc�G��k��Q��Z�V�k�@��XH��o��.���ɤ��af����2j��sV|��MaF����l���$�/9�ACZ5'L�<TS*��(t84�@����r�fp�*�(���J2HF܏�9$>	�E�����o��@��^c�A
f84����`}�n�5�W�R^�h��#�5�c�0#��X�>a�gW����]j1���g?SuJ��hAi
圗Fu�ꍪ*{����N7f��k`x~���ᘢ~!�U`T�j��^�P�?�ek�1PBu�����P����S��X��q5zE�L�u���Da�+������%w�����r	Q�6Y!Y��_Һ5��O�!G�wl�Z�j4"�:7^�E#ӊ|��k'%�֜�SK�R^�̂����s�'Ҕ6 u�5[��DL���#�`�$��@*��s˽ܓy0؎iXp3�����lE�3���)�ϕmI1���8"�ҩB$;fa�D�����T��v�7�w�]	b�jG6-"S!9��Ŗ��Ʊ�@C��*�=ΆX�0�~�>�<�2ݭR����B�h�F�4WA*�kи]B�i���\sfA�%������b��/�?W����a��$�(-n;���a�:�t�$7��ى��K�~��
��$�~T��#��]��ȿ�C	��MHϧ�<;h	��qЏ��U�+-�11Hף�_bh�����~�w�0�4�޶�O3��5��?��&�蒾�H�S-��:Hv��!��Rft\9�Jk�c�H�R�&���T�>l�|�l��5_�k(6���>���w�K���m`
�u?[���o��,ӏ�8�ɏ^����ª�V|��~n�]�G�nΑ�l�m��qc?D��778�o�Q��l7gڃ�dڸh�k�l]U4�����D��2��z\�ȵe� ��u$���q�ǬO<���l?�߳�����@�/w�0ک,�F��ٔ��H����U�N��7o/vk��k���7XS�P��󾩭,�T��Ae{�z`�1?�H��ꍓ�*͡�r��!������l(d.��_�WX�24��#�:�vÚ��(-���Lt����Q�*X<ۓ�>�,�"�������Q�¼9y,Gi5(�f��)���(�L{�I��؈Ȩ~v �N�e��T�Ɂ�����^��V:FmҐi-��ɰ\Ba���b#��7�r�"��G&��j
�G��=&���� ����Y��(I���w~ˇ�Rl����ӓ}�4O����!c�@I=}���*��Ҳd�Eք
Eq�,`�I;ܓ26�K��nN������~O��!�O���P�w���Ƃ,��0In�&��u\��n;�M�s/2ca1�4�ޘ���<`�k�E�ߊ���*��
�����Ҩ?{�Z=�E�&fJ!X
���wu�q��'�N��b	�ڟ��#��Fݛ�
F@�ꛓ��|qMvr|?Ӂ/��}��������O��w�%JB2`�l��p��k��\�AXS�s��l��(G<m�z�~�M�����(9e�;GCÄZ٧�6p�,�O5B�8���?�I����r\�Bv���Y?��Z-!,��>C� �\-�ގ�nq`�d*�L�b���L�!��'�3Tj`r}�t�O:����m~���
�t��ja
�y���0K�7'����|�&��s���j�w��dɩ���.l�ei�u�<]-��PN�����qP�~�E�Ï�� \�g������qnSZ��R�|Yo��#>Z��V@��>Z�{�EfSs�N�7�u�N��~Dǟ�ç��n������2����y�.>d�����-|�d�u�mʤ���K��i-�������-��/׻�r� �It���/������4g���=��'���#�7��8�"��aGmG����HN$а��`)�1u��&q�k{�� G'�Ul��op�m?$bq��1{|���De��Φ�78���2�RA��V��جlL(\ ]�O������E�i��,�~��+�ڣ.�9����L�d<&<��&��nÁe�C������q��}���۲э���~5	%Ƃ��&�V,|����4@
���1���`�R��.$ذ	�Y�[h�`��8�KD�B^���?M�<}񋐰�����kWߏ:��f��)����SٚWޯ���^1C	�IV8=�Nȱ�ɺC��BO/�[/�$�`K�������m����/ N�`�SM�/��l����8�<A+��G|��
h��͋'p��dgp���ܓ�����Q�!U��~�g4�D!��5&P��F�#]�+:�0�L;�����ŏ�$-e�z2��?L�f��V#��]�t��[iqS�/�)I�Xm6'zF-�th�$N�������~Ս!��`밬�*�mM��R�Sqρ���T�'�� wo*�y�+?� ��?AO������L���U�RX�ƙx��y|*�x�9^-��7v˕G;�ߨ�/��'~��Μ.�T���f��xl0�2z�4����3�{�/婇>j�^�h�b�����<�|�?�#'��	ʏf�-��z��BP��R�vO�P�\�Cs��;���q�K<��UG�r�#Q�ݑ�p�%�Uy�������-1�
T$�(��ҁ�8m��-T��o���
�����u"fZ|y���`A,l��8��[ȏe�^�`iz֡�
bzÝ��w��Lcri�ݢT�zy�1mՌ�XC-X�l���&a�@3&E�Ow�7������j����4�.���{X���6f����<��¾�R��=LO�%t�'�@����RF����֕�^��#^����#x\p������d�?�3��S����8��-���`$xy��G���b�[���2�#��D����ڥn63�+gV@6:+�h� ��`Ϛe?G��p�m���TE�� .B��z����YH�V?�����r�r�;�x�w�=Pf�7�i3�є��;��ރ\T2ud�D�I+�S[��5���k?2��O7�U�J�>z	h�M"�?�x�;dn	��C��N�IK,�nΐ�����\���?��k 9����jo����\�L�o���E^7Tt�_�,߸Y�������xA���$��`J�t@W'��(�?��T_T������ ���_�њ&Q��d����������gf�?壙b��%n��Nģ0KW	���ږ���ST�	���m�Q�{�4W5�Pa����uGa�yO��|n�׆��u�XӮ=p2�Psh?��°f�u\N�DCe�	Y���ڜ�rQ�]�q����H��L���62ش�i���%8�����'�^��q��Ev|��^,ԧ��?�ӎ'Lϝ��'RG~R\L���hi�����ѧ��>�B��ܴ��RE���SnD�(kWJ�P'��׹�1��Cd�e���_,��"2�.6'�|!^�6��v�{T:!z���;6�"K���	7w_�c�����#]��|��T������b�¬r$�w�f
�pV��:?�P?���?����I�^��i�*���7�ڈ,�b6`��bҘ����ގ"���x��q�$U��=<�ƻ�.D	I����Ν#)!?�C�iU��N��%�i������V�݄v�Æj�rbʋ�V�H*���.7��)A{�j�i �}��R��h����f7�rjG����Q����9��66
7R��x�Q\��[�n2�����%�ܯL�:�$F� �q���2�#�� 3ݹ��_g��5������$�O��ԃƗ����d����5�$h4��������/5R��!�,�m�@C#�N����#�O�g`<R$jE���~�(K�F�"SH޷��z�]�YiB���ƒu�g�/�y�A���{N��FW�Pl�&H��`��t:��fF^F�9���TªC�T}N���u����<b��N�-���k�ݵH����+����[i}���o䅺���'e/u��~��nŜ�58�t>���"����a�����#�W�H_�-������5�N���3��^pG�.�6����`t����(o	��]�����42����:�UV4�|��`�V�S��Gf�s~o8�V`���2�
�0��ڛ]D*H�AgU�
������`�G������X�r��Hs�=4�<B:9g�*�N�kb�Q�p���o�v[{ؾm!��5: ����?vs�Z��O�9����@3��7'�V����qt��wr�%^���Sy{���"\O!�Z��e�X}�MAĉ��H��F֕L��b��&;�Ք�M/�.��u 5��y�!ad~��=�:aP	/��u� �G�) �t9�3?��3d�%������s��LO�QM	wYZ̄!y����$��7g���)��@Tx,�l+j�wJ�T&$��t	�v���4�|��}��i��I9op�	�NE�`���'i������z�6~��9z�����R����]M	A
�
�棇�i��]аB��L��'�B�;\m�@�h��wR�#=�V����B�O��=4ufr��l�iTJJ�Iu}3��1�&M�#8K]<4��ט���}Rs�v��?� �m��R1��G�Q����ؽ���?9_X�x��#���˯+%�d�����q��\�Vr��;��{�e��+�-�®��w�.�)�ۘ�-�Z���M;�$^:ԡ��b9�e���y�S�m]�x&#�BWr�;|�'���g�+;���4fJVs�ay�:tj�p���`�÷2��nO\�_����=:�$��Z�<�Q�VV�>a
�u?!2k���Nǽ`e�P"
bꯝ����B�[�B��X���A%%>ZO���/��8���7dDO؋�]bX�G|�`�~({֎�[MKZ�%r��D�ޠ61�\�Qa�S�e���:�RT�ʻCM�Vlp����ӟ�^�U�ڇ�|��l"�5>��<�tAm��.�#�!�=4�%��U��PAZ~<~|�R<5Ն^�g@����-��w ��~/��mm���-�\�
}��2��d���@�D��_[A�6ht�x��Z �@pVF8e~�}�Rd�=|T}b´$v���ɮoXԲ(�z;���O�B�nprGZ9�I���9���܉�Kĳ���S��9A���fI+d��1�-x9NEOt��v1�E��:$#�$�����G�IǇSBn�[�P8"E����V�� ���h6���
�?YP�F���&�G:HqѥjO��=���L^�h�����C�__Km\��������R�"���6'`??z�=k��n|�aUI�#�i��
��y�U@Q1�8e�N�)_�����-�"���ͭ�M?��ʗ���r��H�f|�����<kŮ�E���cR#sP��I�Yi���54R�/-7�%ҴZ�4�3�I���7�L��H�.W����P�ф7�ɏ�6��V�=�*����ߙ���];���O����$5W(��n�ib��T��X��@��V }B3��n��O5Y�����V���kq\�\�ĶP��a��f9�X����9��A�^l�T��*4�e�{�O�m��)��88`޻�A�k!��M=f�����/O�W�lF�x:��&1H�vw�����g[,���ѹ��S�(��l8�x)e�J�N�ΓSc+�]B���N#�z�EX�pw�s��-�M��M5q���b֮<�vi�!�������wh�fH�2�D��4�����k	S�*�!|�B����h�<�Y/?j�%���̧�O�v7� ��l�-x�F��=�=�$v ��ʠ�0����I
6���
�%�(Y���� ˥��׷�twsηz�$73����ǃ�� �9�[ո "���W��Rc���Z�u�m?W���0�k�Xh�-��-[�C]#�/���������#�y����C�_��yUe���	$�
�׬
+����7Đ�۩��%	����n�|��d�n����
����"�$c#Wi�zȄ�*��#�a-C���<MiA���ntz���!t��M��)�}�{Q�jiwɢ���
�$��Iz��u"��U�1ҔQ�
7?��u�=d�; *BkQ����Gɤx�I�s��,
ǌ�y¡�������ofޓ�?�!s��Pl�����.X7�S[��F� J7���U:��.�y�Ձ�ڕGK�O5��+z
�?�A���j��:��=�8�B�\,s���SA;N(xa��Ә������%3���<S)�>��9��I�����CrT��u��mf�=F���ھ$� Ԑ�F���,O�b��X�E��	h�u�˻1�]�*�P��
n�%o�f� T�S�Mh�_
>��qtg��������RKsJ-i<t�&zR���5��}�pg�>>O"�{�";#1"�r�$S��[��q�p��ni�������Y��ֱ��<JE.�,m�e9 �2m�������fL�e�U��	����G�eW������ �,i��iX�I��+�Wo

�[*��hd�o�0��1����e��2���0 ��!ڶ�cu�❬v}�a+f�hCvc~[�6���O�mh鑌� � ���k��1���mǵ���_�-�T���!�f�����[�m罽3v�w�\�6��h��m�����K���Q���U�T�+�U�;��QO�C�(�|*�P��	��n�|<�y(:�{g��$COC}/��)D�B�#]�/��fi;�Uh�����x��r��o����(�����a�:F���SH�
]q��Jy�_/z����v�;P�\x���Q��d�[����q����<̄����w�z��јdF*���+f���R�<�:�+�D����%�K���,�`���Ӂ"l{EJA��¥�@��˿�s��/�6�i�O6&Vg�[�J?�ɔ�AE�f�����>�U�e�Q�^����ǝ��ʐ��qFkH9�p�ޔ���,2�v|sT�i�5���8�&51���ҝ�vڜ�:	�`��ƌ�@�ksV����&����ɂ 1�6z��^zu1*��A��('� y�D��8��<*�fx	�K�aKG+	��o��O�L?�- �t��/%q�R�\b���d����7>{v�H'��ɕ�/
D�%�����)���&ϱ����N�m�FJjX�Ǥ� �Ō�Ce.8z#E=�#����e_"���8����r<��qR�� ��;I;7V��ƶ�7��7_pv/�A�Nׅb��9 ��&/�������qW_"�*�9�P'O�B���ђ��X2�V<B�pmj���s������)��!S��}�V��nmŇ��j��b���1��]��]��dd�'��PP�+(�7�C��N��*�0,F�g����G�uS�1;Fn3�O�@Q�Pz:np���:_uc0APH��ʰ9:E/	i��Gk���uIt!W𰱰�Umv��.b���,QL#<X(3�z�nb��3�3�k:��ݔ� �Ϻa�Hc>-���چ�)0��y�2x;�_[n�
�c	%�a[�یB���n�j�m�0b�H�un5Xy����3���P~�0���>@�R����Y\ O�oM���"0dV\5��qv]����YBP�ApK�09\���U\�7��;���A���5eͭ �<-6�ں��'�7�����G6q����{��3Ɔ,�-2���I����	�г[��CN��oH�0w����L��?G�O�4�".3��H��z'��D)uo��y���p@S��������2\�1x?M];�w��$Rk0���ֵ�NXJ�'Ү�'�C�h�����J�vepw$I
h���H�l�mB��j���l=�(N����9Ǻ^2�
����x1�@��V�.(���R�}����)-/��<���0�� ��xt#�����9L�99)|�򜫨�vX9���Of}2�<:�N��Z��A��H~�����Mc�c�X| *M�y"& 0b�ͱϪ�Yx4��ScR5
9R4�H!��	O��ϔ��E�3?04F[�=%���� <MZ���)�A?��Xi���z��g
������z\Q�i�~�B(��岷��_.}�`��ٙc2�.��m�4qT ������M�<{�� T����]l�Q����c�d��@t��=��(� a*�qU�������2A��^ �HJ[�A�% ��ѓ����^b	C��i�x�#U"d=*Xβ�(Gp�_�"Q���Q���=��m�P�f%� $�J���55:^G�{H�85���R�����gZ�R^\*u��7[:�m�<[��� �� �f!@�[��>��v׽;�/�a��a�
N��M���<�y����,��"ۉ !��p:�֦�t��&]��9N})3���ޙ �G'*/`������0[H}#�z�I��.=B\��=��9��Ĺ��H�Dr��n���ڲq�"�4Q�wk��L���x�UieT���Nن�LF"��0�ŗn(CGU?W�Kp0�d�V�>�iU���^7&��dwtDV��/�+r�#�%V�M��F%b�E���ImL���\^<|�@%�$ݡC��*B�	�F/�O���+�l^���I�BwɦͬJ���CQb|;�ʽ4\@�P\A�Ԯ��{]?��}%��c���*Z�:��<��I98�M\7T`C-T��F$��wB�p�(|(��;Y�k����>ȥ��F��d�{�tI�������Mn!W8�͉Iy�qU|5G��]ݩݏ^�G=�J�z}_ǅa�$��6�hz8P�j�G3��G뛝�
��5���p�!�CKf�*aW��p6J�MR�F���9��:,>e��� "�Ys�ڟ�#H��@���e3��U����u����0�@Q�G;2�a|�Λ�Mq" �݌=r�ق����߼��e-��}���j�G�بk[�߻��Q�L��8�rַ��
"�%d�z�x��g;�*�q>򂻴4�-X�*��+��6�x�M������ ���r��ZL��m����X�}�7|P�����i	�N�u0�0�,�$9��9Xa��?8�juU�P�����-�wT;r_�F�?�b%ް �c �
��h/�1U9`�Ok�R51i`�ɛ8�!��o5�8].����o� ��y �~$ㅆ`����-OF ��J�>5�O����.�]�L]tD
��dT� 	b���B�������^�sQ}�y�|2�D�p8�FX����1'��(.�e�cP�Xl!�I�:��	V������ᨦ��B�ތ"W>=Z]c3S����5�KX���{2[��A�ʳ���@LT�R�b���P��'�����mi����_i@���Lۤԏ����aP(� ��/~ )��PS$��)����X�� ΰ+�oLG�B����:�r���`B�u�����4���e���ë�LdJ�:���Lt��ې@n+��G'��xr�&G���M_������k��Y|`tk�[⨮g�Y)���[v�e���=�Ҫ;O���P�x�m�?���0��c�-����N�)(�D#'�1�>����.F[��I@4��=Ecu��db�
h\?-��Y��D����W~qO-�|�`/�i>(Y��N��ǤWĔKj�߈���z����x�ϐ�Zj��$v���	��Z1�7�xǥ|���(��.�I�9�H��K@	z���x	��@�M޸C�F����w%.�痷HP~q%�~�q�RAjC�1�ֺx�xvo��e~�f�����~�|O�Ր'��@��l���7 x�:�R>₶��G�n�6���@�BN�_1	�wi�#H�;�4� ��u�U��pN���7B�9�	��cu�����������0��z3��<��������D\'~1,e?\W\�� �߾�~��� Ԭ�v�B�ʧtL��tbQy�FP ݇����>KH��?���se���q�Dk�=ښ�@�e�$�(e>�� �Ud��+N@�'?��u�����V>��ZIv��$D	_t�v�j
���A;���0�����+�%vH��:��V��� ����2>��6 ��l)%_�����SR?�!W�p 6�T�Jܓ��T����B�+o!�@��k
nsE̓ C�n2ڍY	r!;��x���؃S�온9��ś!��^`O�N/�qk<�>ֳ�ń^�^��	�$,�cB{6���1��>�	��������NLWŰ;G����'L}�Z�!�����M��_��@,�"|ݖ(	��-0�����݇��y"�Ƥ� �!VoQf����7����Q4<TL�Vr-����.��Hp�����`����l"�$;�������`�՚���O��H2k��:̏�ґ�|vT����tƔl��Ζ�EJFt3	���5��B1�\�q#����n�z�(1�efO�ֶ��:J>50�@�_2�B�Ƀڻ�o�m�Z�3�_����PQ/	�V�"@�㍮9$��������LF~ pYH�'���\w��ݜ+�4B͗ko抱�9�l%v�SoE+�ׅ�'d�A��}�~g6�iTG�@G��hP/��eِ�Yc���<�TԔ)w(�n:��y�^�v��ޜ�	�0'e ϲ#�{�l��cn#������	��I�>-6�xP�3�P��h@��1'��̍��<h�5V�o�l�"'8�{��i�vn�彅��a��@�GT��y��hj6;̆a��q���d{�
9Kq� r'�o�mP�gFRQ����6�%,@�H�},`e�q�w�	ǞSk�Ya���JN8�!��p��`*�}����0z�AfE �N����ET����I�)u3�S�sV��$�\���m+�$7�t�u�l�UWN�!�O���^���ɢROF��I�s�Q3/��:�����}��6�q�%�a~�.b1��{�\{E �h@��-�`.j�[(�8�[-b��J��>Z.è�nu�A,}$_b[Z[C�-��'ft�n ��	8 ��	���>��Zۈ�$��-Nf_��]_�j=�������o��>hcc����)NO�䭅U��95Vw�^�<��3@��D�H��1�mV��
rh8�s�[�~P5��Ql�R�p�%��!bm���Ӎ+�$F��� jܒ9[~�@)�@y���YQ�S�OgVSJ'v�o��ORdlޢ��lyO��/&2xSw}���-�k
�����V�]^'�W�Jm<CIg��2���*<xÒ�Y�:�P�p�`2`o�<��wSi@S� QE�{�:������ՑTV4IB�/l��F���OV]���խp�콸b�q�f�ࡕjN�ȿ��]�Z�EU�Q�/�$$j��T���t��DFo=��
�Gȝc���l���8��W �S�R�~��_���d�k���N=+M�X�^�O�Px���'����Y�֊��0<p���F����/��f�JoĴ�wC4vg�=_����IU�����=��ԝ��#|"��;�{��K;	����TKs��W=u�H�;kS$Z��$;�z�rW|�g%�Us�}~ڧ-{
�~���7 �~��04�+'�.���씱�_�TӃs�������j��8�ni�!�툦����뱣�}.��U���5����2�G��%&;��ʱ%�~Yg�C�8�B�J�B�1@�"��½I�� ��Ec͵��A�&%k	���5|g���K?�g�=R��������K�bt����;<��9%#�q�T�8��)+��̔����=��;���04~p�צ�2h���#Q�u`2�w_?�3���L�]s�ߍ7�0Jg#�Z��Ɍ$��ϺRH�M����v��JP�49It������u�/�� ��7�ν�܄+v�5�)|�<����X{��p�0R���l�,My��#5�6��x��s�G;�L�*�i���Qag��,A!eׁ_069���a�#fCz���a��"�"�xb+�j�C�kW~5�}��9ΉNr!�]ҫ�U���j{F�[a�������ڜ�6�/��#m��j��O^dn��8'�9����(��ᅚ�~�!���S%��ܕ矼�	4Fx��'2�U.���r���XҎ��ԟ�do�D�/O�@m&�J�}�,l�w�~���&y/I]��jr��o���ȝ7%u%ReE��Ŏ�Y�p!RN�'T����W�w����:rM��"2-f�R?n�i'H������{�����׶�"9x�K>��]׿�p+)}q>���ҁ��(��[<4k��B$����{�dVc��B��kzE��
�E+if_%��(��H���2͕3��އ8�c�0[Y#Ҕ0V�7���]eJ/pOD��(r;n��d#�;.(�BM�{��j�g��<�uΘ�5�|�%��?C�t�t�'N�AB�Ŏ�@�Ou�Kl�p��,!�O�˙N�^�4r��'�����R�f�'���$����36-|��SG��Y*�ax"��*� �t��VEr4U�Nz瓂�z|�m��V/E�Yx$�C3��n�9�vI�:A�>�3Ǘ��/M+����
kH�����i���F����P>>�;�X���EiC՛�S瓄�%n5L�D/I�m�P�4����r���G���ؙiey�8�c�.��������~q�A��t�����2f�Z;L��_3�F�h.�\^�c�0l����}1f����:
�0�����ԏa���$P����;�%ǝ.l)�='��s<b�#d�S��Iܰ�Ӊ�k��G�C�O�P�gZ�����CW����%޾ɻ�8g|��O���� �\�@R�m����0fuJأ�ם� ��)��x�U���+��@>N��n�o(�<q�N��X�K�)�c=�Q$�� lqh��ƪ�O�X<��d����`7�O3/�*�*�ɧd;&��`�g�PH9�.��mQ5{G���� ã�����r����<�kG3G1�ө��m�	Nd��Δ���,%�==���L� ���b>�1�5����#R��G�fj�y���74���aV�);�v�U��*�a~5 `DLo�"�QT�l#�®pJ��tQ9����.c�����Z4&�*ÆN-_�d.��x�z���NW=*yK:���UNH$�,�g2��~sj���M;Ze ���cMs���>gZ�[�94gY��k:�=��J�Q�����+xz�3���*4�0"V`�I�4��~^恭4���S�����ٺ�Z�Vt3xإ�-��q"g�ǻ�ZK��o=:�P1�տ��M�\���#���)�AؽJ���Ъ�f�h0�'h������]!�ٵ��"LPm.��b���@�ѫڸ��^��ɐ4l���W]�:]�!�f�h1���/**�u��� ["�aee�)I:_��=Z���!H�!\g+F�^��)>�Z�g�������^$�^"�o �0�D�o���s���pF�%_��������߭�Q�}�@I����X�l��>P�:P(�>(�4���E��\}�%,G"�:��O:9���Ѓ
5	'�	q�y�˗na�`xܻ�*��wGM$��In��YBZ�����Թ�_���6��b%)�w?p9\c��~�&���+j�]3֟���������{1%b�y�,���q��R��.�j�	8�:�ԣ�w@{����Č�F�T�i�����)ı~6�E�+�PTP�?<7���@�~�����S`R�	4Xie��e�lVU�����"�
��J��--B�`ᯢ�$�ќ���E!#�;軩WNeQ#�~[�\-G��Mv�H�O�q,X��kO��y��((8ס��~Ɓ�y�rG,k�ڪ�6�se_Q+�H/���u(r��!��{h$�6Vԗ��C뇓����B-�����DU�Ge�L�}S�P����I'�XdB�j�Wׁ�Sd��i����u:��=ah��ᤖ�T.�F�ݔ]�78%3s�#��ǎ��c	��(���8Ӂ'җ�S���u���������x�ߖ�@�o��B�.����[�
M���#h/�_hMKB
j�vp�s�*�y}U�IE�4^�ZS�`��h�(�91���q�pv$�^����
��I����((�o�z"�i��iȥB���mF;D\"�?��K�.�������Y�iz�]���
_���۴|K �)Z�D��Z~'���2(f�3�[��UD�y����\�Q��������h�w���loJ�Y*yb��Q�a��Ro	�x,5���	""�%�rP-�i<V�ş�;�$���ՐoA��ʸ1�%����+5|�x�J���1���Nf��&f�����IU�%�����h���Z�q�w���m&j��t=!'(�nB~�~�-�IC���[D��O3`@�wCgS\z�8��y��X��䀃!���7*����O�Vg���TJ.��n�;+ݷ��*P5�Me?���78��dA&͍����d�9ɧ�^�h5��{/����v@4�M_3^َ�>�g�ܗ�nC�	�xw��;��:߷=bGe�%�p,��8=����uR���O�\��!�60��u��*��I^Ǹ��Duk��������eZ��Vr�E=�ЌO�SN�>�޶z[�0n����;�5̣��O�YB5/V���Ԛ{�?�#C��T���8���!�����WI���[�Ёu� �T��G���[�Z�,v,��)�iE�*�"���J�2��j�� ��Q6e�G��K�uQ��3�]x��*��
jڇ�ߕ&K��Y��@a2�PT���Z�)�@�t��RX���Ey��,v�2̎�^�L�3��OR��+p�T{���1��/���5a9��{Pv���)�M�k���]œe{FxԈ+{���7Y�^8F��b�R:��ԃB'0������
��B�Zx�^f\��Ӈ�WJJ��&��@�8GW��'���}�j@&VD�SJ&22�~�QD�p;�>D,E E�w!�u�TW�oK�m��Y�FYp�ܶ���I>�d����w��l<n�HcM�Y�c�Rf��8g�S���b�>�n�	�����D��f���Dg��D%*�(����[��ʆ��S �bU\�}�����?U�ו� :mQ�|��A$X��D^S�^H�3��c��c8��-������ԭ�+Cy���oki`O����dka�[س�X���P7��^�C��Z{�7����o���漱Yf��d�ޒL�O�����T�?4R��W�4|��V/�@AW�`�k0��n)�3u���+���\�@�D��!�/���B�yZ���Jn���=���&F�A����;��3�"��-���3���+�ŘRX2�A��I�t���y�/�|<��?��Mh'�Ȳ�������|M�_��T�J�9[���I�Ui揅k�G!�&��1�����Mw}0=���M��/W�ў�:�
�F�3&'�|ZEu� $���'u�t�����as8���U�50��?��c���Z��t�[z���c�݊w:ط��V�4�e~4��_ӏ��y�+.�"���|욉qZ*ݐ��^��$ c��ւ�ϾP����ȓc}��z���.���2DE�t�͂L][�U$��R�;o�������q�n�t9���<j�'�f��i|�"��g�t/~�[/��� �Z2��|�>�?P�,ۣ�`�F���E!m�6˄�he�1��<R@�ϞǧH�ݍ�s�i���UbT,Y.�{�����]��\;�R��7��	E쩣Xs��z�J���l��]'�?��[[��7���3F\�owT-ڈ�ͮ��A��QZ�&5&UN����L�!è���L1mR8��Hf�#��Ɖ����x�����kc�Foa���)�;�%�1�
��ǡ� ���,4��6����N�\�p�Z��(h&�u�E=	��$p�)��W14\���zU�@�1!O�ر3�w�9eJ�tr��a_�g8~?�Oݲ�jLg��9���ZC�;u�LXn�����/=�OXàR%�$��N�ܓ����{C�Ԁ�@'�{�� <�Yns**�J�(��*��G� qR��!�$ݧ0����Q�n 'jl�5j(���A�/2�٣]\�����~�IwʦY���c����U�x�C�I���p ?Q�N����b�N�W��̻��I�� ���&ݓ�w-� +Ɇx�Q�|,g�����Җ'q�i��Iq��=�L��Q������a�#����7��,+ݕo.U���B��Zu��4���"���5Ouw���E�1������z�ຠT��~�#>g	7`٨�_���ix�<�&g��`� ����4)�x���ɒm�`���;1M��:��L����L�$�va�m��#~��ËU���4��N�}CQf�2r��@K���g_���$�EH��yq�2���J$]P�<�^�n��Ako#]��bM�nb ���k�V�9�_�E�lDS4#���9����o
my��j�;�:Ȗzi[\�jx�(�gw�'��]OϨ��m�P��$�#�'�v|�N)�K�H�ڣ\�ӿf��%D_���Rh�tj�:-�����b����QW�P��[���Q���@\7���*N��W�7}_Z���Ke��p�k=&�sB&����$���ىA�~#�y�ŦG�P���8(@~~R�]9���?�,K�h�
�8��O"�09w��Xe��3�x�gT_J�v��ǼĞ�L�py�(��T�`��[O3�z�$I��K�E�%�c�!�`�s�=��d�~�O��F/
Esz���
i6��m�\���5�;o��rF�?CU���?�p\��ĻG�8�ϧR�aƚ��{{��pZ��|�E:��j�'s��4���ƭ�I��q1�Wt�
��Ta-�g Ш�?��>��?3Pb���@���t�BJ�]GcIa%�E�)(��d�q��n S������IQj~ǉ��n���E�d�����._�X�*����i�6ɳ��ɪ?qb�4�.K2�D6Z���H��$sC�2ť�Qg�+Ч�(^���h	y8���IIN�3h�f� ��Ό�d�����}~�Y�r�C
^���B���R:\���j<��6�SM��j,��S������K1��+g|����9I�u�+��DQ���`>.ph r�{��k���!�\�j��v$f-�5��M������P�z��	{������N��X�?��j���E��K�.���oQtJ�X_$�S͇j/j�D��C�５�J��%����y�5���ҍ��c��	l	k�w�XӠ���Q���ѻ��H��Ȕ������R��~?gE�6&G��ٵ��~4{�r�YWd�+���Z�R�p���{k��F�E
&�]��� ��L,z���]�6$MN;��BJ�:�����~�y��#�wl�$�2fL����w���h�b�2
:4��������2$�	q�p��6��p�����I	
�&X��Ӥ�Y^T&�6�Xáw|l��.~�3q���F&-�^[0&Ux��9�T��xGR�f��2�_����̍@��8|8촸��E�%TS�u ���Fޤ-n��˴��=2����%���mh�ʡ�DP<JUXe��s�Ì�jB
;����۾Iyw��p�����|�,���R�y�2{]{A��	m �m_�E۰Eĝr�!b�(�L~p�K7/���7��N�p���d��^��i�?1a:ʚ睓���	��3�w�%R��n���������1�1��ػ���[5}�Y|�� ��4�b��ꌨ��غ���f���8Eo3���� �V�ֆ���.!�n����>IM9�z��1�i����=��S�7�mx��f$��/��S�8E�n������р.:@O��me(5�$w�����rˌ#l��l��:Y^h���;�_~PH١D_�9��{�8�\|�	R��M��j�E�t���L7%b�p.\JX�HSн��nH����鄝�O��)��Z4F���:�Z�iA�טy+��A�� N1#v��Ȓ�H���c��25�X_�4�q����Ʌ�(��Ƥ����Ԡ���LfȈ���<�|&�!#��=���K�@Ј�������6U4+Ai���d����Ǌ�V.�����8�et�"�a���f��6�ݘR)p��Dd{3�
��� )����d��!f����`~e�Kb�dqW7Y�c�/9�����b&�����y���Ō ��oYr �<��@�*����
E2q��r���͑��U��%�u�<���e���,=�҆vw�!8�� �$��ۅ�&��(��Dڪu����J���(��w���j��q�n�ަ�a��J�����O-���[Q5!��'������W�ʽ�)h���P����18��F���N�3E����u�⣆;��+�XS��%>�..�-Z�,�#	Hs�w��zL���"6�z���n��a�E��lK(Y��|	���KYR�v��h����&ܡq��A%�I�a��vd� ���B�j�e�GC{��H�������3P����h G���R�ᢖ�a��a.��3&�_!�]18��t�[|0�I�6w;��<��X�g�a�1"��pX[[�X=�P)q5�����C|��&|F���2ףw�j�d�����/i�i�����<�Q������WX� Plh�E��40�p��܂L��I�G�V��*��c?q��3�K���� ����2`���(j	����N6�zZK��d/o�jq��T��vU�S�3TlD��w��3��O�%}0�}ԭe&�s��@y[��G��MΏ�Z��8��;��B�����=<�G���?�@F4�:�k�=�7���=���u��f�k߁�њ�9���iˢ)Ҧ�5(3�����ʥ��e�TA{6������C���-̜���� DU"�s����]\˚��C�䗷t�\�9��� ���J�*���^y�F*�uKPz��<��.u��B>��^�W�����1a���z�
��69���>V;H8�HY��@9S��H ���/���U�������B�j�y��@X��te&�pe�F%�BJ_�|�ʧ�v�co�����
���3���S��b.��T�k}!~�l7�g+��sdn�Cn�L~�Q���X��B|�O�=O���k=j��8����r�u�Y�f�$���"\�6�@*�������Ci���A�־rʷ�+��U��[������K�+)�8LK��j������5,{�If���q�
��oS#ؒhDf��F��Y.؊�յ���!�I~�n���n�HwW 06����q�e�>�U�]�=	�_�U�a�h�AL�o�h���Ë��O`�p�fU���!����섇��v�v�a<�T?�ˌ���Ne�0[�"�𺩤ۉkG���XZ�e32��[���{r���̥b�Y�֓��$!��`����z�M�c H��ȯV�T���j������`֞x�&�=�`i�t�>86z��m�F	'[���V�W����j�/7��f�pL�,k�nr�J�*>�[��x���r�Y�.%�CF�Lև��� 0ŝAS�vy��r��~ -r�m�0���1�"f^߈�>�S��R��
�B~=�%o!�8	$����݅�6$��.�od |BD.q��AbkrF�'>�9��@j݉�,�JB��'��j��2� ��x4�,�W�8������]���qy8��uUd=�6�����|C\��]n{����M�s�D�JÝ��0��Du3�U�������%!�=\R濂"��ckJ���x��$��d�g�O���^9�&���xz��d�/�ɩ��1��~xy~�@Vp���n� � ��X�FY�@���$�r�������N�\��r⊄�V}��8s��A�4���m/��Y�t�]d�u,�ҹn�����)�m@kU���%H�~,��{��_��l���������l�}�W�gx�����W�o��B���&D���h���I��_�VS遳�a�?M���D��\FH�%L�/Hگc���t49�lf�pҘ/����� 㨤��:�t�-j �6S_E\�9'./>��<� ��.��p��.�G�f!�#�?�^�s���wڽP�]?(�~i�U�|.����sKNu���� �~��z���D�Ч��pǦx�9kv��4���n&�T���'�V�]��"��ƙd�@|�`p)3�qO��`��ֲ]m�v��~h��Z$�
�Oc身" 7�×h'6'� m�,S9W��#�-��7�s�U��<BE�u᮹꼰�����S�Vg�|��I�J7��"�?Ǩa����|"�ө�b;���*����xw�)xյ� @U9a���@����I�ֺ��������d�]�H�g��&��<�$��̧�'#/����$B-�Me(I�M�9��z`�C�ÊŲW�KR B���GT!8�d����SWU�OD��e{F�����.�W��Vo�&�,l�i�O>��ر�vnN���=�B��w3�K 1�Jn�������+��Y$1@�5���gY7ݴ4.+I�u��E�.�K�b;�`"m'�T�#}�iPm�#)��K��OD��j^~���Ah�)��9G��'�egp��d�] S1g�P
 �	��� -��?3/d���wప�9���O<M*�BZ�4��.�k���xb���//��M0��{�c�;E�|$ji<��6xJ١	��:kqWC"�����=]�Ҡ��e�tS���Q���56�Xج�-@�T�+ò8�-��|^:
���V:J�cWR.ßP$�0�F��g��[L��nXy�6�Qij��|ՙ�n~�wu���� -������:3=@z5�+.g��\�8��/�6t��z}��==����,�C�޽.A�w,�r��O�*Km	Q��2UJ����8����;�ļ�竟�Ht��@;��n
��b�b�lM��N��R(�m &6s	h��7����k����x3&^�"b~utӆ�d���f���WTsJ����+���ze�����q[�����j� ���S���m6�S��hX��٘�TM�畚����恗T�+�+8?�����g�)o�KKkR�"����JV�|���L=A�x!��b����7+42)���xL�����(���F�Vm��F�����u�v�8�&*�M����Ǌ�1`vg�����pzV&5`��$��F=����b�����
K^�c���r�Q?�v����&�6�5ޙ�CS�"�������y��/�(�����xb�#h)�l�T��kQ�= D.I�D	��䓩7��z3�sR�w	U''�PvȊ�/���^�4vs ^�PЂC$�;��}� ?Q���9�X�f�h*�/ ��^'C�<� ���c��<�"��ά J���t�/�>�r�9/�ݪl-�Z��8
�"�<�t��QY��!�p��:W��f�j]O�˼H�loY�C*!��H�����>���߭$uل2���]l��DG68�F`Uv�68s��Q4�a�MF�f4�,��''.�U?��s�;�f�	���(g# @�������qA~WxY?�(��}0}�g�_M�
;
�~��H�tj�H�8"<�&�+aw�˧vJQ�:���924/Y��C�t�����L�Vt�c�3���n���BQ<*�3�֪zT�O!?{$+��$_�E�Y���5�LR[�ֵ�j�en�:���kHG�T'�5�/�D�2�����]�t�c�|⺭B�cYp"( 7H@��@�>��wd���9�q��Y�x1�W��g�=��빸KDI�Q�����,]*�'��*�h�ꎦ�Iݰ״��Z��R��Ɖ��'�b�Rݽ0Q�� �/��}� �+��Ԁ�^K�7 ����^���5�\��n��G�9��)��53���w	ө&ǟ�\�}�w-򬕇�;��%�h�����@����-�i:��V R2 �ϳ�\�9�'i�Q��ǇO����
Ɔ<��vM��������B�/b��0�W��7��+���V���ND�7��EL��B�ĝ�4|t)LI��{�'��e6�#w�Y ��q�������]-�e�=�'Q��9^h�*M��q�e����QL?.��[i�5��zb���T%�/E�vx_��k9�OG�y�w��*�>���T'f��Gҝ,�$+����D*SN$e�@�t'\[���C����#v]*��Y�i�<VM#�^�W�u)m0݉&<�:��(c���h�%��gi����c�t����U��IB&�`���Z���*!���rE����Ɨ�0sK�na�ۚ�_��X��N�29���T�]�s������/���O����A��a�8���w�kqR9�Mߨ��vF�N���n�G\��<����A���fh���9gG�Nq��������t��$���n/1�9���~�Y� A{�rF`���8j��9�σ�{mQ;��ԓS���<�<n�i}5���*��1z������˨�`u}�������;���*�٧�B���+�'�ܰ��,�g�{��F��D�������^��H���Pk9M��P\E��B�|�cZ�Ċ��iR9�/A|����BO��ڹ�@��/Õ|ܜ�d̹��kR����;����X�)tS������d)z�;=��A���[W�o��U���:�y�܃cJ	�V	Hv�'����C	����`8u��((?x�gG�%6с~{�����Ԁ$�B�h��+���of��Y�O����Ll�;I[JG�h��؂�Vd��RӉ�)EZ�biwpwt��V�JH�ֳ��@0w�.� sfhD�7z�n�l(��������1��[�!�4����iu����i*6jg�H��7�J�"h#j�IEHC�#D��Wc~�!�tԶu#�g��#�����!�h�����ay�y�Q>��Xdy/
~/d$��I�[B��}���L���m��e��`�x�Jt�}�A�#���$�q������rR#^�7���a3�����0��2�����TO���jV%��O�^�ͦz�eY��F��~٭o�~4�CC�5Dxv%���@��D
���c��B���Ҍ�9H�RF�c
�g�·q��:����v��b�x��"���/m�H��E�Eg�H���h�4Z�d�hx����v�]�� ;w�\���4D�"��Ș\y�Q���T'?������[DĄՍ#� .8���C||}�ұV3��g��&�������H�D���~y����������ڶԄL��-�Z^�z�G�iJ������(֢p4j���Ay'ŨOt9΄'�c�z�U�Q�%n�IJ�x�ʻ��w����2����!�S�b�-��T�@�p�@A��82�O@[&���K��);B�/��YgVBs��
�?ZӣfN %���\��8-[ m'X�1�PP����ٸء�՞�'A�w�]�/�h�W�xG��}*�\�!��}M�����y4�W��b�g����KU�x�G�O~ZkaK�"�b{_������#JCD��S6��ͣ{0I�od����zO�j� �]���$l�Ta�<+��ߐ�n�m�o�#��gn�0%G�'�=��C�G��[rZ�t��	�'%l�r�=ᤲL�|D�^��5�!W)l��9� N�������㈞ٟ��}}s���6�K�M��=w?k�����}�S�WE绗��'�NT�z?C`h�<*�ӛ�ev�@���i)���g���Y��"P�5uV��6�{��:W����U�M�.�`lYdh��>���/�d1�D��W(��ȸ�x��.)��
�q�
��bE+xA 9�gh�w��1�����>Zn��yj>Q���9MT��F>��K��� ��g&-?,
h��8�a�g�#���a[�\�M ����L�U8m��]ڤ����%͞u���	١�Sq�#^��Ǎ��n-��%���$v ����F�0�\��Fa)<2�,��
َ:�ʚ�m���3P_�r�5^j()�^�F�q�2�}p��2���Өb"K}�a���^���zx�-�#4@�r�J_���sض(�9�BN�%- �j����o�Ŷ�-D��Y����ڠ��Nd�2���|���Oq�V/�r���d���T���tk@�蓍u���z�O�'�s�Z<���l�c��x���5�G�)�J��Q��3�����WD��n�̛����ֈ�L;�f������wS��Z*��9"(���5�?xo����8����n�?�h�,��]J�eGmU���PQ������^�^.�2]s��>�����{��Uh~Ò���8�V��pm1_��� &HdwF���p��Ҟs���C����w�� �EB~�烱�|��P-$�'K�h�X�����/x4���Ӛ�/�N��u7S���l��-t�����B\��ؚ�<o���f� ��Oޡ`'Zڋ�KM�_�V&X.��H�xj��Ft�l ߧ�D�={U���|T	j� 6?�+y�����#�ա�M�xïH��ύ���=�j�O�|��z
y�Aw���(��
.vT��OSꇋ�/)���2g�9�	{ʴh�3:���S�s�jm��h��������fF$hKA��IC�.������p�Pam��tA�?�<�h29i� zs��\����n���#��d���-~�1A�崵���(纯Ҿ8��u��:�ݏ \UU��U�D���٪Ћ}z�P�j�m�cV=}b��|?L����M�aGupT���|�0�8Gn'�a1:$c2����u�D�he�aԨIj�z�����:5�g�PԴ^C�<B��Ɨ�b����n�9~̤��r<Z�:@_���q��=��GIo�{��3��0F���d�T
=���䀯��(�p�{������/�Ze�x�^N��f�)��:�	,��ι9����YU��r�cZ���(�v�G�~|*,FD�� "z5?a�@����+8��dE4��_i��&�@����t���orؙ#�z���l��
�&��D���.��T��G� 5�D���iR:��~��m�v�����{��T�Z�B�t/����C�e'*^O���d����s� ����i��D�Eϫ�٫�K��lc-ʚ��H���:��v�#� b5�of��"�'���1G�E\.n�c�C���才�n�0F������QM蕱��mRҝO�K�,̷XH?��XU,��|���ʣ)|��G�E���������⫴�nq���x�
@�_ �����₨>l��Z�����)��t�!�����wb�]I�`�����.c��Ħ=pJt�2��h��>ߗ�����Ϊg4~�Y�­���*8�6��V�)t�(�E莞ؘ�Q�C��	s�W��{��?��E�DӮ@�B�`8��9,~M��]?�T���ݠ���m������ۙ'�#��~�Dza{	�ښ���#&Wb����`)^��r�m3���� D���dx�:D�fL=�,�� ��;����	����Pt<�!�pq7
�T�p������6�1C'�7Q�?%^V���F*��ȅr�� ��1�:�v/�tsol1'��e�e����w�5Z/�0޵O�j�J�Lm˷��=�%.A��C�*�ڦ�;� ��@���4EL�����q �rZY�	��&�gG:I��r��׉�m�Ytn\n~�qd8⤳��� dv2g(]2jn3��9m�nU�,�I䅸�㔌�����o�����s�6eqB߂���˭�d��J�>���.�I��otM��g��%"<E��ޕ�u�������"���DsΗ���M��递l�ŬKS
Zq������1L?�B�ᠯ��IB
���?�6�{��H�Vf�4u����v��K��&�T�fSp��/�m}����#�,�H�m+�K]X3i�G]�W}z�E=m�[dWZR3�n��q��Z7��Ǭ,���� ��dAf^�uJk����E$0���%�"$� =��zk��+�Gx�v��Q���;�M�7T{�����wcm�aT�UT�k�˷UE�GM��J���%�$62�J���Ú�x���Ʃ�^����T2��>CdW{��jQy�n��%��V%?)�5�8M$)V������$/���;}Ч��+.y�5�-�u	��L�M�%A���`07��T���U$6��D+���}n]S��{������eՈ�𻐚[�}`8JBo��L�AP�9����f�9� �K���E���/�Y"z$8E���O�.�$IA	��8��A�}M�����,#l��1�WK�s�V��3��#c}�(CS��!.c��D�f��`]�+�=��6<|&�/�X��Jo3�N:���Q;�آ
��%���2�����_�a=�t�����\�~R��B�L@�*Q�ᛝ`o��i���]�-y�WiƙY*�Cёr����
�f���7N%���@��>x��nD������,�B��!���2��,o��̣�N�Ss�T���U��f��F&�u�c����'�N���/���Y����пw�� ��Vb𠆙��$��*��?*;����]��J�Zu�c���ݮ&����WD&��Z@K�&��r��^j<�(��<D�S�v��)�c����8V���[��a�[	�qLTa�\L���l�â��Gg��b��qɹ)��9�(�j=��1�aܔ�E�ܪCp�����j?Q~�Tʉ���^N�#�myN�*T����J���ҡ��@�������+Yv�p`w�f���
`����P����R- ��0��;Ȓ���*I� *d�J���d1��7�O�<Y�?���w�=�����M� έ�RA�V���ۡ�����@,s��B�`��U3��8ܔ���嗆f�.���KCQ�������1��z�ٱi����SEE�eT���(��O!I����4ud9���}H;� L�>|����,Ӏ�n\S��Ru���i#�"Х��c)���`���a"�X��\�����P�Z9I��a=#s�3���_���h�Y��r��Z���m���
0�ެ���W�qĳ^(~��^�a4It?��H��);�!�ؑ��*.��36L��7l��UN�Q =)��q5�`^�A��|b��\l%�ie��xj��X��kNY�9���՟sfj7jSNf�.����B�o����n�l���@����&�Lk���b��Wf�rb�l8p3U���_S#���5z��C�X�'�U����|�;+:L���0|���`�h�9�a���Z�J����,1n�-�7<wس׆�zq4��$���5���5���㰾2f0�L��Z��������[t.�����x�BeGz�Uu��^ �V?�.�����*Sm��!s��11���㝆 hl���_!4'޴<ʝF�>�����eWA�����%�2,X�}ܿ���E�T"X� C"ut�� $���u4ҦA?�U��KDVs	����j;ͣ��쯥M]hm��	7���Eo�����1�p������Xm����"�j�+�Ā�;5R���:}�U�����k����#d���a� H$�T70j�J&����6]�)�*f�
S��a-�+Ӳ���9�}�wHL��{��Թb����`c���T
���,S0_熥,W��G���=)3�ƿ5鐇�οF��WQ*L�5�:7%W7�!��@ؾM�?���Ȋ�V��]R�t\%ӻ�z^��8�b�s��_��KL|�6�٢�E�F����wQp�Z�y�T�� <쳽�J�٦u����j�������>t���W�"u��(<�1�xA�j�q��&70�0G��8HU�B/�o7�2��>c���<���p�a�1Q;�Z�Ȩ*}����L	�Ͱbm`�HUh�½��`~ߎ2�C睿�����G�.��	8�vW��n��ť�]P���h��ZP������릁�X���yk{�Sz�X�|�]�,Z�%��h�O;ކ�W�ɨ�@,P=@H���/�VV�[����=4G9�	�|�P*��ل���T�)n(���%8{�e��n���c���T{���K���Y�&�#!�m����ZD��u�ۻ����Ƭ<%T#�j_- ��'���_U���f��$*��R/j[Q�dM��X��d�g��lk��M���W�"�h�0�W�< 8�r��0(tg��bU���>;G(O��i 6]�u�k8�ף1'�oi����T,�!ª�/����tż8��]�}�<H�m������`T�����u��)��]��"��x[�^y����_QI�����x�0��f�#��d;�Km�Ćɐ���@Te��N�znS�>���-E��-d�Z�C�6D�����K��a�CT�퟈�!�X��o4���@�,��p�';d��� ��psE��.�kj��cŨޢ&�q:�.rv\l[��:J(�[:�Yt��)[L GX��)h&�s����[��D;*B��Ok>������M#uL ·��,��gv��m�{����vO��G��V� ��������rt��v�(R/&
T7���^59���՟��Xd*__��&����9�O�(��.�i(�z��	GOS�aR�l�]�^߂G���������G��d���b9�UhPF޲�ٶ��q�.gkž���tf� ��W�q�\֩d._f�y�����ġ
��y�Г=����Fg����i�
�U�DX��:��9��!�a)!��:�K���`�����N������*��;:�t��w��+�_W�>�FW����E��qƣ���]��k��j����m:���*�\ظ�v&~*���q�N/�`\e+eǏ�N 7U7Ϟ������ְ���x5�S����k�%�lb�.*�����<_fA�ֶ�5������K$�^�9�"m	b#J����=��o�uq��N���s�:Jry.gjיW��hqPWNЗ�����x�Yɔ''��֊X=���-��)�h�U�v���1�3S��`��7��>��� נ�>1T��Z�$���� ��ml�w� �'� ��{V�E�%T17����GZ �m��E�5Gۀ^�J�g�K	����L;*8^� >�q��̅�}w���?��ǵ'����1Ux�e��XVEp]������r0�wY�u���S�K���އ����*:��d�z˛��z�?¤/�z0Sn����2�kU�J6�!���_���[σ���3Ώ_
�>����p����%������&;�������6��Qa-�7�@����/�
�v�&hPs�F�uCOV��m;!�ߘ�K�P*j���v����sGRf�����8%�X&,���9wR�MC�����I�6ژ�Q"���\Kd(E��|��:j82��\��Zi���z�C��ON�G�8�*��aP�e�jE�:ݤU��N�.�����d#�ø=����]��c��9�{��W�Q���Ú�w�3��[��X�[p�-L[L��	'Z���YI�Z��H�E�ըu@���߻?O���`�������|���5��x��\������%��|�i�<lZ���j�����WRց� ����S�hY]R;�٦�����F�t@�%���5��1�[�ᬠ��t#��F�6�:�R��#����M��4V��p�JY�Ь�����~V�Q:�Fv�Ю���-��+�ƛy��wҷ�[�����8�F�P �ᇜlil�_�"��`1ᝃJ?=����i�U��-ep��A	L�T�z���S{L5
U�M%O���<�@���?;�:
q��.%E|������f\���������FЩJ�y�����ǫt�N���L�<��|����O�z�E]����:5�F�.jI�{��Һ�9����,�/�y#���P)0��E�W4�Ї������V8��+�z�XA>���й,��Z��{��N�г7ܼ37�U!���x���C�V'��i�z5�<���hKܸl�Q��e����,��;�U����\�d�J��Ж�E,\\4\Զ�6����yE]m��)�[�HRA�Xf�P�l�3�.���ۋ�Z@Gy��e�a�TZ@^V��6���(v"3d-k�;4o"�Y.52��A`�Nȗw��w��,���X�i���vfǘ���Uג+OI^����J
�.~Orv�ѝdM�`[�HV��!}��J2��W%6�'`Ms�0���o#'L�c K�!߁�nS�XV�l��~x�U�<?8^��-7�c:�y�/���lE��7��3n�%�_q��m�ǽڍO&�l��#�=٫�7�LŬ�w�Ȱ�PL�׫5��_�|���ʵVD*��`�:#�s�^��u5����i�d��9=a{�p��H��䢔���	���pFl�����wK)�Y�&��lڢA7�31�S�-�/���-�{,q����JDU<�Z1)���^1�b��<?6��< �� �C�f��<�b<ij<��ӑ�6b�����V�ߪ��l^zG�d�̫�Q�φ@�7W^B���d)�W�$&�Q�n��ȌS �{�Hn�,��S,���_	D"gRA��BK�ﴁi`%��k�&=�c��CǗ9��:Vt�oC�Ϸր���dH��nۜ�����b|����Tag2�+�oY��b�a���a8��:�Fz���V��f��O�0�KW<�� ����x0H.�"��5��dQ?�M��@���̅8S(=�:���P��/�"�}��:߯�
U.g�_��-�b�w#+�}"/�~3���<�|�L���,|�9�oV`�o�s�@�wVtIUy�#x�T~������$0� ���ٵ��+��W��T��&�w�?�Dw�/
4c@gJК󲭎�L�&��L�/QU&�٬�&�3��a%o��p�R���T	�O4���F��畫܎���B�
��|D3�Ѯ��>?��V�*_Fx~	i��W�|BYc�0���D�uA��a�Y�H_�Lm�0&>kz'���޳C�)��q��7����Zϧ��%$__�F\�\�5�+��<�nj���)�K��;�?�X<�Vauc�Nn�\) e.y�9�,2�<�����K#�;��F_�X�8�e��s:�StV��@���j��_+�u@L ,e	��ϓZ|�
�#t��A���;4�>z��qr���͒4<8Эfj��:E2/j=$M&�Zח�Z]~��:4����P	p�1�e�C(�)6Ϣ*(�8
 �%ó���f�L�wn���AG$�ر�,Y��2�3�����<�Vg�^.�N��]�y��.A�
$Q��!E�=	ҟQ�@d^q��+ڸ��������`	K��;�8j���5�v��F �GO��ܠd�*�'�ef$���5��6D|��R��ĵ�jA�����`攧�s�	jDi�&0�F�nZ׶D�o�o�zcb�����\��z��G �<��U|{��1�ITj�A��d�Co(\�����PW9b��)VA��iT��|X̆�)�r���(�L�=��v�$
�%Fȳ�H��ӣ�k_S~��~L���1��SE,P�}��2����A��=��f���mi�8��WWV�ŀaƢY��1�dk������j�*���uG먷�?�X_�0���Z4Hn�����y�����ł+ZV��W� V����l0St��Q������GƑ�U��^���M򢔘0y�
u�^(�c����U�~%r�K����.y�ػg	p�0�+vu>0:����)�bl��+����y�2n\a\��rJ����dp������8�zn�S��W)�4��P,p�/\��T"Zŋˣ'���~�@mAIm��r��ܢ��/��P��R70Gs.�� %�:}����G�������G)V��������_���S]�-q�1mqmq��X�ַ{*,��vq���ڵ��$UhOdT̏$S���UpN;)S��m�����T�T��v��S�o��i����B���Q\}�4��_�1b?:���ͣ~�ݗg�"#���-}�y,#��{o�,;e�ti��3N�<�U�f�t{lD�� >VnO�?렢�&�Pш�����}]2�����`�G�yY��Q��[�[��/�1�W�~Ӝ�Ec�1��dǞ�bK�`�,��w�����J F}l��/kU��4��B4$P2�����O	���.�h�(� S�EO�'��ɑ_mѓtNy�r|N�����onԆ�L0�mC����(Wif_��c�sUQK	��җ�X���b�$]��xm�ɥ��E8��OO(>J@�E�H뀇�<�VsFs�}��u��H�>��Iz�T�.�ھI�+.#��R�v�ޚ�A���t��%I��,��檼�1qJ�,]!�-@B�r��tj�b#�e�+R��N������)�-|i3��[w�����f�vq� #*�t���h�H�C�<�(dƨL�G��a�B�U��?�A<�x��
;P)�*���}�=�����)y�@�sC��G@���H!�+�ѧSJv�1��t�So?BW�C|ݵN�Fr�����Է�D���	�}E��1���IL����wL.�MU�W�O+������}>�;`ZŜ
���"���&�0.#�іT �b��l]��'9o�7���Oz�'נ9�{5�#�/��^�R"g�|�ѯ���j����#A�����)��Il*��a�p���E���'|E�l�_ȧs�I7�a��G�*s[%�M(�2`2΁?`ѓ*�ʅF��`�a��p�vP����ߟ(�K�n<��&�WzW������QvC�����t,ں�6��F�Ʒ ��/�>��	�vtb��弶6F�8Hf�V�!�bS��Ƀb��UA�~�|��c�I��ɿ�vq:}��	��y|��O��e�5��sQ�g��1�"]�87x��V;Ec��)l�#�+�	}=��w�\a\:���6T�a,�����X���/,`���{�mߋ�|���:P)k�W�����J�8��d�
��3�uD���β�U��B3GT9|`��~�&��t|m��z��׎�7��l�s�Mf\z&����s�����"������qA��#tjF7Bu����i��=`�Y��څ>�����7!��Wv�ȗ�V�T�i����PI��?���O��}V9^������e?�{��#y�2(6����a͉���#���z�Wɟ7��_�:FK��Ig���vY�S�����˼�����Z�I7g��iv��+:�8ꘋ�^�Qy�w�L��N�a�n0�E�(]�&�1as� i����ל.�x%��sm<�����y2~�b�~��"(��]���k�g�2��$	��祙<�z������s��7��=�g���E�D�n k�?���~��7R�KZ�c���?��+D`�~+�+�;�U���C�2�f׿`�1B�.|�K�f�\�l�s���d�ڰt�82��`;�ā�* a�Up4q�f��4��ڴ.�v�QLg�A�a�ȫnҦ`��'h����A���������zj<��bز��|�#;�U���>�e�q��c�q��o��?���t���m���f�z����b-�Aw�_Q���i}��/}�}Tu�U���M��ִp}�M��Q����������'.�t���s9|4��\���d�J����[,G��2���r�k��"I�����#jܴ�}�����Oқ�!�ᐰ��7`���C��L-�x�u5���L�v_r��_��|o'�h��b�d�}n�n[7-�+t�/У�k�uD"\����U�88qn����:�ǥ����B�A�+�HG�&�_���m��C���d�G�����*�Sz��f�����6�Ϣ��A~��ޑC����i���H	���9�I�g6z!d���,�^B���K��2����PY��~&|�V��;���,�U����wSq�Qx�h�?����ÑG�&�AQ��e��*��;�)Jd�h�?�Rl����y�Mf� ����Ҍ�f����d��.�Dc����9<�S�h��l�C=�-��dJ_C���=�3`"CN�J�K��;�糢&o]aH�?R�dS߁��DL�%�,<:�B�^��xsb5Y��Q�-�*���v�cR��h�v�~�C;��<��ś[�ܸe/���Ly>��dzqut��J�T5�`��R�Y)�E�:�b��w����Ø�F����)d��2Hٞ-�3*��.�>��?����-��KB'�Nă��B±���(.����k��]�Ƕ�Y�`k�����k��\�~��?���
���wʧ�=Q7AU�}_c^�Z�����a�;=Z�AW}�{�V�������{�  T�`��-�HȲ���0�]f��&�+��m��	��}���|f?U��@��gll=_M�t���g�Lg�su�A�,�W}>�|aE�O� Ԅ~i`j9J�[�^羂�&��{vW\sT�q4�����ͣ��
�%i�FW�#����"6/�5�^�gb�X��]"�/��<��	��G����j�f���d��&���xB�(W�����������ŃB� �B��a�gS����O-��]�kV�2��N��.�����I�
�4���#�lV��J�8��
g�)Ld����V`�)ùó��蓂a��b憨�ԃ����2c"'�CN��}�ҩ�%�D�^1�`sݤqY�����5�G'_��I#��lb�Yt��4�7��{����w������7����H�m�Or�
��L�]�a^��PA5*��'�ХR��($��_}��UϪ����5Y���T�<��`�����2�ٜM�jtԝ/��q��+��3nR0��^�u����S7,Ԁ6���������䷣�4���^�@��{�l?�э��<�<1�V�Y�q���n�1b\�h�Gu���P���Ѳ�����OC/��0���a��M�@t]}Thp��q����8 �oNj	�E�>~����v��)n>�w��l�#f��������o�pȊ�n���� S�O)��0�Q�e��j�n�bT_Td��N,{�D+ucd��/�8_�y�'���릸��N�,���+:�IEe|��zw,�aA�@/� |�d����7�aW��N�9!l����4�w�`N����bI�'ڻ\V�T^�9��El�:���7����DGyAI~���]d% ���-J�eO�d[`Yd��~x4q��1+����V|��I"�����seya����T�Rg��P��h��4/Ԏt�x�j����[w צ����9 �ٍ�5�r�D���I�D�$̸�ܖ�1���1g6͓��8�lL	k�Rj/�����B�d� b���)NWP8(>�H8k���(4Gx5|�d���q�8�w�S3�w [����pL���	�ްF�f�8� �Dk_����N=�f��!��(��
m�OY�����dW��d��v7�ZRV+_f<򷗿P$Z���PK��ЫW�C�K8�4+��r�qlc��/#:7�i�����O,�9�j[m��=��|	��m�o��̛9f��V���fg�ڌlSҀ8�ܹ��׃V�a��}�'&U	�{��@��H=�����#�A�v�쁆і�HR6�����,���/��*���"p_qd{9��+�SkV�ßo2��$"��&E��F�� E�Ս�y��CL1�0�V�ޜ�Ta��IX�/&_X#ƪjH���6��X��� dx�ѻY)u�F�79�Q���+�I�"���9��a��}�6�'a"<㉊�L�� �2�߻ϝ�9T��6_!K�>��jҬ����q�'�?u֧�i���"z5�f��kJ�nAm�k�L��G��8E���,Bas����e�pEC(Ɖ�Ɯ�s<��4�{as�Ǥ��Y>�&�����(�֦h�2d`v�������3�+�m�G��y�Hb���o��)��]��I�������8�{��"9Y,�qǟ�9I���Y�t�m$����!o ��7�x�AP�'?�W���N���B��d��mw�� 9Ȼ��9ǰ���W�G�j!(U����=��9"���'.�R�Z+��H�)WŕZC���y;�dgT&��ʈ�9�9D��!�m������{-w����_�aO[���|+���\��% �v�+���1��6��P��w%%�.i����E�9����xI��-�<�.�A*"����$�.��4�=�� �����b��B�$s!Da�	���kUoPE��ߜ�K�4'����b���Y}�����dy�����\�����eH���4�ܠ��
�#WoC��#��V�3��a�Zj���O����خ�?��e���w����g����&�<y�����
�� h�i +.
]n$�
j��aF3d&�
*�~s�'X��G�A(Rz�Ѿ9cV1�]��
��p���)ߋ�2J���QK�'
�ݬ,\�����R��i�x����ҦO�U	/���~#���j��
MlLY"a�j�y�b𠲞�u�p�=�b�d�����ݟ��r;�b�t;��[Jz���Gz-9����e���2rMf��î�e��G�X���3�eR�Ԟ�7�V�����J@�σ�	��L*]�>�F�.�k4��ii�yR���t�}i#����-Ř� !��hb{E�<����1��]��"�@�b���r�ޢ��(����V �� ��<�����o��sgp�݋�ho���>E�e��5��3-���"��h=<�J\G�Q���﯑A��!]M!Q�s� ��������AȦ,��X,ë�"�~2�:��a>f�ng�q3��Wf,��m�����!�"r¸������lE�/��S�+������eN7�B��y��5�t�r#��P�}���d5jk�'��s�hl[��j�M�>�_�g*�kF)����9R����.��(�^���ex�`�~~�mÎEky�A�*�S���+�"\����Ky('��ÀT�ϊo�f�T������u�vY*v�(�S�*Zp�h���ҩ�L}��B�U�Z���b��XI���ܷ���r-ݻb�Hr����g��.{��	����N}a�V�;�x��u�6�u-Pn��w�Z��uu�M����)`bp�a�ħ��8u}2�W�F��a�lL�Ia'�Z{�����ֶ��0���ޅ��S��a�1&��ڴ�>I�;}�D���}�"SΑ�Ν���ܟ�O/]R��l����x����F|� σ`�����VƬ]M��#�U��������G�]L���jo����|[��+l&���c��5C[�pq��_���{���$=+��u	�?5���sF���L���R��Q�6aj*����[���l�