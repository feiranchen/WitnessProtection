��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�6�q}�v�#����q�����֍����N!Ί*b�aW1/����9�����`��<u场�d��'$1E��>x��2liR������ k�u�؈�C� �����&�C�~�9�#|48�S�=D\�ЌW�;��w�sН��Y�;sk8�nd�W���n�Zm���(��,^(k65��W���6Q̟̆��U����LΩ�g����n<]��f
�KR�SN�e��#E�H��Vn�~�NQ������j��������"(�Ao�Ќ#3�j���'�V�T)!V�Q��}�������x��*�l[*��ݘ=�ݻ�X����� 
�uMw�]�K�:��N�f��DN���W�c�ox�MNlǡآ�&��H�m>��~�G\Y��<n�U��SiUSz���5�B2ܒ���[p�)����p�O#U#�R��8^�G���):[M��\ӥ�����0��IӍ!�T�p\ృ�*�.�]�4�f����`��s=q��� �T�8��Y��F['�3�#��4X]^��ǥ���-Z�wغ���W?U�r��=�w�	��N`�6q�ǔЈz�q�SM+i��o
��8a=7�g�w�B������gtk��5bd:��K=>'?S�t7|�Sd^��n��h�O�Op�:�d6��)^קbiT�`%�}җs�w?=��z�ΐ@M
cX@7�����t�Q׀Fe6�T�<��-v�uEb��ߚ���f�f4��8	���y;���R<z)�i�W;�����goʾj@�H�T�8�$TyBw� �߫�*�9]t!�n���N� �Z�Ekb|O��쏒/�?}0�e�A��eߍ��6E-�k>�������2�����b8���+��e	h�w�M��Y���9����j$Տ�q=�г�@�m<^��]�ZRȻ<&��E��6��ڦ�c&
F+>17Y}�{����r���'�*Al�]����".�*>��vݙE-]����/�ǈ��pN������%`M&���D^���*W��4��������P�[�r��#�{S����jI��B��7m��eZ��|��KLe�(���M���rW��������u�$�k����Ѵ�; ��=0fG��%�ё�@A|'�_�p6��9}��8�W���Y
��&:��oK��h�
ū役�����Ĭ�zgM��j��:�� nu�Uvµ�8����DU����ϖG�<�$?,��>{��-��bw��(��V�����ߑKp���\nax����PR2f&?[�!58<�>����%g῝�RX�5i\��C��Aơ<bAǥm����|�̓��5��D�s�K���~���ݽZ�_�ŉ�L�r`e&�[z��S�]]��o/K��<��q9�c�$�ѮpE�y5p7���Y��X��p��p^-ЧhK�, }��s��Y�����I����&�x\Y�����+��^�;<��'�6��,�*W��y+u�����9#��D������,��M��G�HKJ(�����<;���p
)c ���T�)f��|���S�W@�z"����:�跂͸��'P�h�{��$	Z����������!��MO�h�2xi-m��Y0_q�IX�e�� � ·������ل�,'g��<�8�C|&���<��y�b��65����t��0���Ѫ0ژt�x%w��Yf��-�aXt���`t�_�g�0(v�X}�:.'�R�M���N(�]�SF�I�v<N�L(y[�t0�1�@�\f���҇���ޢ��֞����l�w}�V����w`�s\����
��s��~��g`�bw���o�r�k�;4妶~a�����B��;��t��r�+u��b��v�h*5�)0��pu�Q����P];�j���I�^%e�4|��N�ֲ1�
��l�϶|ύ
�*rB!�	����\��ۉ�@Jw�����y�D����x6*�\$�m�Z�LG��T؟P���_<&��o
T��`�H��.��e�9�����j�?g�CI=�K	2z����r8̺/34��J\�ܚM��f(�/G�?ƭ����o�������4��� L^ȡ��\PN�l#��ou�D�C�+[�?��
�2�dX�iT�� ݃K���1�l�Y�-��S;"��r�ڇW!�qQ�Ѧ}FʕJ#��@wL�uf����̥^p���|D������		�B�7�STB(I@������B&����7��pG_���&Xj�C��0^(֜�d��q,�2���e80J������6�ij��"8��p^J8]`�^}���c���w�4 V�����.�cO��
f&׮uyK�=X�)���ok�u��Ę5����
RO�� ��]D) k�{�ە�PJ�y^b����ݲz�3�В��9>��?�Z8�.b2y��_�Z��0��iQvWgXx�}��E�(-z��k�� v]eѵ�$k��<�v��3��/���i�L:��(-��3[�n�a�UTu�uEQv4��=��;(L�EY����W�lO�g�d�d���+����� ��s垠>7�Rbd?Jҿ}2��{�����tl�������~�Ϙ��Ek+1���e���$�x�����ff�zK�� qK��R�N��!�<�G����/4�$X`2Zȩ�\Z�X/�_��&ܐ�<΅��j)v�ԁf�W)�W�V%Z�3O�S�}�	Դ�������ns;~O��:���9�h��3Kdv��PlvvVN'O}$����KoS��F�����|�&������
�s���(-��}��1�Cq>�Up>v�1�/5�\��ֲ'�i�Y9;����
p̱�� �ɭ�aJ6�D~Bܼ_��u�q6�
�&��zՙ�H &n��y��T*�_���V2���e���Zĵ�?�����;<2�V�����.�P��g�4ڱU���˴�MP6�?�{d2�܍��}���Q"��d��_��I3zz�����x�V�3D��e���O���JN��2�&��;�HvW�TLi��
Dm�(��z�Oڐ��t-5H���-󁔲��LQԵ�&Ip=<nG�7�}8>8�/�A�L�~�2�F��r�PC�sI�#枺����=�U`[�؉P���R<��8�\.�=v��K (}8�cR��I!�	u+_<S��'�B�� ��!���\铛�3�6q��8����4hw�LĬ��]��g���o ��VH OT��m��Qt�(;�܀3���g��c��J�7'���B�]>�%ͧ�>��z�B�����u�R{>>�'�n�<�P�;��c��>M�
�9�D�#�?M2W5|����G�'RǊS2*���ɯT4p�PI��6��%[�� 0b�3*�4����ֲ@3�`�Q>�^(��¹9�#�!`�{倜ʁ[׾��oOOf��Q2ݩ*�[�*�����͍mW��H��l�"9O�`q$�w�V��/'�2��-���5���?E5
?�v!1�0G޸��/\�J���L8�cꘂ��KN�R��+eWjŨ��(3?�/����p(Q k�_F��*���S���8-�[:�'�����R��!4��K���d�}�}��}���'0�:s����^��+������3g4Ȼ1tFC���6�[Sr�)�l5|f���Ֆ@r
پ\p�ߩ��W�)K�.�̂5��l~-C�0��C#�J��Z@^A/�&��k��7���\�y�f���٢��+�wT��c�C�e��E�s3�����Z\�x��d��.��u�o�Si{1�Lk	tV���B��9? �����՟.ҳ��F���lȋ�t�i���I;�h�������NX��x��;ԣp�tr?9���q!gV�����#���zq��]�C�By���.	�x�g?�ץ�����ʧⶇx��4T6�c�o�{4DZ^(p1�<��t���\�{�{b6����-�i(�-�[2�o��%��˹�6�_O9�5B� �h�Y�d���K���}��-寗�F�)5��|��?zx<FQB<��K�ᜣ��5q"݁L����Z�U���T4+qBCg� }C�n��*:p�*�j�X!�R�4���>�UȚEZ�4Ⱦ��@� �M�Y���3m��"�d��L�9*v������{�7o�8��Yy�Yy@��>���v�%C��x�L���H�].��1�&���*��fe�
�ת{Ȫ1߃x��g�*WE�� ��8��yu�7evP���
	Xd\���3#(�*��\�$��d&˰ G*(?�{Q88r���v��;\���p�m�p�"�I��?�R��.���6�=�o?�3۔�!t��VxQ�� j9��a� �@��i���&��T9���yJ��߾�mKY]��J9+�=����u]�60M�����㊯��96�<��*10}ׇD����yOJ^S3�u{�gM(C��5��i���j��d�t�U8b���
�c�v7<�L:ށz]+�P%�eJ�'#�3����#��2_|%Q �r�I9!+WlO�3C��w�4����������$A@nV���t �E���E�� ����F@�<�jM4^�]S�6dĭ��o�vG�ź ���5tԸ|aXC��c46}���0TA���s��vν3{fk9�����C����?Y���.���1l~�QH�H"�!P�[�ȁ�w��R��?�0��J5��Tx?̡6P<禿�DV���r�jK�해�c�/�z�~�E�&�Y��=�M���R?*��8�h������$�? ��ʹ��.�/���7(��Y�#�n3j嗹+Ҿ����8 �껷�8w�=K��%��+�
���XVp����ff+"V�d�@�
�QnƮ
��0cc���_��P|50K�j��n �Fa�AYJf6ゴ@�2��"�}&,���;�<X�}
��{Ct�nl$�%CL�ѼG����v����4��!���E�g�5
�'�y��Hjn\���(��>M�y��l�5'���Wɢ[n��_3���r�`�$Uݷ��+O�(��62�9
���Y1
�oɃ��Cg�ii�F�����Nkg��m^i�l� �C'5��Z��3�g�'ʠ��,Kk790����,a�l�t�VW�0o }���鈕��A�"z>��-����!������#N����k��ko�c�~��QOg����2\ĉ�|���b����m�P�_��9���[g�Х��[�O��?F'��������&{�w�=���P�>�����x�k��?gs�x �M���֚%}k���P4"D��J���g�[NDi�0�e+A�O�n�buð�'e	�����1L�wCr�Ur�(�L�<s@C��ЮS
	r.�l���u_\�9H{s�O]��3�T=���[4e�j�d�}2�H�ʙ�@觶or�H1T�}�aȟ2}\��m.޶H�1�a�,g&�dYb���?���0��4e�EC�H|&�"�*.qu��x�@�.𠞺�g��4=��Jӱ)�7��?���q�9ͮqZW��o^W�h�c_IT7E�Yu�-�����F�Ğ�F_%��N���:�T G���M9��$����EJ2��TXj�0.d�	q�n �K<�͉���d
z.ݩ!P��+�i�p�U�:
4�1�Gf0L�a��R-��K1�f���t'��^W�ǽ)�X�ÿU�(�U���l�(�?�A��oaM���������K� ����R�P����;C�-���I����i�c{�%����N(b����N��$����ﳋ�-�f0Tg����܁!�r�z�*�,#��F>mmC�}5���m�v���(�L��8C��Ѳ{2R�SІ�����:��1�F2�s�NQ�zM6�P& �'����0�b�e*$T�?�ϐ=���1h�Jٳj�nQkS_���`��#��_�X���.�v������[�S�Wꌛ�US��;����W���.]S)�,ĥ�����($��`V ')�E�ڒď���ˎ�I�B�2�G7�
kNNP��ލ�� c��Z���"dp(�jv1���
W�Ş�V��π�{��ŋ&��o�D��2�8꾮���쉺�����W��Ly�,D��Cz�¿�핲�t߁�~Uh��q�i��Xqъ����B�W�ed�c31�����%W��'���S^��i{���@�sר�v6����U b8y-���pI_YZ��7�h��54+��v���!=v��A��W#�`J�}���{�吏�Q'�n:"�� ��|X� �O��I��<1q9E�6��"cD��Mq8��wW��G(*�e���Lw�W��\j��8��8`�)�-��4�5$��av���n��sy^2Q�Qk��W�P1��j�-�ڪ�K|�!� �K�ٓ�u"����;��2I���.�@��{^:+Mq��YUC�
&2�Z]��)l	P�p�i�+����-qg������j*dZ��)pޅ�����Ѥ�	�-�����ɡ��09YGjEQfS�G�D��`P�I��J�#�����5��Ъ2�%Gh�K���,�
(����멎�������<{H�MG!����#J�\�h��8��ǐ�sVÎ̒VO+�簵�I[�%���������
Q@��Ć|&G`��í"lDB��4R��E��T;�N	1�_]?7�ݰ��=�s�^�_��9�E��5G�����Ǭs���F�
�Lȝ#�����:���Q"�e��*�#��
��a�(j��n.�]�X�)�Ao��q:��c2Q�W��fk]s����O����5�A~ؿKe:�A�J�U�8�+G5!q����sQs~�{�f!]Q/j��a�e����+�˥|0�l!R�
��X�.�(�l6:
��da5�Vqw�Nև�D�T��'���Z#i�Z�� �k?HAf�疶��6����9E��	C/a��)�k�O��u�o[(��\3��ź���'��C����>�x�t��+b�pi1�FF:L$��v�SO�y�7*�Z
WRw��������w�+�G���\	e�lÜ���i;�'��c�k$����)�5��e�r��	��Q�=ƣ�����|9G�"����5?����0��v�[`ԏ53�ڗ�"3V`�o� �Fցi%踏�Us(\�jY���4t$�����ȁ4�`Y@�G�'�N���LM�vC%L��E�bt���z�G���rɯ������O:�]Q|i����ϱ��eB� �XEcjo=l���V�UA��-�}��;��H�O���g�#� R��6WÕ��y��O�{;c�f�egΫ�x�&�\��w��d���[���S��Crt�~L����Kwrui�'��O����U���c�O�/�s^�ȶB)�2Cv^��$�양���r{�n��1Ә:�a̾����a#��It6���&hX��D�^��>ԝs!	�����H�����&���H�4d�ɫ�>�KÜiQ��N�1VJ�#��X��s絿U(1�ƻj������|��h�3��P��"6�D�+���*0�C��N1rf�j�
,��y��(��$e:��;�M��@����N���,��j�N�ma_�����{�P�)s�#y� �2Y�M���)��F�I�,��= \�W�����p�x,�	}8A�Br�uOӅ�[�dNdc�g񋍟9�-D�%4Tfި�����`�a���x�C��o(�x��8�P<�� g�
�"�8"!s�1]"�Q&����d��2��[k���Vs_�����^>�������0������C���{�+s�c��y;���Mc�%�pZBy�%:Q:�1<�7�v��ن����,���G��Z��x|��*,<�;9���ܡ%�����Kx�hP=w���p��h��$����/��Md[Ԙ`��Е=	i�KfF�Z#5����Ȣz럝�ʨr��`A�Nؠ���֌����4���2	j-eB~����Vϗ����h�kͽ�7�o�<��5���E����ZK�A��3`���8����'����>�L,`�