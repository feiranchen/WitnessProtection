��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��4#5��
I��q��7�y�J���K|.ׁ���	����f���|P��q6�c˷(+n�C2�&�=[惢��3zI�aΖ,,���� ���Zy�Y:�$^H�% �s1�=)E�9yj��7F��t.G���,=���؃Awޥ�j(>�G�W�w�*�\� �^+I��.����_|7(��y�S���DW5g��M�Lu�L؂�j���ED��rF� ��n^���b����!�4о�8�`�����i^̅���`�T��@nh��' $��j�Ց:!�%hRL�����'[T�b�z2��w�ĉ����D��� 6�'����ny�^i�=g`B
������Ҋ�@�s��F�Z:P�f^n�#���x���4�t�Z�F��.�F�o��0�ʾ�n���:�k�Q;��ϻr��l)�P���œ�<�eN���$�(�GH0�� M��hՂђ�h_y6���/f��Rذb3�Y����c���2��%%(fk��A�	~yS���E��h_T�b�̲*=���x���v4�'x"ڹ�K�aL�1'���c��5�ے�`��o��{���ے��Xr�k�*�*�(�m����w�c�[[$�B��jC��LK.���N��b?ҕkK?
���L/��
�vq���̵8Cl�<����ڌ���}Ȣ���uB5{ Ej��PO���&��,t�,D���C��Z���iu���=�����-+��&��[J�ⵁ�<��� ��m������=2���;.��CKY���=��,`�4�����"�(E�h	GI� �xJכwo����. ��t���E�Z��Y����Ye�s�5��)� ����>RO1O�L�u�7Uo�~���j{��x:�
�x�I
�b�%u?��l;�3'�q]�#룰/���گ95{�����{Yq[a�Q� E�w_w\��i Z=7�Y����)��i�h�վ`�RB����5\܈���v�d;�i��-GI���\;-�Ujƥe���#�e|��A{�ROɱ��X�1���;�3g�0� >�L?j��@�@�a�2�p�(��]���B�z�wɻhC ���'�c��s�ٮf���,���N)o~��SU���P�(j`�҇xx)EmW���s�]NWsV~�e<�k�B��Ȼy`�.�!xD��<����ɕ��e�k�(��5�N��h�Q
��y���%)�7��FQ�40?���.�����Ub�`B��q"�l	/˴h�P�,]<I����d�& �'��*�;!��Ew �Ÿ���,����|�(�w
Q�JYW�^7��ԑZ��"�>+�t/��`�����(��AնM�LHZ�:~�������s�����Q#n����r,�������D0��׻ F P2X�4�K|�7�ޒ��H�?����n�w�]��B�|e-z{�$�~Q9v��F���F�.<��rsSЭr�#ށ�d=�kqc$ӌ}�d����Ս�|@}%�#��U�&��:�}d@A�����&r^	����X�uX�k��,�c^��RD�1握Oֽ������9v��Eqw�t��H�vR�H4�]~�lӋ�%C
gL���|�l�n��o�7>U�D��z�$��j|)��xeH� �>u��TB�&Ѥ����Q���JQv�- L�q�7A|��p�rm��'��l��������\��]�+٬�{p���|�ӂ���@�
<��H����L����ЬI�>��'x/�/@����A����C�|�Uʼ�|'�L��jm�9�{R&����@�,�Oܪ�v��pLe.PU�C�{ף��	���ڬ?ј�;�mTև��\�{�.^��Pw��m&�q�%�3��&ep&z�!{A�uYRóp,f'��ܠ�]�K$@�i�P�/��P,�������)h���F6�`轶�6V�t���XÇߨ��Oy�r�
/]),��3wqq~�rt����TӰb�TOYB�m֯��.d��z=���J��7N�vYy�M�㘴e�^����R+�KM^�Q�U^K2��| ��/-5������$�|����T����/����:ep���챙���w�hOu������܆I�3H�qj�Y"\�'h,��v��h�L,� f�<�4���w�SԱ��2�U���,̎.RG+����Sbui;	ED��;}�����7����iG`�A��H�E'xܺ2��C/�ԣ>AOOb�W������wGB`<"}������'Un�E8�/At���}�ܲ�5�D��`�ڑ�X�G,�Z�L�gH~��t���wV�۶�3T�B���K��E�G�YF�fx<����>0�k���qx����c���y[d��q�_�s��!��hAJw(�vk�m&aj���&���=:��i�մd������0��?>o��q��N�MF0��y=<���=׋.�y9���p� �`�qt�L�\P����"�G9�����f����c��>�k`f��z7L�{���98��?O�l����㹎���ۇ�gd�߅��K�!��N�W���JzW>�g������򁼕����8Y�Dף��J�e�q�q��^Kd6�TU��Uk���as�'p ��,�̆���z�x	/�>��8�G+��ɱT��t�?�T��u!��2��a�J�o4%? �U*��m7�-�bzj>wk�I�l! �ǋ��E���Ƴv93��EY��=R�c*oÇ5����e�Ly^L���jR?�=D�2�Dy)��:�}>^h#�<��A/��Kz��.��0Ghѭ&S�PL��x2��>�K������*�>�l��;���z`Y�G5�8��Ȑ��f�܌�u}�\�4߿���<~I�sx-G�M��Q�`7��;d 2x�Lnw"P���Ox	Ip��@�|��υ,P'!��˯���ڹ��jA�|>�ٕ�!�b��Zal�T���TK�R�\�s�0o��%	��&�()�����<��-���y��k2X��$�J	��trD���W�`����6X�`$�~Е��΅�Y���a�-Y@1[��N�w�����2�0�8.���q�5x�d�=A��2?��\��cD?�SO��� *�K�#��}wIhf�r.\�۬ X�^:�(aj��_)`2T�X3�f��!?M��v�ߜ	_��a։V�؃��wfl�"���yc� I.�b^v'�5����B�"5[��V������#��<45�+��	�8���\1hV�ucg�w*2d�J�U��)9_vN��3�k֌8*��Дt�JAt|D�����H�����@�n�j��Z��f����5Y�	���a��C�᠈s�Ң;�����-�Ve
�ɲv��&/�f��>���� 6���$�Ю�w�K�AЇc�r�'�rBk�{Ӆ%�~g�H�y��]ߪ:3R��1�75��ǌ��&��,ڡH�)��uY��rX���Xn�'�i��?�ݱ���xF�~�0	���^D�B*���",Z]&��8���2~�e�T|�@ԉc-��mtZ����,z=b�җ�������O�)��~y���zp��{�0���&R��6�tx��Dg��\�u�7Mu*�i�͒�Ј�
�79�C�&���UM�Z�"�1�h�����ؔY�~j������9�*��NYS�P_Z���-9@H40_�1Ω�er�p[xW��`pO��'���z�X�@0�{�z�1�cэ�!B��X�$
���y;$����Si�9{Ⱦ�D!imm��4^8��i{��U��EA'�Qͽ>�6�/x&������im��wy!�U�6��p��7�e�U�Y|��C�h��	$V�������O��_0Kxb�� w�ҽ�,!�y��<sA����[��|��C�@;q��A�8'9�Q+塰�����c�4��ױ��aϸ�u����m�b�W�!�<�P��;`jQ~�����/��l��2U^�Z���56�zi�!�k$c�[�t�1�gݭe��VN]��	Hg���"?��)]���=;[�c���)��k$}�'�I�9
��[�IV��}��=���^�9��)�̹f��ٷ�;�MC���Z����0�"�)�Ma�7�{��T����v��.���I�*9��%�`{t�qTΉW�B��Xg�a3J$��/ȸ��X�NO,�4�,*{7�V�ޚ�6���*|�fے�@%޿�\����F%qb2�D��|ݥ�{�"��c��ŮiM/�߆bV}�L�5X�s�mR�fV����|]K
Y�)p�F�� ]L(^AY8J'=|`b�<�c�J�L8���6s�T��/VMӝ��O�,����^(��8Nސ�:��tj����dL �;K����1��qy,t����)p���<����&����l(� ��ԙg�OD�JYb�6����A�N�M���X�uڮ-nH�2��6�>��ǦivZͳ�Y6ѐ|Ŷܠ���V�RR�ǀ�T⟩�X�ͣP;���D�˩ �L��'��b1�5�kV�)��VƘB��:��Gy�h��j�K���������
l � C�� zn×�B��E@,Na�Q�-B�	��+7����$�eyՖ=��c.+9��`.>
����. ����_@�`�Ovs5�1���60(eO��Y����j��˾6$b��$�,.��q���ܑI���h1nVc0�!4��0�,��a`��.����<L��#�|:k�,��������"��J=��|���UʡeÌ6K�顩�>�&x-7O�mhz$s�ڭ��#�5I@�\p� ̪�0P�a��x\ڙ��LOYq0bAߧ?>�^8���D���Ĺ�U���
_KO  
����O��d��=Z~^Pz.#�`�V=�y�Y(zL�������̊Ց�pz��2�|sF9�DT�y�i<�_��8C��k��5�c'��>�uT�{��˙���2-��dx��3	ژ��y����*�D֚�`\���aFIN��n��Ǥ��5BԴc�Orr�����l����ً�P�l3e^[�Z���ڮ";ٝ��4�OR�� ������%��ŋH��.$�.EL��]�/�o
�<��OȪ�$�-�$Z���Q��Ⱈ�N�;�?�q68_��B�e��.K.��*=�8W�l��e� #�n��s-[t��q������:' �K�u��m�7e{�TO 8�"�[�0���6�M� ��'���������V�=4x�.�]�m8h�=����/��X(��z�ȉ�X��:�Wy�#*���:$��})�L� xA޾= ���7�]�V�N�!��N ���1d�����;�D�23��w��{2��=_o�� Fֳ�$�ݨ��s-n�(1,�N)3!�j}��g$��Sn݃�]�
��^��Z��n�B�c�D;�J�H"��
q�`Ӥ+�06�/���s��ߤt��s�����XPJ��a?��$9�Q�H�
��=�>o\�G^�)�u��=��.���#���#�"���ǚ�A�9���h�8��d�{#nE7O��\ɶ����0��[���mkP���l��N�.�gq�D�~�ᤄ(s�q����$Aw����7p�M��P�y\���*���,����J'������~l�L����qM�_N���y��^��Xr�Z��a���pOg����4gǱ�69w�a2����L����n"J?���������G�-A>��j�ō#�p�!u���c�VfQ��'Y�)r�!��HE�l��5)��\5�YJ2#k���M������J�L�T�y��'�}����i� GN>�Em��ޯ�Mzg�,���$CRB�T��֣_$N��4ҡ���0�����B
%7�� ������=',���c�s�i2��F��?DUt�D�;�s��X	� ����W���&S�L���-:��d��+��9�h�L��ܬl���P�@�Bz�_[󎘂a�gJ\,PS�ݻ���b��W=rA-��&�����O2�N������ a;^��垘0���8��6x/����.���p^�����M�H��xNV����*+�xNuQ�~s��Ǫ!ΠTh@���G]?�o�=�`��Ǌj�в����ٯ����qe�S��m���K�� ��K�$t ���R����5D�;pN�*�f>��f�Ho�����ٷ�	��WG�_N�m�ز3��ʒ����F|*�%,Ш? ��� 6��S-'E�)�L����Õ��֪(<����W���X��@b���j1S����ۘ�"�I��ږk�=�$p~������[�����:��W���CE�*�s�1%4����NW£&egI#�%0F�*e�P@[J��)����n���ǰ�k�V�f����X¾_�f���Ї�{x�4�C\Y�7$U�V�k�}ңAQ��"m�y��H�9�Q���3�w�1Ǻ�`���7=�>;oW5Z�ٗ�XN��0�;��t7kO�E(j�Y�ZR�~Y_�m�C����������ڏ���h� ����XƐ�S(��5[�����khy#�x��8Y��3d|��;��� �Xl��I
��R�Lՠ�y�[x=Q�GʡL�����;�Թ��>����\��|��u!�*{?��J.\������M]�]h���ɡS�?�֧KH<�+�����`]����8��P+�P�:W�����u^�>A;���D�ϸ�%���Ǖ��)RpA*�,�8v��d������ ,������~?:qC�p^�K����L9+^B�q������!;n�3�6o}�`�2��7i��ug�e{t��aSL�o�妻�+��PM��O ���#e���QI���sf)^ކYcJ��JEa����>��pʚ���.��hG*���?ȵ�x�������e
.z�I�gCX���v	.�Jac��lk]�$3d���Τ���q��q&���\g;;�h�g�l�q�UA|R]��
N�@VzW��W9����D��r�'>�}D���h��4GZ��۬�Z�q�T"N׶Ei�����'Κ\�4	�
ԴӮ�6��沯��U�^�V�������ɰ�|�� D�ǥ���=�+)5���i3!�L�oЎD0jk����,p`�hP�����h�)�?�
Ɔ��$��7ifX"�dm������*Ӟ�{,�$2*�/����7��F���S�1�r����V�Uap���`�uf0�׭�&S�R
4�!ij�\��-�����x)m���Y�ͪ������/7���!��I)�dU�M	�~�1�R��vv ��!�ʬ�r�Ed²�e)�d�*x���5Fr-��$~�b�&��=��X�ĵi���	��U胵0Ĭ�fTcb���Z�������P`M����>1��|��6y$|-���Ҁ��U1p��`����RQ=s���w����Sf���#��y�t���*o�����B9��E���,�!|��:��mY���	cI�(��ȧ�����7��C��N���y�ˡ��2��B#�I����&sf������=�<�|��dF^e7I���+o�z���p��zoz�l���,_q�(P�����ԑ������`�Է��B�5PC��&i+�v�}�^I����� �u#�6g�i0#�N�O�w���V@k$��p��X	'A��2�5�:m)@uJ�Z@�q��ŭv��Iϕ�ۢh�ј��z4F��vq��u��;*�����bX�ц��^
��k`�Ie
޿XBӁ����vpL<�Y����C�S�'�b��t�Q��ջ$����Ƒ���:H�w.��b"'�P2V���R�	h��d�w�3�[+��&<� 	���-+-��5�A"�d��'�m���uW+����
��V����սu�R�E3l�;��R`��:��}_K
�j���|�6H|��呞����l;9{�:q��:�!�`���# �Z�)�u�o'����Qj�%aѡ�?å5����2�"c+���F���7��K?I�E���V��;n�$k���~�X�S��C�B���?��iV��"x�� p�xlT���fwtO�23+t۞�mM�JP\��a�"��ԁ��߱}U[ �Y(ʺP��O��-��ݴ�K毾��"�rF�����t�*#4�Z�_��[5����D��Iy.��V������t�l	�1�'�){8p>L���kM�*�n]�	� >���r�"��#4r*�r��pr雳[�q\0����f�j�>|�ܛ=d)��rd�n�V�6�I؏�Ş��X-���RJq���������-��v��2�3�AZ��M�Q��j(��V���u`,�e-�!Oc+��"�g&ݬ!��PF5���9��gƻ�=�-�����c����CpÝZ�}dg:sXtF;�Y���<�=P�C[:�0:0�T�	�O5k�ӿ���ҥ��DX�2�N�.pƠ��:26CyTȧ���:����,H�/X���A��.��ք5֝LS��l#+�W\=}ݯj���Ր �%��4N�Z&j4�����0=�'M�;J���Y �$�Zn�Ng���3�����`��D.�k���wF�u>^��;�8&���	��3��?Vb-�E�}|�����%�4!�����5=�u?`�{�k±uF�Z��g]Mt���pќ���'?H�[���ޖ�0G	(ӀCu��f�W���횪P�Fxn&,�ѯ*b-�������/+=U5BD�,f����[obqG%IIQ��P�U��ᎈ
�
���Um54%�=W�6P;�C��������C{X�#l?�}�����u�g�fN���a�^���b�j�3<�4�c���"4Z���v� 7�7��´]����d���A���
*��GWwe���_�]�z�lS��M���ղ�����U�������>�n���T�����HM�˔����4Vnkt��Υ,Р ��\+L�
�g�wݏ�����R�]1(>N�	�J�ȃc�<i�~|�iQ��8�K���K�{0y�$G%WS��%��_�o���Z-6Z��5�%G�6�b��+�ƨx�$�H�]�˰�#����.�U�d_�3.�򸻜.���B��=����"��0�xڜA\=ܑo�A���>��ǈ}���j�Bo"]�9'c�.}��(܍k��j �J�e�F<�~����r$_h��V���$�9F�����5�Cgr�E�@?NY�|5A���C"�a��D9����:NC�
B��u�BR�j��S����6�� ���j��:��W
��Ą�lx�}T\B�;ݨb�E�lWO�2��mx�!O��Isv����c+�q���{��n��Ž��3����ʊ,Q{ќ�֤W�:v/Z�[����v��J�!�`�d9*26��p�z	��b6�wN$��^�@�x���|%�򳽃E��2�B��tM.�hKN�C�y�!�l��J�v�(��eKa��9��U�����x���t�o'�[����ߣ(�JXrCBL%+�k?]!���=T�c�T�?�I]ۆ�N��;�6R�$��l s��d����g]���ѱ�d����5�9B*oS�x�dej6�R�a���v��Fy�M(UKx��A�t:�SƓ�Ȋ��͡ײ� F�ۡ���M�,�s$���/_�t#U���&t�Q�E������+ 8�ݴĺ�g���s��a���Nݙ��|���$�������,��{_�*�-%y���m=����х��/a哎w5��BԲ����bsI������Bo����z���~_���'~�6=����u����#�%�!��M���A�÷F�ҳj��b{���b�<��T<_����R�YV����Ѯ�'��w�"]�����[A���U6|�ip���	!u�D�T��!N!�1�;�p��i�ɓ\:���4�/���
!�y��A�Te`ĕ�¢'D�+�rcj[mdY��(��C�&׺�0���0�-�W�p߿�����E�H�ڝ��#��b"�Y�A��BG쩡f�#a��ʚ��n��z�	ˑS�]�1���C�amǓ��@���[����a,�2y�^^��������"�����&�֒ʊ?����'�Ȟr�2��ə=����:��,
P�����RGI+�]�ʫ��4�lI��}$P�e#2+%�Xyϰ��Ǝ^V���̭�0$�}��Z��2�D;FY��Kb�O\�[�zC��H��$i2W�[Ϝ��6�l�褾uvպl�["�,)�3�W_��]�3���g�E�Ld 5�U��ux��&X�5��d &A�"�%dz*�(,#̴��׸�Fv���J�;1��~u�����W�|�ǃ٬iU��ȷ��FP�!=9U_��Mx��*M|P�#^�s��۲QfJ�J�,~��?G�]f���(�� �.B��l8��f3B�I��h��:�D����"<ޓ��=Ws�?��s���|����]�G<�S�h�BA�1��$l���O>�����H�C{
��QĮ$e[�	tt�n��o����/��Gދ�Q-� ��"%7\^���߈�+�
�/�Y�ig��/��{�gX�Y��P���7��O������n0+��6�Բe���؉(Lk ��/U�+%�ub�
է;��W,[�8���I_ꢨBd TZL�����?��$x��o�!R��#�o�Ii@������s�����ʣY�yN���>1�%�q������:�A�p~�a\ĴKm�g��Yeie��B/:A�*���0���;HWԜ"tD3�<E0��8�\�.�$+�2œ��G�0��]�<]8��I�%/D��MH��`濻(Ѽ��`�Jc��*2�+�؍W1"�F;��Ɍ�Md�(�{�J9d:���G�[-����1%�f����k��ˢg}�#�x)�'{1��������j�6ԕ�?���p�yzj=N�Br@������R&4?ZUVh�5���%� �Ց��1�5w)0��Q4�r	��{X�H�)�`x�xկ�MN�-bqa#�C�c��?�	q[/��6c���u8m�O���$�oXaL�3� ~���Xq�?�!����6�b.Z&y8�6�	G$�$�+�9�Q���3'�-�&o6��'J����e#H���5��n!_�&f
�HY�G��n]O�W'�T*0h��ȾG#EP�D�I���L��c)���IHY��Pݛ��'�G�8�����@L�|[�5v��燱���j���
�mGE	pޭ/+޸�	�]\�ѡ�	!
��'l�.܍��v��xJ������� 	���А����fǥtk��BsqQ�4J�Y��(
w��= h~��T���-)N��/m�9}w�^�=4���e ������y����r�~/P��rf�r�XC�q���ך���ӡ#i�4�S��&G��;�{�1?�l(1T����)����6�"��̪���\��� ���kw��@�b͌a�j��i�j���Fl��ݶ��ʱ�u�~$%�@-�ʿ�Bj��N�W�(;Ajx�AvT0!C:�P�(��+������d�ܨ��S��!��Xǋ��o\&ٮ��j���Y�PI&t�gr>�;z�>�a�
��N����D� ���`z������I+�.	J���(�Ma��l\��KR|@��l�GA��M� ��g}Z$��&`0�5���C�Xo����0j
�//�]�aL/\��$��B�K\2Q�n�oh��֤ �RW%�z0��U�j��7.)|�i�7ʋ�^}�I�7� �c��3x��ʄ0��Wٔ�N1��=�nz�QŘ�GṂ�K�K�Pn�i�	�p��Rتp��ִ�=�/�:R��J��gq�+	�uV�~ld��A��.2�Ut~/�<�_��o7朴Cd����9P*������UZ��Rp� Syb6�@��(
�.�0�J|sK)ڀ��]ç�7��?�IGf �F}���8~s����/��y����@�B�v�x�ʖ�yޥ�m�o}!U�O���e�����$/��}�e���ˊ�]�fJ=��>�BS���'g��U�/h)���0�}����~�{Ϲ�s!�b��9��7���$���O7�ec`�@�U��ˌ��k,��5��v߁�{[jӫ5\�{���!G��H�;CR���V$�Brz�����V6�����f�c��9�Y����� êk���m��=k#�6�?�+q�jg����~A���� �f�Dϣ�:���V�D�1��K������ �rR��)J�k�9p/Z'J��������5���y�j�ɀ �w$��2:�ک F���/��y���g]ʑ�)d@<i]�_�V��s��~ƿ; �?��b���7G��p����⊅��]�n�Z���;��G ��>�闣�OE����7t���RZ�w�i&�4t$����@�Uq �EM7BP�	K}�/߷PL����?P�r��E�2���}�7�����r��I[xI������5+,��m�X�N2�����o�w����wZ��薲���h��s$MjfaE%��>��5nG�)pyY�7��~���?�[���a���1H5�����(<��&�C��uv�%�������s�d Mh�ߍܰW̗�dB������ÖITE5���R$��P��O<�t�t�Yt�Im�2Ha%�/ͭM��*7�=]ũ�Rhu�J��m��N�4������'j&_&s��$D��eKn�)y��E�����o!����AgZ�_D���C���ye/�A �ņg�ٳ�#8|�چ_V:L��nr��J�t�u�+)�|1�l�$��E���&��
�O�y{�H�X�;���`�EZ2y�6I�ϱ�&���]�e#�6��i�5T9�^�|����,�z~�i�ݔ�x�_�l������C�@�[L�U�;R�*	�:��J���H{h�ߖz=&HZ���{1�t�������R��g���*�e�?i�����81`�R�6\y���I�����;�@��\j�I1�>)�����T����e5��|BZ���K\��ו�&��v~�ԭo�cs1��n��������&>{�!Sٍ�o�;�!�IS��c�Tp.b�� �1L��r��h��Oo� jQ���J��>���I�p.���n@��ۃ7���m��tK[��+�������z"E2��~,\�.5͒XiXT�`;�=k. �jkH�h&�8�`�>+���8�p��!�nCa;׍����xdQ�qgV�;ӽe%J���P�Q@9%�[q�m�l�q;����h�iؐ�&&<y�V��5���f��
�����B�kHl8+��'P[q��E"2���>�,RŨwJ����]>@�&��\ީu�8qg�PY���I�Y��l�\�,�<�K�X��#�5x�Ơ��z�H��٘���}[sO/	�.�v2���W��[<���jH�	��[IzUO@a�@nG`�EMJ�hA��^�C0W���U6X�*��&d��L��5�ΫT��.&[��ӟf/�˓�=R���<�YN@�-8 [�v_�9	� + V�}�ޡ�y�?+|���MS\�o
������|t�Xs�8b<�(s�flI�Vw<TGL7��P�B�U^P�v�9�Q���������BD1�'(:k�^��֒�!���'��/���'�����C$��K��`�V+��="m	�t]j�V��u>����7��� �׾Xx{K���t!�;��G��bTj�9��q�wɆ��oI�2�\E4�t���D�|֣7,S&8�{�-M(�I��]�G���0�N���Ah�g�.=���Tt���Kw�׵`߱�|��Kvw��Z�>�n��IҪ3%��Zw_L����ĭt��9�N�6�P����p�L'��B��njM�Tq�Dh��2�Ի)\Y^��*�Y|/��_��*4�+[���U���h����\t���OS���[�u�q�_�w'cW`�����.�Eyj����3�~��aq�~�۟iIU�3w�Ѻ?3���k��[��#�P����b�F�"��]��} ��W^�G��x��{ql�a�}TRx
W�MLM KE7���Ws��V^(���0��i��8��X<�d9�jp[�u5�������w�"���<p��.����U.�����_�A��$�F�����"1�5�9A�qṅ�S�\R����^�7� �0��F�<���	�/����7�*�I>Z�����QDɔ"�ӓ�Љ�s�����;Ռ�T��T��Rb�Pe":�������9s�9�8��C��!�������r` EI�$��?����nY��Ĥ�
��I��H\��H5�@ٛ�=���+��'�L���P=@-�r7�۪��V^Vݤ����RArM%��!k��m��_�1��]�E��F����~*M�mZ�8y1�D�#)�
��)�˩%@j��l4����R��D��`:g.�^�v���HP�f�m�\ϳ�hգ�)'g���/b��
s��xB��{Uϊޙo]��+��1D-&�j�^��X���7��w7$ȟ�b�ٳ��@���'�`6�9����S���>o�#Y!����FF�=( 7�bK�L	�2��o��(5��["����3{�R:d����j�{|9+��M�&���l_�N�6�y��X���I���/x]ܐ� ݊�1r{�W���^:C�  ZN �g}֧�	��cIn�jGz�k �ӟr5��X��� ;�����`�_gbb��=�=� ���[�+����;��$,Y�y���IbL�z_ŗ|� �����g���w�IA���D��@J��_�^��2*�i��n^Q�]��<;�o*����h����gN��+ND�W�-"#�l3�jRWb�� �ی>T�X������{����`T&-�:��t}K~е�M�MY\�͋�jd̬-�+���Ӳ�{��A����,�@�:^�B��k��B�*�6;��F��,��	E��O`¢�I�=�r8<	6�i?j�E��Y��0�e���Q�5��q��P�N�̪����U"��J�f��3l`�\���@@�Di���A#1<�]w�@�7-\ZmV��5e�D����&Ǖ�+�g���[��s��	Z���eD}l}���q$V�toF+k�� K�����?�)�&�w:=%�R�4�cs��v�S~��LXl��0�)e�+�|Yګ�HdC�'=��e2�v'%K�o�{M��s����#!CY3���pk����M���>�^�2βv��l��GfJ|z5h:󨠻c�BfC)<�m�JH�b©��M#&�Ź�+��c�2�qf��6[x��~��C��Һ��j�~hanxO[��Z�W��TJrl��_ր��ċh.��j���ٕ��*����!��i�`�(�d��T�ْ^�l�Z.#�H��h�~Ў��YP����N#8�[.!:~=O�l����u�1�↨�jޤ[��Ӣ�GSqNje_@Rkh\}P��)��z��ι�:ɲA�)�����Qw���O� ǆ��Z��?�m���L諀>򩈃5��j�aܷx��(�%nh��zY>�׭J�M�Ɂi���-��Ū�H:t��~z��U(��&�F�{%*�Ƒ�L�
�����*[V�켂"`/�b��g�}@�0�:6@t�J+��+��i&<�h�)�'#�r�xP==3��qȑu�E�����Q��u'���
�3n���.~PV���6~��jS�����F��g9�ZM�te$� ��j+q��K��-�p6��X*�x/"6Gd����(�=�z���3�L,I&<�%%кKK�ߖ�ȵ��o�"+؊�γ4po{���f�ڰ�L��ڌ�a��aZ����2Q�
��WupC|�L4Xis���6K���\�b׃M�C�d6��l�l"��� "C0#�@Y�b6Cjh��v�u y9݂e��V�P�i��UM���:;�J�B�o��^�Ҳ6�җ�.ȵM,W�ER���2��]��Rre��}f��7Gߘ��K9��g�~$�o��Ze�K� Mu�`���~�Y�ֶq۲� N�1���ڨ�Q��Y�S_��ːʜ��{�d�����P�dV�)p��
����%�נ�S�|�K��Rh�47�x���M�c9�n`p$��Te���S"j�@lql��n�D(����}w_,�(���V�Զ���0�Csf~����r�-�I�.��@�LI��Ps�jq���b�����|݂�h�x.��~��j�X�{�#XS�$�p��`���3N���b�#1�թN�i���F�!/-#�
I����7>�����2c�p�j�C��-�?9O����p$��o��r���_O�.�M�kk�r��KL����Y�=/�D:�[�a6��}��$S�A��Up��;���z���T��E�_П��,hz&Ѻ7@w����G�u���#�m q02��=}�'�	A���/�`aFP���O�6/C+�AY�� y�|�`�7xP	SpQje�"�Ǥ��+
A��Iz�+Q��X���*&�t¹ܑN��)dL:]�C�a[6�����w)EB�H���-��g�<ۃ�6��"P��\�LI�	0#���Ġ�nJ�3Ry�&�D:�hD�KEh#����JL�����vO�I���Q4� ;u�^��
$��12����7�¼�Կ����|�H[���-��?�e�`�4��EM��;=�-��:�c�e��x�DCq�L�ۮWF\_&��emC�ze{!=��:_K]p�ݎu��W�z|Vp �<Z�R�&$�6��!� A�ɛ�=j�-w�~�Jå�1�����.#��!7�&����AfE�5b@��cPa)�U�#>�V��
H0,q�÷��8��]�[boAm�K���i�EZ�TXy��r�G弍�ށ��'�sߞ?��z���|�����Ng���`0�y�q"?#'�ӂ୒ ��h���D�w�4����Ԅ�xX~0]<�i^�����1��QU�7���*Z<t���'Q�*����62ĝ�p�-lHT�'Mt<�����7U�?��dƅ�>p�'�`��_���5�E����ԂOY�/�R���C9#�a=�]���2~'m`z�@8�sw�Iñ	Qlk�U�\w�+��wޒ��L[4Ya���'�2 X����tQ��c�{���c~����l��q����A'qw�����S���pfnĴ_g���٘7hV�,�\9l1��6	�� ^����_�9��1d��)�����qUm�wҗ< ��x��� u�"�ں߄�@�]�@iq�D�T�!$�e;G��ĝ9�/�W��v�����lj�bR	-���Sj�U�Oܙ�����OD��j�h��]����S�s߱��]�����^�['~���v���lm�ո�1*�ڌ��_HE��Zx�GCh*�0�M����W�:i��d�u8�T�A�Sx�Qסa'g]>m/Aү8�m���"�&���8CF��F8g;T�Pk?fcB�W�I����PU�+�	�Fi��ݗ6����-��_�"S��F	XM�=��lʒ�g���Ix�V6�����S�J� 	)'�"���Sۊ3p��^�	�V�:(ЭI�����f�ؗ��W�;In����"����|�|%�Z����֥ �ow����al��"=e{H �>ᾞ�c���/	jK�c_E}n\t�3N{�WOe��]}��ꌄ�=���Dy�i�����D�����a��`09��.�~th[�rxK2��
;7� A1��8e$gF����_��1D훹��)�*��a�j>��W���G�n��yPB([�D��l�"X@�@�x>��Q�T�g�1Ms��c"�S�4c�Fw�B����t��0!kbPR\"�ki@����e����)G��L����6��|��C�;U�ɓ�`g�A�Vm󧾧�1D���۱t}�����ڏ��m�.N-5��D�>�d>����qY3��(�y=+��'s��0�yu���()���<�vTh�䫅��$�j����B�PZG䚆�P$���]��죯@����gr�ӯ��.Ms�	 ��SH}�s�7��lmB$��%Ŵ�h��X�\��_2L\hc�wO�Qf���0��/�E��g7��8����b�G���_�*��춡����)���g4s(({��!��EE�=�N��nL]
sC�B���l�`$��s3��B��0�
鐬9��<�#{Mҵ2ĩ��I��/PYw�S�35M
"걐槎-�o.y�v��'����T�"�VE�У�W�P7�Y&��J$]ʪ-��4�L�l_+2~Y��T��X�p�k��	�t�F,�o�98@�'孑}���9��K����/�"VQ�av�k�k�8������	������!]�1���Q���Kıa�G��M@�����%~3!a'T��"����G��h7(D���b'1B��j��[�gH�z���E=M�ְ�č�D�~h��o�C��+�d��̢��pWu%��DN~�i�u�>�WFfm��.����"��� �/�p��T!��,��0̶[��!�8��녫?�x30��z N�<l��[x�.��L6�>�xVF���D�����=`[ᮾ5�1�,'�0-�o��0�WS�Z�c�TYW�jp�R�S�= ���q*,�&F���1��ҥ���q0{a��g/h�9{V?���u#?��Nt��j�C�z�ݡw��0�ϞlK>O0N��k��+��-��
�虫�x�D%DXE�n�&�P^�ew=�g[ӥ�q$���ryJ�7��F��o���H��:<1�+j��b߿"�����&��l����8M����䳵��@Vf����h:t�ê�{�(�]��(e�k�j���~� S�e�5�3�!c+��M-�o��l㓓� {�^5#�}Mn�0g�ea�T!n���d�٣e�K/Ë�r
K���x�V�6�Ω�0ab`:|�8����Y�Z���/V&fz���^�D�K�u8����91�By�x��k�����>���_cU�\z#.!�z
W*X$���r	�g������Uxz�G;��3�׌�M�F+�l�b7���-d����U���t#@�Z�5�RB�b��pd��H��L�+^"u>+p�#���_�x��u=N҃���˘%��(��f���\g�Y��4���m���V��=�Ƿ�I��w�>G��?� �͙D�,Ũ���]����^S��Q�\z�;
���9�dl�>-�xG=gxx�Jw�/�8�nG9����~�y��Gp)MS#yyU��:��N޸L�>u³K�4������t��M�3d@�{�>�#m>����\�/�� �Ԙڝ��g��{ȥ��K�0�$g?�����Eq� �X �h2z{7P:�S�}���qrXZY�1��n�=��_$���Y�s���6ND�I
��CkD� &���2���88��dխ��C�$z֧�Q3�<A�"g%�q��-"�U�#�(���H�q�b��d��X��ܼ��,Ԓ�K�XRc(`4� ��iu�;�Ѭ��	HaF����)�������qS�n�&��Q�'��ZcI6Ozh�aL�����0��{���;���爰9Ai��B��ٵF��.��f���s!������_��"��o\<��b2��tq�� ��uG��PmŇ� �(=�N��������:�h���􌉲�:��#��Fi���a�rhG{f�^�c?�!�9�@B4�q/I��_ԍe�=wa�8YR&L�L��T'g�X��o�<ڹ�:�4B�?F����B��>Ċk����*z��#|2`k��!n%�@�w9���������^i�a��^pM��fsh���i�l1�b��Q�4���+���W�������w�4Rz���Ƶ�2���5hj��+:b<&pL9a�@�(�-�]�b�|��Y��c=�U��%ӿ��H��x:��Ne�;B�TK^���J��?�uB���4w�1]x�-��А����MnGZpS%�k�
��qѥDM
	���ݧ6���CN�Z�r%���-�}Gj�@5�Q�N�@�+�B��(Ժ�C8��R���?rh�u�j�D�AU��jDPo}D�IXS���s�L�v-��Z����&����@�A���_4�l��t)ll=�X�+�~i�uҺ�%Q�m��O�:z�@ˋ3�O�;�ӊ����B��si����a㺑S�g������;�9NW��NuAjvX�2X�X�� �$xY��Yb�*�T��Œ��5ނ��ups�Ň��vm��K����2j]�876�������ĊQ���<� �y�����Q�%+�1Sucq��]�Z`V����pf�=�G���)�őA_����Jm�`��1����m�"��0���y�4��%]�kv��?��;7���Gw}��1��Oi]�1�}��DÞ���U(
���& �8��zȘ.JA��l@⦐��[������~5�}^�)��ΎO�:�sll�
�?7�����^�������$��/���L�ˀ�/�?��s�o�c��\N���n1O�A�Ԧ�a��ɘ5��o,2��9#Pq�"���f��"�{�I�
	Q:,-�!�	-��?=Ա�S�2$0m��[�˼[x���������FC�r]<ݧ�n�ֿr�(���>M�!�.`��f�
5� ��r��cTUd�~������r��2�']l����f�I���Os�=/�陆(z;/n�a��X�� o&��<=3��y_ߩ��	
��0�}}bRTA��[�a �2�`��ޚܝ�WWz[Y��3��3�g$�-eq�:-��6��>��./���F��öo�/�v���Rj;(��?8���kj?h�4���k�M��E�a���+je��l�:�(j��2q^�D^z\6��Zs��~�4�&���7�u�7Z�~�Ai�
G\m?Z�ԅx�vi>��d8M�1�HеY�~�*�.g(��cq|�J����)��8�	I ��<T�E�����]�O@�	2#t$ ��|�NZ�~#�oT�����гU��&�B��v�уһ��6;h����Ţ�7d�h0o�3���C��o��}V��f�%���޽��s��?�P"�*oS'��4~��"<��8K#1����c�Y�f���g�����H�ř���욮<ޙ��8�Jo�H6o���(}W�3�Ǔ_#�*p0��K�pH��T�ti���V��iͩ��*a
�T��]b}	G�0	��k)۔ķP�F���s������J?HOl�I4�����]��A��uY�+�k���a��`��|���zO���C���,��1c�P���C��KfVD�����<������Jn���c��J�cGZ�'dn�$�>ۤ[k���˴���S��Z�Cy�?1�kn`�L��͟�c%'�����5Vp�
��˵�Fu火A��������h�,�T�p����t��6>�ll��ƹ�t�tlv,�	�q�M�>�*���A�k�@fY>J\pt��{�s3ױ�c�ӗɋ'�!%Չ��+�b5���v l�cQ7�V0�:���S�D	6է��m�V���ZDs�h��]ew��R�B��r�%�&B�7"e!ުcGQ�._�ta؃��  �B��O.ZrX+�Y>g\Z߈�F��_�t��LS����jF�<��Y�i���-r<��Z��g��Я/��du����¿Zb!N��2�;U�4��_P�a�T��)NQ#�YUf�/k6_��w>�<lb$U�9=���!�M��y������U�#è�j�1m��dn�D�^F�%��\
Tn�±|�,2�)u�Nx�T���h�zH��B��O�"jK"!a̒��PP��0�=PRZ��K�f_�r�2aX�)_-��#�X
8l|��̬��{:f��Mm`&�ӷi�_C��O�˙4n;ç�|&�jGOG�56H�R���3�9nE��.�ETm�<1����"�a�kl�M2�������A.-Ŧ$6L�a�v�O�H{�q��~��Z%�PDn����h缅�E�v�j&V��g1��U,l���0.�^9v��ԉ'9�5<F�4�� {r�U��?z�M�3;�r���������Bpbm}������- .���<�9G���m^�#�V�{�Ǡ.�f+�gR�I5����*D�!�[�?����6�_0��S�"��c�<�����4�ekD�'<��W~!�x�J�NmI椫i<��l���^h7T����[xm �>Y�b`���j����Kj�����R� �<@G�2�GH8l��%ʐF�r�E?��NY�����w�c�;D����1y�L��R=PS�޺�z��H�f����P'*���bKiw"4�5�������a&q�S/I���B�z�ju���Hu�ݎc��������>��'��Ic�����^��0qF�m�ϝ�w��^G�7��=�	W�����ndm�����6X���)v��}Z$~�Vo�{��0�/�U���'��[7�;�D���A�i7d_�.)��[�)Y�	��3�P�E�Uʋ}�h8~�>0��o�c"6�%��)��p��K�/��^���i��b1��W��ڿ�%W'�ñ.��`e�zAFGwDGW� e1�`�I�I	w\��[�9[`O�qä4�vMi�T,j;���@�����X�cb���b��pF�u�ݨ#[�z�VO�CEV�M�����ݛ0��^F�-Pg{�|���(��'O�U����?^�TOoh;~d��kdG�Z��+�W�_obK�ER�������v���=� ݯZ<>*p�5F���D0|��,q�͆Rs�-d��J���p_^�`�O��4N�`�9���w��̡���j���h��vf�"�D�^�p��������L�Ƚ(�����^����m�O�l_b��D;�RH�mX�bt�-�n����ݯCc���~�{��.�@��ݝ[��E��c
��?�br���5:|�7�]"=Up��wϦVL�2�^]�R�I�j���t���'�|+� iI�g0��`�a���Y����)�agC��|�9�P�9����S��-��џ�u�����N�/�������S��􋀑������������U�ҟi�(JLS!����y�73D%��`����S���{�f�5|1��L��?_�F��;qN��͞�"γJ�����mv>!�\C�u\|�f����K��2��D)PM��b�$ĭYukV��2�!<��m�`��jw1��'�;�55b��!���,��;m�	�+����I)�W��m9xVI�T��jlk���AW�ƃ��+b�(�;�1���Y1{ktIdZ]u�E�&i�lLx��m,z�	�\���u�K�
S�J�xd�o8l
�Y		��ߎ��Jt*�S/o�&$��N
Ǚ�G0}/�ӍQ .y�F��a��h���]~�$��(����E����7td���dީ�LU �Q@7��E�����R_�^Zf7�J IB�9^¤�9wJhÈx���x�F��s"�Ч�!�e%1P_�Ɣ�󢡋���Ƥ �03/���})�|�R{�c�^$�D�l�ŏ�t���n�L=��_�ۇ�2�=װ���v�a���W��F�o$��	��E���;�V"k|� r`�F��f�@������1��b� ��vw%������y�'���;��m�ɬ�&��L��<�|n�]r)z�b����G��M9��S���_K���˄���?���j����^7���z�8�G�k��F+ԫS�}�����uc4mt	�u�J>�|�N��)_]w�c)��ttp��A�p�a�d�Q��� u�i�����ݠo���_xl�Aa�R-A��>��~�>>��J;�����L�_�|#�	A}�6����n�6�&�0�T�7�O�	�L��	�7��<`\����mb9��a��	���_��7-U�ׂ:0O�y��[ke1�
�#�(�SA8$
�Rs��03����UGH;]7=ѤYS�����!)�����I͘\g?4E=�ث��XWB}�@)�mn�XNC&��$�<d�&9�L��D[�p㣖Fj}��R�\��@^�}��+"ɽ� �_�]o�%OP4��7�!���uԑq�6��_���7q`cֹ㿱�GVEm��K���󔚒��^3��Ɣ�T�D�(��"ڇ�Ql*�gqOf��=�n�'��3\��Q�ZRTR�`�G����q6�f�0@֑-�ѩ��p}�PF�p. ��p��˂=3�}Z&?�#�s��s,z�2����F��A��r酣��}�b��փy����s���]LdM��X�6���]Ci�iV��o��p�%���'�������p���ʐc���NW�4�Q.�a�h�X��q��+��np�o�b��n�*99�&��]7��p�a��Ý�w��"�'�u���b���]6��"Tm�`���엮i���WU������(��d��������"��,�%Y99UX���*��?����]�^{urx��۲������ʋ�Q2��h%�����3bz��T
�"��˨��&�c��	�lzD\j�!2�h�a�Hϫt�H�%l��n�����_��{�q��=M�m�]-��?�%Xa��ͦ/[��:0��|]C�Hf��lg6+��![;�;=5~Zފ�ո��� "U1�������B�Bo����a��&f��3=r�ǿ�w13�m�9:��s$�J�k���4s�X���~�Ү�'� �X/E$��`���p��d"���*����.��-�����\�Il8�� �^��5��RTڙ�Nq��_�ftQvW;�����Uc�eѨ����'ͰV��-��aڄ��I8C�d}�H��ʂ�����Nv�����s>�:8�����25۪����>�l�9	ܬ�PV-��.�h<�U�XY#j�x����ϕ����5!��Z,Nܵ���hm�a�̈�mᕑӋ���U�(꺦�
	��5�K��0�|
���.�^}�sl�I���dH�՚3���e���}�K�I ("��;Kc�Y�+ـҡV���,?0���[h�mGU��
AWA�����2�s(f�]�J�(�y�.��6��Ly�qSL݄��]�TE�z�u	��ɀ?�"�N�CL'������yJ�2Oo��d����`m�R�WX%�tm��Ʊm�o"jf�zD s���Խ��U�̱=��A���i��&K��� ��D<V~����ޙ�l�����G��>	�0�Y��,��5���tv��;$?��C7Ec���Տ/x�{�P?Te��:	�]��$UL'	|��O����0sڤ����������Kq?|L�ב� i𣧋�I�"1Vc����N�rA\��rU�тȅa]�KKU*�7�C���P�@��2ҋ�L0�kc`�36q*��h`�S7�2E���ۭ����j��4u�|��JS��A���͍��k�6���W�v.�=dǴ�ۛ��&XS�c�-�k$_5?�(PA]�{k��Ng��$Lն��s�>���៬�<��H�@O��"u�!�-�"�u1=c�>�z<�9i��1=]�9��Q��R���m��`:\+Sm@1{c�Ke��������u��� ]���.�&Y�ByWA��_e6����S5�?P@�zҜ���xIʕwq?W_U͙�ͅ��u��d��v.
�����H䏺4'ȼ�� %L�&��	�{�V��C\�~���ĭ!����c��J�2m~-JW��?�� S�q��F�R���U�W���ie�l�4���8��#��n
�f����^۴�H�G-��Ҡ�ݦ;�W�--(@7�su�F�r���ؚ��srՉ�����`��{��=�s�v����ch�b�Y�����T.�䆍��c,�JJ���r-��#-״��֣=�]�/h�TK�o+���Ο�?��N4��{���-ɣ�!�����oJ�j䴰�rr����̄�07�̒$��iu�����b�5���VԆD%�N��ۧġ����i�  QQ"�7�(�7��>4�4W��m�DG8���~����M��	��l��bUސ�b�j�)zjA�1�,x$���G�G��6Lٰ�QtC��ir_%Ð
T5"��ZIe��#�!�"f�g��;��r�zh۳����1=�u.�l�SWANᗘ�_O�����Aleڝ@��J��~���	���T�FfIPE][i�C���WV��ѭb��u���](����8�SL�]��h6��:�|�y˵����)�E��rddS��G8�B2���? �(�Z|��ϳ�'��' /T7�M��w����=����j�^/_q���C<�)�y
����?�%����ۇwJrO�"�u"iy��olG��K����9@��b��bi'�+0i�o�>��0��� �ִ�~i2�b��D�z�����:1r���L9NE��e�4�hCХo$mNT��Pб@7�nbSү�6�a�>v�%f��qf(�)o�S��(S������C�QOHw��GM��S)�2jb4�ЦWGJn���/L���*H�*����J�$��L=.3�du��v2��7�B-;y������H�� W��o�>����8���1#��H�M���K�אYW]�p�=�_['|\�X�@��F	e7ꥥ�0d����RjrV8D�Z�7:6-���_��?T���A��