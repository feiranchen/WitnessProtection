��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f���*�x�����?�o'x$L҉�#�=xWSRϔ.2�ZHr������{}nr񋪹us���:CJ���w&���Z�}�Uə�Q�f�m��:&rrFבȂ�������V`��MU�-���ryyO�]�p�޷`����g8�'V�����/tS);�d�svo!x����u8@6w����!3��$��#��#�S"J�."��3V�I͑S���)�=��?*��wpS�ҘPN��0�K5�%o'1qu���xTad��*��ض��]9{U�3Pp�y�3���|�\&Z����-�\��	�_��M�
ۥ�e�8Ҩ_U��A��[S�e7�͚�3��LQ��iџQGՃ�����)XnI%�]�զs��5׫c�6r�~��4M}ؾg�Df��#2�}	����:���l��Y�A��Bf{(�j|�]�Q/9k�rmb����;��q�dO�J����ԁA���tQOM�a�����5/5/�-љ�&��u���6�sl> Qu'{�T�D�)w|D]X�.�YG�B��I���&}�{��6:XҶ�f�a�]O�n�2�@J:"̪(�4�ҀLOE��\-&�>�n=�{,�R�����j_��v�����E�
MϔO\������̣4?��f"���00#2��'��4V(�۲��A�A���T��Յ۫3K�3����������E�q��i{0�>Y�y��b��&0���/��5o��X��_ ������Ě���čH�M�P.��f����ѱ��ep���̡
-��I76��*���:�^����z5��A�e��*L�9u��Oa�-���,�y�?vXm�.\Y=OץE�i��\�A�r�{�U���ǁ��دZ<�_�$��޻�<[�~�}ŷ��_�x���žP��2ħ��!��ۘ���B��1_j]� v�����(�ؽ6�g�-�{��7�7���}���7X��,���E�*��qa��g��C����:(�-�NS��x����sp��cͿײ��e��JPGת
?!�������
�C�}x�[�`[t����u���82�O;	l �O��`��l���r�4B�s���
����P���7E)�=�Á�U!��$��'q=CS�F�O�sV���u����c{�����+Z@���[D4 �>!�b�#�f�s�t)���/*vG6Y�Pt�E{Ժ�R@���V��߅�B��a8{Q�i���,+��&��ړ�$��՜�F!2����+Gj�3M�!�j�ͦY�-c��<���;��g�:��(�E.)�E����D8�����/=B�v�@��������U\��}tRgh��r7# v{@��BR���<!^g�.�6����8
�.�D9�j$Է�m������*�Y��EZ[�ܸ�u����8�H~�� �����zv��Yg�^1�[iX�T�
޺�b7��������xF*� K?�� �)��(��ECk�<i�B��~ _)~�w���Ȳ|h�'=�d�\E�ƻ� z	���r�Ru�x�6��*���8�������>�����,�H����}ܔ��r��'j 1���A���G�\<�="S`�����u�.>6�VOBRiJ���(p^wr���=+d9��W����@�p-�^BJ����~Vf�G�J�3��	MQ�e�T��t�x��I��/��q��
:�MC�MQ��	��no�k���<��@�J�	� ��mx�,���Kb�$Ԏ����!Ҋrã8�B���d�[�a:��@
�<�;/i;s7hp#UN��RDȾ8��#H����	��G�ʇ,�A'�-�RU0���� |�{AI�� �@՛�kB��l�:z���j%>��f��S9r�b+�P|�����Ԧxl�O�7��Ɠ.��1>���*��'ǝΦ�1[���5�����@ø7��mXM���5a�в�����2;�)5����}m�A�A�["���ux6��
��T��P�}�l{���zv�F`m[��#�4Gp� f�
=��H��l{n$&,;�0���`P�KF����h��'K��vf�%�>�����T�-�������~���0E�%�]7loT���@(��Z5KB%W�@D�{��ۭU�)���..�2�G5?~��2��jxh���?{WlP5z��4�PT|A%�]���J�Zȳ̥��."�LZDj��C-�>�|9��"�ep�w�po߱	TӇ�	��gJnD��7p=�����Nc���Vc����г᳐P�?����ZO�c���҇*9 ��Bpc���/t-O^Bi�gPph�@_��؇�ƭuy��;ȧB:A=��ِ� �C�	vMJx��8�uLm�P?RiR���d�zMQ�?���:d��ceY�#SN��f嘠
���������z�v��Q<�����|[���7ԺN��:5�ǯV�{�|��m[���7�z�4�(� ��e� JX?o��wپ�}Ǿ��䨧��l�l]�
N(@7�L<��I��l�$間4�P�����g��A�B��k1-�M��g�W{?v#3������@����&��b�_gA�l%���lک�?�k|a��kď�$@_#�͝��F����u�q�$��&q[�R��<��?�?%m�J��2��P�}k�e*��vq�����t7��r`��2�/c���*T���	�[���8 �n�S}z�c��h)��@��_�zm}Z��CP�0\�,�{�9���Q�?�y��Oy��P�6<�>�eOu)�f����Q�t�q,�$�n~�s��-7K��'���]rD�<������ީ��)4 K|��?(.~a��P���$�Ka�LE��7Ӽ��%q�뭿��5��dPLt��-����dRn��.|��͒����(��7h�j��闃;n� �O��f�G:���n�����\O݊�	���[]��sż׊��絣蟆��KOy���.y�z��MC���kzwe�A�a�&ƙ��Q�u���\�Wz�P�4����Bh0�~��n���j��}#�fg��#��Űb1�a�I�gb�,/�G��1?������G�f�K��9Z 4��06Xk�!{l
"�5
���r�@TͲ�Z���˓��Y=R��U'O�d��;X-�䴎=���H��:�\"�
�[�I������**��ONuP��}�7�L�F�)��@[�_z��P]�N���窽7�G���(�;2�|7��w�" gE
(||6D��1��i�v�{�b��_�&hA ��8�t=���+oS�Q�I����Τ^��0�٧9&�(Ҵ���9�}������,u�D)Tߌ١�3+��K��O�Y������[ԛ&�<�x�,Gg���Y��\��W�-�0��ڪ�<���˩�z/��B�L���F
}��ev��B$���r��=�s�u"H�-�\��
��9��7d�O���_�Ӣ���t�! �R��#����^�8G4���}��� r[M��~?����Vt�~�('ϔhyt�X��]
�G�x���8��0�!%Ar�� ��`��_p�|��ª����4c�?3|}x5�%��*O��eTdC��5��ڤ�p�Y���
�Cv���p�i���?�r�Xq�h�RC�F_"�Ɯ?E�ߩ��{���^K�k'�xy'�;S���.w{�~b��|�a�[�{�e�%~�L~�JI[˟��֙{�G�e�'k1�('w��*����r2��fp�x5w��.��o�-y �m�����n��)Ò�Z�˸7m���'S���������r�Fk\��������>��F����n$Bs@茓|��%�V����H݌?P��<M�@6�@>}�l\�Q���q��x�xT�r�O��t����>E��P��d;��Ђ��ݖz���e��i�^���Lu�žB�mQ艔������i	eo���Kc)�0Id9�I�
��V��f:m�P��\k�N\��3��bP1�%	q��d�m�%dVq�b�M��|��2�e�[za�l���n�g�@6�i�O��g��.E�jM0 f:���Co{�Ȃ�!4��(}��tA��9Vsp���k�<�Qb�lx��0/��m�pff���4yݧ>�H�AS��g=��l��7�ᚶ�M�F��m�U��25���4+��ݺ�2��}&h��20Tv�Z� L�w���I��v۞+�^�m;��g5BZd���@�v�/>���uxJ&��grdH��O���e����gռ��o$��H�4��NF;�k(�|�Ax��+e���e����on���D�� K��m@���g���Y�zZ�����A_�-$���m{�Y���u7�c+�7$��R���1��ŧ/U�#�[����&B�
6*��x��gv�L8:�.[��P���ͅhH�k��������7p���"�2����������Z�ǌ$��dm�Y���O�b�mY��XT��Ԁ�-�N���/��	��bK�߃%H�Yn[qݜ�9;�RSn_�B%q��%�a���m'"�ꕧ��>T�%�̹�4.Ęԉ�I1b�j 5:p�N���C���kkH*��d���3�j�&�V�����ԑ��B�Z�ƾ��?WX-T�}o�\��]�z ) �SQ��;�*���`�M�u*�yB_RnW8]��O%,@^�%�QK<�[��J{������'�(V6�$���3yn~��mRcG,.+���~��O^�`�OGA�@�B:���;>.`�p���}� �Ǉ���H�+�1��	g�,Z��=1e�\����.c�K0������茌aItE�<-Ğ��bi<d��"���P�R0
7�?&Գ4�.���E<Vp"6���\U�N�:f�s)���t��1��
������ڠy�W$��b�RC�~������߉uy\��I",ar�B$�Ð���fY5Y��l�j���A	Gp_�j}�F��jZ�k <�MAK>͗n�Uf,���Z��3��ټ*�sEY�bP�\zx���y��Q���9�X��$��T7^�~eٵ�9=�%CpѵQ
A;�w�*����96U���؜�\e�����75���Y�P���Bb�K�˱�?ҵ��q�'��f���=8{b�������]���^_Ãʃ�FE��F)�iRO	.��bZ�P�YbEH��<`�����&(�E��������sO�4.��`K�ti��Q��*)���ze�$w�G��h۩d�4���u��-]�OBj��}
>)g,.���I����_g�����[�R39���T����&s���Ӽ�q5=UJ��GWѤlT5�Ӧ�["�4hr1����G*�_�|�e���p�c�"|�N�(�|�
K�3�B��b���W���T/}��F䴨�{��b�����\����������͸�FD��lXh��M�1 '_�.ɘ,��#�����(:��tSN%vMi�{����%�{n�] ��Q>��֘t��]?�T#i��nr�5���:hT�ۑ����H5hV����]RF��1;!���i=>4��g
�`�����7�9*qa���^ץ�T����J��l���zM5yq�}�􁡛]v��u2���_��L���rI�I�����?���~��7Q�HwL�-b*֢p_/�x���N��v�ꗷ��2	a�]�ȟ�EJ�c�G���Y�6Y�8�����D�R���� �4Z�f���gN3\0d�
�@!�5�&(�#�v�9J$��`��:��j�rt�	�_�f�Zu��ud��kV,�� L���I8�>ݸa[[P�i��8C�!����}EٳAt|�Ub�+��q��g�Rl�N�)�@�?SeK�ɡ�T[8?�6Yk�A˄�]�l
s�1ρ!��u+F�Xk���_�C�V`J��F�`�ܘ��*~��M�+v�/G���u/����qh/�C.�c�oʦk��#�u��$��u�i]�K��}~>�Q�E`��������+¢4�>3��zuGuk	��C�{������Ӫ��u��]�ô�8V��Tb�O3��(%�� v���#!�4.ݜ�Èo�e���
����lf�I�w
�5^$Z�7�qן.��H`8I<�D�>{%�d������M����K���О����7�p���U�L��X ȃ�+���iv6�t�R,�Ξ�9���ʴ.��^����x�NC��T�Ϊwvx	1(H���<qYt4���.L�t>��Grf��V���^(��ԃ(8w{��^Z}Rj�ǎ�/J�%E�Qi{�@����O�_���n"J��G���2{���Fb�Iut��p�$w'��ͥȚ2<����}�@��+���2�a�v�4���[�����Z�yN��<�"q['u���ɂ!�����7o�TG�\g��iUe<>:�_C$�Q���G�AD��=ob�}���E���8�a��^�[O�]�>;����x����'���>��ҎXi�wGzO��K��Ղg��&��W��0���)���^N��%��:�SPh@S�����_R�<��C�[`è����[��1��}������YdA}�ȭ`�~�:1<`3��te�A���ək����=>Y�M��KH9L9�*ͣ��Y�@.�����B�7Ij�x�<�Ƅ(;�;����DMo�x��I
� ��Ʊ�%�^�Q����Y&�q%OS�g`��]�˟�P���-\�S�\����O�w���(ѿ~�;����4�:�^�<�O��<Q����M�w�,����ʷ����m���L�3iH�ïs4��M�d]�� $���H��-�����4��aS$���´M��&�b�j��h�l%&"��T��?7�+��*�ӂ���A�6yӷ=<���_rⰬ�d��whƼ~p�@+�)�p��wO/�f=�:=���:����1B���g�����#O
b�����#��z�҄ ����[2�J6༝�q�rRo̐������l7�#"�6�Ku������g�6��Զ�+����%��h���V���`�4���F���ۿ2��L�w�R<�j�H/8b�q��L ��|w	I7�ڔ��g1��<�,�`�FʯݨD�j��B�b�W�p�1��^y�8xȫ��!t���lp�]�����U=o�=��L4}S �n_ rV�"�ԵM8K� ��<�3�I��U�659'��\ՓL����.JAK�]��\h�
R�7^�Db�%�0���� ��i����)5wl��]i��f 2�4�&/z��d�.�%O�&_�&�\��p����ھ��OߘY�����}��e!'�g*sh	R�=^_�,�0U1����)�e@�sy5�QYn��!{�cmB�8X�_ס�Ѕ��t(��}J����5��['����\Z����2�����ٺe�	+�sM@h'��(֌Ax^�C�m{؍v�o�G��<O�[jM��+袪ɠ�A��쥽;��L��[b�� u�v=NG[�ah�A�W�J=�Qthۧz�C��8�O�p��z�l�X�IR�:�Yl:�[e�w�_��!��Re��e3WVK���i\��~� ������l7��I�2~�����2d�P����aAF�!��þ��R����Ӝ �_�5� �N-Z���i�D��,l"��gYB�  ���S'��6���G��!Xy��Jis�gy��y���x��4��w��4n���GF��C��um�t�4�Y�������6�-q��7�fWY�>��nHu�MxIn#���i葚�CP	�C��b(xx�������2�� ��#byQ�'o�s9sAj5��l�3����_M��9{��=~Y���޸�Jv���d@�&=	$z�ׂ�%+����w�U�t;p.�H;#�kCg��� ԗ���g����F�[H���nY)O�ت������S\�AC��z��ccw�"n��; ����ۨSL<�u��,ʷ��q�bI�=�L�l}���RmR�a_�r�){��)��G��$�aV[�B��ld�`�q׉���6�9jEU0��!�k� F+[$3r�c8��X3�{�Qu[v��<���]����p%�Lf�Q?�W@�&��(�ozxdU�c�R�gY�ݱy�\i"e��k��w�g��_�X���do-"k��B����}���f��dA8�^|2p���Ag���:|���('@���#�L)Ӳ�9 *�{5�!3z���7�@r�{���՜N���։��� ��Y��x(oI�ԏ�z<K�.�s�\��$v�.�ţ�9ǔG�`�	v5JI��8n!N���^����Ő,vC��(��b�o��]�,�_XaM}��C�����5#�1�@�d�l��5�ϫ)7��ዝ�X�߮;\O޼�ߍ�[�Y9�=,���(����bMy�1��̓�,��%t~�%y���{HJ�-����+�/;E�{����:�n�:�C��>�q�
W�c�o�c[�P�	��9"??[k�
�