��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1�b��Q8�u��� >�h�t:{�\�DYz��:ϒ�L��uf�P����r�Gq9GJ���F�5�^�'#�t޾��3D��h��L$���vA�O7�~F2�n �D��;F�,XM'�Ct���o-�k���e�� +ڋ/1_9�c}l��K9(^*�����h��6[>��Ψ�2��C�����Ύ��{�qw4�>�'ȹ��ID���K����@}���Zَ�h����QL���c���.�(k�rSXB" k�����[2K$iG�6}�����2�ش���3ޭѾ����d�"&R`}Za�_�W�aNK���n�/~����qٹ���	o�2��z�*���b=p{}���n���n�h�jB��t�x���(d���#��P=�e}T�e��z�y�X� ��z��I��#�X*T&��<s��=Z�	�)m�"6tk�F1>�zFU>�fQ(
s��!0���V���WӟI1���pK�̦�NW��>�q=��
i�3L����h��..���ĩ�����r�!�2%*f�<[�R&�	�Q�pQ�!�=a\<`j���J���
W(��z8����U=M�$����cw�cd*1�T1%��<!IJ����`��ɲ!;���q{�-�!����8毞���߿,%R�����@7.�з&�s=�^��z�f�{���:�L��nH���
E��6۰�F�@ҝ�F��'H���9T�8�C��H�����25.	�AރU�ZKfy�<��xj�����c9)��.�,iX{g�=&�����a�8T�������?3��}o�g� `����{.x4jr�a�.�e�X����P�"� �iRͧ�]�Odʑ9�ɓ[^��ϣDqS5k*��"���e��TxD��f��	���W�V��=�^����.B��MyW�W׉�� f�������� ��T��܍���Lԧ����rFX6���˕l��Cs�\���~V����d��16$���J�[�kx�l���`C�&��9�iK���dt~���=��w�V� �j��u���{;����J�U��˜3|�)�!��:9���a�_)��}�= �8�2��T,ȅƪgo�����[@ͼZW�H�@מC��ԃ�;�Y�}��4B�3υ����#��A������ @�qL�_�-nǤ?Ę�`�+����U�=��<�P��Gd&�p��������iz��TaʣY
�2����Fl9/s\�Єi����<4ή8u�m����J-���-,�ϧ�?
��N��RYĻ�6�3X%P���~�.���V��i�k{�����絹r��Y��Y��df
��8yx��T�9�5an�ΡG3&C�l+�Wt01מ�4�F���#�4-��R�3G�"ƌ(7����f��6�`0 <!����*�\��K�5�T�"�ĕ���ԟa��7�V�(�m_���a��g��J)�x�"O�	�J�NGN����(4q�*Y�;�c���}�"�.g�B�Z\\�&�!����g���
�e;uMmiߴ%��>����<�D16Q���Jx��IyS�yC�P�hB®;�M9��2���!�y�%4e����e���ܚ���@u�r<�W��i O��<�V��u����GA���[7��v�� �S�}{/F-`�3d,�p}���F�X��.Y����ه�|�"�<͙�"Z��ƾ�q�:}y*��C�d~^j�)����1���X\k
w�_5����>��?����ڝ���W��e�9��T!�ϥg��=l��nY[ɇQ��s^��k����d�崨l'4š��(G��#���>eՊ5wv�����D��)qMs*���-�;�^?�ʲ)C�~�>�C�jQ�5)�(b�ĵ�[�!�d��q<�9�Ѱ_��b[�a�4K��gQ��y���
�P�g�� m=Wˮ��Z�e
�J��DpԆ��5�˶�d�O��R㨚<��&��yo|rp`Z��*X`�.���k�DV��7��Z��s�M��C�ZI�Ս6�U��|�ڻ��1���2�Xz��!]������j�'��"������ɓ�;�͕u!T䄅��%�@�3b%u��$�F��4�Ű�I�M�s�:"0V��
�f�*�]��'J�=�9�e���䒉�p�]��$��#�U�
��� �/����
�����(��ɒ|GB��e��f�хZ7LS~���c� ���6ӏU��JZJ�e_���?�������{qcA��%�uyz�8����.���J1���<$���Qe!0��Df��N/�[�ě﷐�>5�E��p�`�W�����rX�<�ǭe�F)NKL��V."��cC-{�<bB*o�d;{^���;�>ݥ2��k��c�B��e�X���4�:����_��ξ��<jI�+a����p�hr��Z����3�_({l�A�����.<5˔xX9e`���X�@�sr�"��0&��[��XWom�|6��_vCe/����	�ٶ6f�֥T��G�˶B���
!�#に����=࣬O)�&��y3�$g�(�\}p�R�L�'֔��W7���($W{�U�pji5*2��@�m]m[�%�,qI�>�)����/�K[S:C�«K�V&���t�m��c�b ̒01çs�+�T�;���$l�n��8��;��&Y,�B��G�	�t,�T�Ț��)M�"Л�fY���s�.e"a�se�w�<�fo�� 3�V�����ӛ:�KX��%�ram�e��cXDR������`q���+����0AhĝKN�Zی����a��	e���G�-ak�R���ͽ�[��$U �f�(u��[����Q��_	+�G��}*�g������m�N�<A6�j^K��'�-{ڹ��D� 8�� K���&9�/D�� hO��Uf�iv?cu)HV9I�&w��ej���-x���Y��#�$�ܾ20���j�h����_8\��y�T�I�(�d�)_��`���CAy���q�$h?�9�#�v>�N=M.���ӝ�#rZ�t��A�{��m�X#pR2粭3!�w�g1���4[�/�l �k�+Ѩi��%v�0�8�b�
P���]�i���Li֐a���y