��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z���"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��`����zF�0�P�:��d4_���S�Ǆ�/cLx�XP}Xw��l�Y^�3x���P�$:%X��|'m��JQd�o@A���a'D{#�3y�aGw ��251T=�]|7K1C��ة�I+R���Ġ��h}�#'�ԔE]��J�S��8&�:F_��5��{�<yP �$a_�o�5+�D�u�>rNZ���6PD����}L���y�ƈ�o��[=3���Z.L]\x>`�H]8 ��0�?6gjT\2̗�����U�A��;���c�@{�뙯�Q`��y�{�u�z	���Gt�	qK�S�.�8��3�͆��O�Žֻ6P��U�2C�
��[g����\7[h3!ʟCG�*Mۼ�Ū�`ka�_j����\�U`���pHp�&�N�;s��=�rľ�oX��J���?��]?i�u�������'q	��F�ص���T�+PD�إ�,|�8_r`�)7���p>��X��t��ߗ8~EZ��b]�Ef�o�3�:t���3��-����DD3&�Vގ)�����Av����w���S���9c6u���G}	l�������l9��l�(�>E�u��h	$R��R�������e��!���¤"$��T�#c@Mj}���$�E`�k¿�+gn7р&�i��)�����w5;�n%,M
�����?�c��K'�s,> `HM���B���	�sG�+����)cǪ��:����d��ѕ��|��/88)�����S��J�K8��ژ�jJj�|W�����L����Qq�H�dT��ɷ�p�'��[��5���&�or�Qb4��%�[qīU&���)�i�������~���n����=Εj�h�l�<>��p���9)U��TjF]x�v�ʂ?�sE�r��
o����V���F�/\Fm����;lF�)��_��(ȁָ��_�^��yL]a�'b1)S�f�b������Z�ss���n���V�s@�&aPT�YmY.�����X��T��I'B�D4�B� �J����*�jA�F�v���҇�00��t�ʞ>�yl��>�
��I �2���7�����?nϱ�����L����)��n���m����|M�r	����7~��������S��7c��]_�OS������@ք�����Q��-���L��u����j�3��3mi2Fq<�g���5C���9<�~,�>$91��kue-����VN*" �󋺌�@6Z���"n��_�2��%F��
�Y8e��h�2���F% ʋ��?��������Q͖��3��$��~(#��	.Ϋ��h�sqR��?̅�����1��>*������+1�|J�5�1�4`��7�:0Y�E����S�-'6�����
�� ~�WR��uç���Ӏ���� ӇS�;�R�kC�,��g�)�T�oN�D*�ɏtc�_��IܨG�������}��M�P�� 37 �|7�L���.r���Np�Χ$��n�SZ�p})�� ���,�L`SDNk��w��)�=���N�������亲�a��H��ZQk\m�k�v���ZA�϶�#��a��)!`�c$�M��n��HZ��i�I�OT�ݗ0B��@!p�W��GJp�h�\5��ؠ���({�`b?���ۋ�~*�w�H�R�`Ńv@+�g�KLn�պ��	d��n�f���q�ϲ'�R aI</�_��l��\�3�3�[��;;v�4��wZW	�:�./RD1�汷?Z�0m|�G�c*~q=��MM׬�����}k���_j�a����w�NsB�K�P'��co6Fc���o��4z���ȟ9g�ks�q�<��@9���^H�FW]k�X �`�������9�v��=r����#IVy����9�a�;/?RT��dC 1�X��|?:���k+��zENo�	������iH��`�|?�3ֺ��2
��G�`[Hj ��%��P�NNgW-�t���]j5c<)K7p��{)!�G�ѡ���q,�n�~�#յ �Կ�S4`9�Y��ITkO-|]q�~���)���8��E07�GrY��#���x��R4Z-Ҙ��K��:&�pe0��u4�k�@������R�~h c���48�i�
�ު0@�TR��i�E��m�C����+��炴(�+�����A9KHL$� od�i#�5ǿ�"����
��;cSU0�_]���)���AWp��k�b|�M��?S�'"`"�F������TNQ��j�J/!�`Xn3��V:�{�q#��j�{J'�2y}-��&�{"�k,A�2x��w�9R�UgA��xW�_�˗�����xxb�|?�N�mƇ���F��-�D���=1���У�'B�9��F�)޾�S���#�>8�X��� \M�S�t3�)��/o��|�{y��)|��'l4^�r� _q��iKY
�g\B��{���F>(-)d�l�8Kv��^�f_�H���qdO+!�M6g����`�t#K�\��Q�8֫�>
�{��RW ԝ͙`I� ��M"�~ߞ��Ο����xv�����0/�9PB9|��aK��|�w�	���gZ�.��;��Ցg�&�L���1�������i�2�F��̓��:���Z�������@���i��5CX/�+io������K�9���f[ѸIн�`J��F(���Mg�ښNDl�tS�uh
C�\��m��q��t�����1�:�g�{ߣ���*�_��QW�⮖l��qp�f�G
l���z���]=Ԕ]����#��L̄#���6
�F|<�т� C��)���}@k��:>n �u_T�{�'q�Ӟ��r�v����GU�!
;	�z��y��`˘�!�/���m3����-���PHj�b%��-TX����]3i��Oy!jͩ/l����o��+�Ʌ��F�	c� ,zl��� ��l���~�p��ڝ�F�� ��#RՌ�Q0��\e��Y�q�&E�	�I�F{{��;�Wq{�M��d1g�*�,����ƃ�:W֬y���.�� 
"���;5��_T�B<lx98�4�K��OUl��ș���6�L�u�HX�Mr�*��zw�6��yl�]�Nv��p�� �3� 	�#�KH#��u2��1b�3r��x���+iQ^U�aO^�N�`6e�VG�����*xr�+�MKȝ(�(�e|5�J�p�p*u.zY��A����o�X,��Q�:���d����a��x|2Ҙ�ҶƑ6~����ė�t����JTdyl�G�[��d:
49�pJ>��4:���y)M8:Z}���!<{n`�<�=�HE�Sy��cmj�_����?9S�
�pV����ށ��tmRpUwt/��_4-G���`�z�B���9��Vo6��C-�G���j��o��`|Y�5���0k*Or�!ٖ�h v��;\@�����V.\���xȅ�*�v���>>"O�����mW6�	7�o&����1T>���|5�V43=mB�㹒�N����`CZ7�_�l��%]X��~y#Ãt���+\3�(��A��Moe?��Љ����Eݒ�l� ��s��n�v�T-�E���Gƈµ�{���2ΰ���\�ʬ�e���fՀ��\c��B�s���qX,
�=�n?�3�Ok���#F$�qk;Gk�Mq�����]����(�hQw#_��ıG{�q��r��$K��ߩ�@����0x2��O�Հ?>&�7�+�
#�	�;�ix�^!i
i��f���/n�>5����;��+���VN�&�nZC�Q}K(G)Ȭ��+� �V�P%g�ӻ`�kA��_�u�f�9�U�o�����)h��a�]�����Lb���C�}�	Yi|�KE�OqJ��iA��}7����]���TY��Azq�����{�n��o�7g&�]a�v��#��,�ݢz�>�z��d�t�8s\�n��$/L:��p�ؓ�v��Z���=2���O%�=�^A�<�V�,`����Qy�.�N%P�J4��N
f����Ģ�`.^*c���I��;�;�Ȟ�L�.�{ᣅ2���ڂ+��.ߘ$r���j�C;FuA��j;�v1Lݠ\��Xp��ຆ����ﱝ�ƹ�ނ��ȱ�>�x�ub�
��	��b������%�9T�%�5�u�I����)��C�M�.�U�`D`C-��ab�@�B�pl`�\XDA({ �z-P������;���;�N�¹��	�5�f½��P�)���ٓ�p�2(�h���b+}��G���h�:�7�Js��拳""�
{���=(V�b��%�o�ӏ^�<�qD�#U�P�]���9�_��㘅�b�eB�^ kH��Vv2��C����AJ՞)��r�G�ߐWu\3V6���߾�I��0�D���%��/�ㆌ�7^Cc)$0?
�RA�obퟂQ��h����$s���.���,��;;&�_~��h5�iVc�om+�?��x��ʀ)c>��I$x�ȩqE�GE�ǠD�*t�,
�pe��%�ݗ�5}���]7�x�z�#��HQ�9�_A��̓�����oҮY1ۡ�J��5�ug�YE:��U�5K�����Ց�&�eZ+�l��a�Z�����Π �S_�}��9�e�v6!t��S��(Y�\�����\�7�2���ƹ(�� W�A�ū��p���:z�G����Ֆ�s�c�j��k���]��s΃�~:��Im���R�;��>�^��w�j+UDwE���9�oa��h�f�s���Z����*/��:�v�B�hv���Դ:��Z�ug�#���A�u%Y)�d>�RE���2�(3�M�J�-��E�`�\�M|����,��L*C�� l���ѣ����E�=�=-}6�iE��c5̹흵�����ą�3�`�Ș�o�,�z�s��u�����۸����`�x��?<X���{���o�ט�i���݂�ML��zK$VC�(�ǳb��J�A�Joy,S:��a��hD�(��s0�&�gm$��F\f��@35�>�݈i30w��v*fx�]���B�ֽ�?�0.�/w*��JF%�2�[c��Rs ���n�IH:"�yc�����:S��Pc���AdEÝP��{R�~"#��:"�U�'d��l���7�����HG��O��zl�/nv��g�u�d;U�	�Dy�$j@�n�����%)�ȟ�*@F/�������U�{�zX`~�F��������ׂo@���"u���{ vm�?�X���/0-g�ֹT�B4�?l�SU�e���o����ד�z߉J�a���Y�&�
��@��FAׂ*��Y��t|O`=K' |#�e�r��n�w���_ɢ�wz�6{Ƞ�ho��$s���h� WD�����a?����I릙~H�g$��yO�1�(�Y�z�K�J�f¨9��W�hؕ'����5|zBd��"��l������I�<,5�A�5�Z}��# ��$�:�8\ʱ�cj�+~^�`d�P��s��툉�Ι����_�ɛ��/ L7�箑�b�~�V]���J`�NO~T੔=U��X�4>�)�8�<���:`-i،~�Z�wy+Hw��a���A3��*d��@,��hI
��3HZ���=E`��v'�nQ�M(
��@�Q���ߍEt���&"�#����� �k_l(���Bb�1�G�����``<��@.ͨ1��2����v7��,���YϺ�B�;j����*�,�� �>��H'xZ�[�����pA��q�'X�傮�ϫ-��U�T�ۘO�#�Ӹ�t~���E����M]${he- �4�ǆ��]k�;ڿڊ�P�?��v�z9}��cj����1g0�r���Y}�-R���P���zb+�6_��񐄈~&����M�}QH��E:�M����Ta��6� H-���Ԙ%S���2�L�<���5��+$�g�[�ǽ�D��V�ȍ��'�n8�՛��+�\���o��t�径��Q,O~���Բ ]�W��Zǿ��|:�u���N��i�מ��\�n�*�;��ú{~uU��v��B��`L���%�f�[�j�'gy*����!v�?����f$���p�j�<�� ���Ձ}9N���a�=�G���iŊ��TBۅɒ�(�R���߷шã�ؑ�(a��{���ok���A�W���=�06m���a %'ېn�c����d���PB�����Z�!��f�縕��PE�� ���1p�jl�H�pKI��=��حp����	�L�\�'��S�i��m������SL�A�R�폁pbLc��5�s?�~�^@Rք�C2�T,�X��������"�J����i�3��`nG���؞i���  �a �C��E����]"��۾e���"�����vK9Ys*,���K�8�{Yj�G� h�n�Fh�>n?����Z�%���x��=n�����A�K
LA?9��v�Aj�٩�7�/�� ���z���;u*�h3/�: ��?Xw��q@Z��:J.�?o�l��1U���"&�[���K�K��D

��v�6�[�/��Jry�■D3�?�0qM��ŷw�Fd�2ypK��� �#|鐅�v�<"g��ҟ�oѾ$�z�X�wel��MFXnf�C�����;� �G��M��"R��P�[б�ڑ[�/Rq4�m>F<u��7J�w��"����������I�6�7+��@P�m-�]P"ksy�s|�#�Nl�\�.eA�|�/��=a��7s�M���=�SI��	`
T1[����Kt��!�eUtܝ�>�>�*Wҁ�1�o�{�? m�d\�ǽ|�z/��S��D�y��ob��9�)Lt�D�o� �7!���z���R^��-_�j[�*��Ƥǫ���U����w���0؍��F���2����&�<������T�u���;Wk��b<mG��� ��\�����i���J)S�%�st��g��e��/笅��{�-�o��Ro�Jܷ'3� ă��F�*̔�7���A)�D,c����]��!�I�|��C�(q=R(HUr�G�p���|E��K#��w{�m)ve`gu]A4I�#xl3��OND�w3���(�Κ�?#�j�����D EU�*G~D*�lk�����x+#B���UM��/��lh�ܶ���D�m���ʳ�)x�}D��ĳ��4�S��Y�4م�;��=7��bi��E|���v*<�p���(L�f�����C�,�j�8��������:�Tᱬ!���a��{7iS䴮"���]o)�LE0�&��f�O�ip��gԌv�Yzi�h2�ymϊ�6jB@�jX��$^�����=�ߤf���۩����ߥ� 5Bm;�]\'�q0��E����YW�\�12���de�����bo,�$���<�}Bխ��fU�f�Ȏ�`�'��̷��b���Zu�O5��n�g|� `н�B^+�2qi-��9%
ov~��j�j��:���N��C1kQȏ�[��B��tB���5þ�d�C`>Ѝ���NI,A#�j3Oy&(��ovIfGi�+e5�PvkKC�p��	�$x���|��֣A\��Tv�4OR%/������򋿯���^�v����ׂ�|'b�� �j���s���Ԃ�7�8�#�.�ˤ�}�Kt���"T��H�)	3Eo QU�}FU@���������ܺ:�M�PR�͠��ACa��a��8YℙT���CP�UHhe I@6ڣ^�/^�㤀�b1���T3�4��������o� U4 ��$�)5Ę����e4�Zﶆ��������D�p�S�O��1��|z�q��۠��#�{ހ�k��F���<L�:Y;��SF�� �l�ώo��5�[�|��7�/��=+w8
քӠZOZ��kn.�iVg�,̉�WFc�&D�����C5%1�� k��.Ǽ`�=����i�V� S�?���5��d�!�_��"��Q	��c%&�mm;�R���n�U��|�!<Y���8e#����h����iy�8�DR���\W<C���/,. ?%O���e��&�d#*C
���o�@���Z��'?�/�]z�J��b��
�ܡ{.�t>ڸi�*��:/-_2)�C+�ˋ��NY2�[��wW0*��Y�$�_�S�G�Pִ a�|?�0Y�l��.�x󛯒	�L��8~��-<Lrق��u7g;P4���G]�|1>RW�%�ל`<,B�w}�*�)d����pRp��N�ʴ�1_o�)��l5����gq$I5Q\��Rf�5&j�i�	���;__H�&ID#ͶC[���3��Ì��u���_��i�ː@��ú6b-�!E����ݬ�w��;+��"����7o+��T�N����o�L>xA���I�[�Ȑ��Lktl��3Q&�b$�~�	�͆ou�<D�@h�0�D����B��Ņy��1��f	�U�̀5$w]����M����4':�䥯P�-��jS�3���ۿR��_�A}�<>��CV�弗�+jl�#Еa˟����2uQ�`�2���?�b�Iq��?�e�D��5�'!L��r�2��Z�Z�p2)��`�e�?����1Tţ�CQ��#��h�)�pƁ���L��'u2Kb��UY���е	�f
@�d�{_��Ԣ�Ǭïr�DUn
���%��~�Q����IKD��읮W5{���R]���恰:J�0�HY�B��d �/��BV \���1�s
������z7��(؀7s���=�)���͘G�Jn��(\��M�ko�6z�@�{��g`Nqf`��|���Q���`L�Y�&�7�T�$�� ��|�,�U 7�I֘I�Y��U��~a��!�c��)g�f&DI	�O�C$�r�xcE#�b`��_��ك�z'd�m�a.5	�/���1ˇP��D�R�nj��]vD0����,�B�}S"Cc;Oh�%�gH�J�M��烓Bm� 3{�?���:��4V����@VA�݆RyT���1vϽ]W��uW���"`EX�=�G�O-6��z�N�em�C:tW�}i;�ی9�YP���t�@�pj�$)�t�/~�7�	�ͶK	�Xhj��̈-���m�|݋��d*��x�ڮ���4��>�"P�J��{7�c�����q���:��\�]w~�t����Q��xJq�7��'��*�R_�s��xkc�����`��� ��{�H�q56�$}�e��j=�P��Kڅ4�C��Oa��;13��/�� ҵ�ի�c����r�F��p��+�^�w�,2�9���P���
!��p.�U�����{m@��Q�H����'@�Қ��6����}��7{��K�\P�����4���̯�MR�-�/�k��n��c��!������E�ݬ����V��ԣ[{��ep���$�:��p���<���"	��ꚫt�^����[�!}�����rq˺�p��/��?�����c��+E�����N���y��� �. �������Of��m��q��?��8)��	jdA�U����D:�L�l��XT�,8K�=��R�G��M��r�.j*�V�A�ߥY=U-=���M�ǯ_�8��7��Č�+U�.r�M�3�m���F��ք���uX���)�c�Ǿ�s�������7���BԝY����,�#}0����h����`_1O(8a,�KG���ly�d�`+�@��ouU�9�i4�Oo�\gK���`*��K��0�R2i�c|$�$cL��k��G;'���b����q#C�v������x�-K}d�m�|�樢�E�����W������n#�'v�L�t�e���'�����{i�S����V��r�f|�Ԑz�8o��zD��TK��&߰FH�"?�\�d�����YhJ~�H<�DTy�%ti�po�+�=^d�C;�`�lq[�'�m��x�$y��H�� ~I��(-,s�r7�?1.p�)��0$�Ͽ��u9����3���
�_��%�{�)p���%�o���fL4�S��u�����@� j�v�H�
���8�</<���!�����t�����7J��{���Q�4vp0s{��}(Xl݅h �
�4a1q�=u{�ʸf��"����X�
gP���,[}(�
-�\X��,j�z�i��n��T^T:���0�k.D��"��V�fűh-�>�#d�>MŝⅇQ���o�9`f����
&CÂ*�:���Q��\$�� 7��[?o� ����M}w�f\7y��Y�פ�@ sN��"��3�(PT��2�L�.�}1��wf�d״�L�I&�(?���^�Ѕ~��	}~�ܾ�s��r�J"�ح���R��	�����ܞ9 4Ƕ�V�)7�:	!J��_E�N�T�Ȭ��{��1dm��|�6K�>c���*O� ���9"�`Ϫ���aR��Ճ��?1�B{�Ă�5EbxT��5m�S�9�������_͎���f�>v:�I�1�;������&V�Q>%���@T���`�<1oK>u���i�d�u��̼4���2=>Gd*�`}AZe@�l�yz,nPJ�;`�0(F�A�\���]کg��S���iN�R�)駴P1��5�w>V�D핝�e�u�h��ס[%���{���B��˼��f�R�J�w	�E�x�y�ǋ�ĝ���QF�7���y	�4p�/A�F��7�B��á��M���$���ڱ�*@�H��WvЅ���)F����M�\�xSؘ��*���L�Yp�)�c�5�+�2��3����Э�^��GD��I�>�v�[��D�nN�Ӭ{.�hY�R3���� ��@�d��x͝/��� �����d�p��7�VS���1B6l��DS���/���P_f��sC$�]�X��Ӄ����x���F�81�4r!�߂w>�$��|�����j@���Qց��X� ���E,�Ei��8$8\m��
��%֟�7��+0��G���Uyu��I��2�~�\�	����B8k��9�Ӡ=��bw߰ו~��;/ǃ���t��*�(��Ԧ�A���Jj31C������� o�q�X3D�D�R��^���e\�0�j˄�1Gԃ�h�&�H�:q��itUڜ�'�
嫪��UC�&('�dJӲX�ޒ�P!�J\�4F�|Xdb���+��2C��~��,<��`Y�RZk�٢���ss�&B�0,�"�E��u�QU2L�b_E��<��ن�G�Y^�\ٖkR Yq)�%G��֌����7�g3��I��xq9v��e����}�E���qL��J��G;z���m�t�Ŵ!����^�Hm�7�J��S�����ۗe������^_�GE�
TX�o� ��&��ˮqG'S�PR6'q��5��c;��C��g`x�e�N[��b�'�q���C�3t_�]eb�G�l���̕���Yk����iE����:T����_���6�����3[G���R:D��݄��cAB�%^�����/�d����n����l����b@�ݻ�4s�������I5%����:Q30�@��T�E ����3�$��<����\Q��o��;�I��Y2���8U6���X�J���b �VjO��ʤw��Ǯd�����:�T��!��*�W=�i:ސ{�r���4(�"	���
w���ֆ-_�P�e�@�n�~ͧ�Y���z�*��K*���)����x�Z�0���vs���� �=��=p#����Lӈ{C�&B�*c�SKx֒?����	I���T*�~2����x�v[)6m9��;IS��|�R�����W�rj�uv{�3��=V�	TG)c��-O�̬�S'v��K���6-����§�'�/Z+cת�Z��K�e�Dxw��䄅�;a.���LjM.C�ꍦ]r�:F��{�N��o�N�-�y)��6}�yX@:PԬ�r\{29��kD�/h#��@��or��&@�󱙕�;��Cv�L�ju��e"ɥ�4nw0>
��1�h�{Z<o����P���.�%� #2׷�ò��Vm���J�%�.		6��8'C������[�MD�K�
4�D	�aU�h4�x��Gغ���b��ω�S�r�
m��[��G�"Fu�Yu���ˎ����XbC�[��cF/)>��`�%��BOy`�6ʮC�ܝR��[7W�Ë"�"�+��U�p?�`C~t)49�e��HRp�偀ܞ����4���y6�cn�RZ�A��j�ifD�~��׮@��	;��A��a��i��?M����jm\���$�� *e ��E���̞k4̱���&_�u�x.����aV50��@�`#Ӂ�SS��%c���HQ���]�JtAzYZi�C_�����雓9Ag/]���"vPR=jvÂ�v��-�|`v.��T�"��_ uU�^>��)�v���5C��1 I���fb���K�=]��҈M�u���|� ��W�+=��ao9N����w�=r�m��@��R)�B��������X�b���E���O�@=��pq�`�z7����R�x�"L�U��p�v�
� O �Z���AU�`�t�Q����K�齷`���Q�ր��g�x>�2z��e����s,�p��݀'�9M�Ju}x����UGp)���E=�;�F��l~>�v��l�Id�;��|��i�>)��	˵��Y�/4�8R���u���<FXTpq�ր��w��|����=UT2D�����D`��So4r-��G������t�� ��by�h�[�0]���Ó��bJ�?b:{�	��Op��geh������w�����xŜ�L�
>���pJ�C�e���!I��V:W�A�U������x벖҅�C�/�K�=!�1vp݉��wNl�mh�]F���tAr�=Q�!������u/_3�����)�/���`�/-Lѣ�G�u2��Ķ.��\ԥn�@�ݾN0s+0��ҁr˰�$Q!�y)�*ӕ�I䰄��*`���}7w�/CJw^�h���Πu�bV�`��-m���d�X�^���28���%A=���7 ��l�	�?l�^���I|�� �& �tF������U<k�}�Ke�=gG0�\;�+P �)�X��1��O&]�1DD8���Ur��*N�܇,��w0%�j�W"Y��8V|G��"��ZH�v�)��,�Dl�`$ON�&�]I���+u�(ZP��9`�!˜fճ�	��)�9	t�'H�Ow㯣0�7�ZhW�&y]��9��;ȭ����7V��`��1TB�� RI���z;I6od�3&^de�K�ǣ��+cq)���C�nX�X��g�8��s%�M�9�h��q�[8ִ��:�6G'Z�!������-)��Z�U�tw-Wf��q�Vz-�v4ت��*�����(#(�5���������f,pw���$٧��iBv�>�J�r��'������ܖ�+��ۧ���a.�M�zk>\a�GM��	���)F*<��6n�����Q�NI�O��(.!~�	��$B>�U����}�F���0�r�M\�Y�K3�4Հr�0=�|_~c�!p؄B �_�;�= Q*�?��!��8���z���}a��d�ށ`�9���a�쎚g	r�n�B!���B�j�m�A����)=�2���[���%n|o`r��E3�����0�LJB\W��8d�ƥ�r�i������Z��;��XI�����ȶB���tw��e�0,>�f&��q������I��_d�բ�ΦrA�V�R*F�&!d�#۞Z �G��G��s�\Fe*�[��.�j�"T�N���4j3	Ғ+E�zÑ��J1h7PAp����4�P+fO���"�{����eM֗�{�ǵ0	�<?G?a7t��,�;xF:���s�~�S�J�R��B ���*(9<8�M{ry
�7�i�薌�}�,�Iisoسsl�X!�>��9Px	�ڈ�Z��J�iֵ�(� ��\`�z�w�!bP&`�b��k�k�j�� �8Z�|�$XS�M��ޠ���$���	�)�0�t^�zM. ^�vϲ�+˾a�m���esQ���i0<# u�x!~#�u��,Ls�{?K�{j�a��j���$���E.����J����o�G��T�m�ʐ�����l�!8���J,�v@e���Nu2\�S��nOR`��0ԭ���5Q�c����O���� �4W�"��6��AZ�uƎ�,�Ϫ�'�ˬ<1@�-�s�2���t�SP���c	�m�o�Eڠ���l�5�2�Skd|�b4*��Jn/�E�W��Oi��|�5��HD�v�R]�x�Zy3-�C���7
 �݈1��aI�&��s�t�B�z̕�M}_>/�:E_$+'
'�Ů�c�\���=��ȷu����#���]tIgA6�@B��#cЛ���Gl(֕��$%�(ehi�I�=;;J��r�	��0�z��9�)s�]H�q��'{e�ޱc�->U=�
S\��V��|c:�n�n&�A��?�2+�ҾPk�U�h�w�v�p}rOk�����J��]!���+Q���p���H���e�P� �-^K?_H��	m�
��t��u����QX�RIPjvV����f#���>�$�֎���h�
l�?���MtW�b&��QM욖����p�o+��;_��hh�F�ȹu���h�7`�6
��7�ߡ:�R��o���b���V�Sh^W̭�t���x���|���?�Y|�U�52�s��v�?� � ��i�l�3O&�i�6W�U���:�
����(��Bь��46�E�)ѤWBK��y�a���7f%"*m`f;���4rV:od��C����%L��@?=�`.�ό6��L��T�����e���fbm���.��L�������N܀*�pC�R�r`ì��ġ��h5���S��0P�>�@��n>��-|���r+�r�|�۷�0��nLD3��f�V��Մ���#A���@�ÿd�%}��XSp�[l�X��\���Y\�ܭV{����
Ծ0lfp���>n�//���|��~�Ƶ��ن���Z�RR5�I��H���㣐T �ф~$��C�}p	<A|�U���.c��q�枮��u���eɕ��[L�%~�~��>5�6_Wws�&R��z#��cLH���2Ķ�aIy���Aª.�n;ʭ~����hc���iK����Y2.��w�);s���#�p��l�C�Ba�O��M�0aeh�hꝒ��5[�qU��u���F�+�fwb�k���W�E�Fb�A��9��(��J��B�ERh �r�& �"a�k,В/畢�fo��&�2"�Ԙ���z��j}J�9q�&`��E�{Ր�o1Q+/����FB3�u��U�-���[���������ݫ.f0�ї��!s�нR�0�\���&�N>S�����TL��8�*Zm^��>��Z�Yl/���������]�7u
r�c�t��Cs,�����Ԩ�Ş�6���s�0�-��ˍ��4٪K��
A*�>_�2��_A���<�@"b�L���|l���#ʎ�B�c��=����=cML�7d~)�Ռt3�?�ߙ�ϷW��DͮTW��޳t�+�-x��C��d�Tm�D6��5_E.}V�<��v\C�n��fj��2?�1�� �V������λȳ&7(8aRCtZ��X�Y!���G������~*�,!q���X�o2�U6*�A�G�M���j�[�Dbv�&{�uTt*
��hȏS���À]|^�L�G)�<��)���d�RnsΔ?MG�B g/�}��v����<�sc6a-Ȅ�m���71��fխ�Z�X=
>��3����{)���r���M6�C<���)�@���[	��C��X�y�Noa���7�Lf�Z>.�ޖ������Ň�GNNb����V�^?v���b'/���)�?�Ws\����e*S��V���an-2��Ȭ�#��`Ŵ��*/kXF��b�le@�C:��)�)v�F���'/q;4!�s����0
Dd�'Ynsno�``�>�;H�$�A���O���fuLc"(жҷ�J�h��qn+#�z�9|L~������D�'k���@w�p��o16Z/ss��F�#(�]9���T ��6��I���=i��#9ڻ�∘#[DA��� ��'�<�
w�Ҙ�[��PV)͑BX�6#����n�[ʳ���Ll�>e���A���[n0�Ƚ�	E�b�����|��?��>c�$E�$I`�9ciq�5Y@uB�����ܮ�
�-h��ox�mZVM���H+9�YB���5�U�}ͷ�턯�ɢap�g���>�ouT��M�;�9bߑ?lA�(�G6y�,���YN`��*AEr
�l{�[�cl�5���(��X!�Rh����t�=}��CKZ�:c��=|E���O��d�33�kEt���{���i{��b�l�C����fG^b�[�I/��v��Lf0|�<�0�yS��b\�g'/�gS�W�L��G�st�[q5�rR�6�"A�{K_iծ~�ҡ�m3�f՗�_��v8D*�1o��Gj��8HK�[�����=��	qU#h�Q���O�Xz^�`�.J�i��qCx'τ���v���n\p��gWХ���!}V�:��R(%�j�����������N����s�0d��v�mkj��/<W2��NU3d(AЧS�E"P�q2�=p�{6�� ��x�bg����|}+��p�iQq��f&
M���	k�X�9��r� "n<Lv��&m�	:��'G�f&]���D���e��-�O볊yk�q��2'�o�V��G`��{�"��g��n'����b6QC��/f��iN��5��3\5yUz�(:�5ɻ"���'�),��{y\{�F$�����E�-X �)�9���O�%nЋ�a��T�����ҋ�? �q&��+\-�|�+�����8��*�C�=]�u������$��=�#�\��C'TK�aq��9w�=�oC�)�l�kt��q�/���]JH��_�� �&&�t���0�=���D�&.�_7}�!���T��%")��O�PH��Fñs�DuO�Ib_;r�F3M��מ��%�%��LEG����9��!�I����Z��-�~K'_�xҰ��.3<Y�r��q��j��3�ֈ0AD�d����`�˽'�dUZ��ݮ:
E�I�V �+�*%(_+n2�9N�j�Za�֠��|��'c�@)ht��z�A�ܙ��9��,\'kI���m�����ʶ�A�=�!�
l �Q�� QMG��t5n�èw�x��r��KKb�K� <����;�P�`���9Î��z
�b����S[C��Q��z!���-NȔ�>|��,9S�Й
����αL���$�.�����-�>sK�)�.�ud��"�5�o���B�g4�{[�߬}��G�1�/���GW��� A��R��{�55��bn�</�<�:�\��q �FC�p��F1aQ������pn�ı�%�ֱǓ�3�.;
�������ڷ��o^�����s����^�nŊ6�ҙȫ����S`���b4X�� ��l^����O���}���+v�㩚��F�6��Ƣ9��t�/����@��I�%���}u�fr�Y/�O/��-�2�7�T��L<��]%�vM����K8�R��'c�����<��|��=̉+Y�j�QEQ�H�t.%LcD���`�����~����P8����ƾ�uх�o�����⬄���J�#߿[bP�G�}sz����|<l@��t\��|W�GCer9d��~������:��3�s�:���	��dN!��5TZCCՋ>�W���P�1��-#x�,q�/��Z=W"��RDL�� ew����/�@�/�� PNX����������@�-o5�*k�1�bE]��Vo�I�h�/��!�>�5�x��8b�о�J��q,����?��3�����krE���ƈ�:K�S!�Z[@��u7x�E��8b��h��#�4�������5��I�iOԮ��,�Γ��	���T�vU<�p��iYZ�>�9-�2LS,��#vq'=ca]T� rљ�B$��:���;�6�  _Y��tm�V�>D ����{�X�娇��t�S��61z��9�(+�n�fF�(��.���"8�ԓ�jԙ���n�<�Qf�P�Vw�%?ة����:̂�T���Q����(a<+�}����ɕc��L� �oU�!�l�40m�0qJ�T�WC&^Ʈ����cT��W��[q��O}Wd��}�@��^V��E�ûv���g��2`C�eT�"Uo���Hi8qx99�3�L��͔-{�b�\��cǱU'��^��k2 ��'z}����F
�1?u�pA{��f5<���]�1�ѿc��B߁(�Զ��n�R<lƱ` �1��;�S��g>"i��, � �V #�ⳑ�����J+V%�_��c����q�8�����Mi��a�l����ҨW46��j�2Y�
oo�����1��3���������J꧔�M�����eԬ�n#�pP.��M5{�Z&��\4άo9�{�z+�J�IA�+�o{����sR�6�����."�-��[�j��˧2x��;[V��M�K>�5� �5����-?�
cڏ4J�H���@Tne�f���d��tm��EI3�c��ٙ�	����^-��Kv�4�=����IH��]"�����m�~I��إ{U���>>�� ���U��u�?eSg`|0A�R'�Gd�>�9eg��cH�q��{ h2�}����3��Vrev�D��4FA���F�%���v���N�h"�KE^:�Y��x%���p���op��KPv$���]ƣ�u@�-�Ԑ���̻�qm���� BN�:�vguǐ�m�l�'����zn�3y� �F��+�4,�
Ea믝N���mG�����YJ˖��s�#�g�w˙_�w'?�'i�$T�0�Ц2Ć@��a����d����Y�}S7~5-:�2ܛ]��~��%�R����;�/5�a�-Q�V ����S�x�7V͍��7[�A�cH~_A�A��������������Do�L;�%p��qA"qN��?w{<�8�ڞ@?�(�0;� ����[�3sa>?�3�®�Ϟ@��L�\��V��l�%J�������[G0��7A�[}J�9;�\ {9^H؋��D���:�n��`�=���S�a�F���A��+@4"J �v�9ܱq�'���{;�Ð�䷃[�%]h\�!�1�N���I/�rq��S_����J)�S9%�m׸��o,*�#���\�(-Þ��.�p!�yo4I�+{@�nĊ�J�ҏM���	������DJE/�n#�~�E$u9f5O��(@���C���~iY����ׂG�J��b����j*W��"v��-.df��wH�[�W�+B��Ĺ��tu20������9�/�in�����V&��6�i�Q�d �#T�ͳ����`�����h�UXlE�J�r5\���)}ۍ��Ri�:�F�$�⤙��w��a'�ϲm��W��1qP��	5�F�'V�s�z"k�T�Q*��<�GS���?�}�BB��6;����?;B������-�=�wa���#�7x	A�=AK!����Z��-4�l�u��c
��)B�c.�Ūԁ1��r��#��U,Xbk\����A'��7���Y���~g�#m��&}$Uٝ�̩5�΀*�y+�j�s�*�΂��pf���:��*G�8aߩ��P"V�N�� ��U�\���\�H���qZJ定f���rEh�r_c���Fjhb6x��Rq�^�=hV�����W����t�g���q�mzW�F��Qu�Gx 򏣸�N$rj��B<�x��hZReP��Vv�@-�}h�6��q�6���4py����#/ s���;�I!���t��s���2�&Ҝ����Ľ ������SHw�'a �AN�wC{T�l�C��r������z�}{����������y{I��ݕj&0�e�0,�����]]��?"s4AW[c�<���p\�HL\ތ^$��&�u�:��٠���h:�?-�c~D��pT�.츗�-Y��+���<g��Sɉ'��/�?��2��u����l��Vӳ�si{�u,d���.�g��)pW�� g6G8���t��N3����n��2�{Bc~R�0?x�q&�S���k�ѱL���,+�Y����}��fN�����6�U�9����cpá�ux�]�a� P�j?j$��OG���$�#�=�����`"�n�\}|�D>��^sG������(�S�+;'N^*�;I)l���uX4��rCF�Ey$I�� ���M4<���Ao�橙"��%����J�6#s��n��w~�1�_�m8�W���B�R$�+�E-_�(,ȁ¶�z?��+,�����`���[эp�]u�F��6?w�U��ͽ�`���ۏ�H��~�f7��x/#!-r�H��Gzw�Uc�'=�s17��A�uu������}q�06�+G9D-�jfi�IKg^�0�ע7�@e4m�YB�x��W�D!F��k&��$T&���=N �w;�_�?��g�������R�>{��ٸ�k�����,3h�A�S����v��#�iB���=��v���F#Oy�JWIFE��F�~��AnWzh9����.h���o��Sb���Rp`��tz��J��sP�tS�$��4݀�e���4F��"���". ���b���Y�����'� ��q@
j����e2|.6� �"x�A���Ș���_|�#H4�=0�#6�#|x�aC���U�۞��]o�s=�(������geYI����-�I!R
����h���B]j�x}Q�vb�y9��I�����;�A33�f�����߶�C�ܡ���i���,��0d��N�7�[�|���q�vd.�9��c6�����p�P���Yl9�a$�9�"+K��ԖI��`�=�����Up�a���@���ճ:oNԅ�e���������=�m��eT�q����,k|��`�yN�����WY��mU߫E�,�N5y�� ��EE�����b�~� �@�^�5�D[őn�N�c�	Ϊ@=䝣#�v-�L�'�H��(i�ͧ�yU�9 .�#�d��(�X���1�u˅����͇��|vʘ$��K!�}y��7��7Ě[)�G���S7�S���O9�n��۪�����~�Ņ+,UŠ��v~���D�%���u~L���$�J�Y�2��DA�(��&�]9�tu�)S*l�H�G�b��9�Z~X�=K5��{�ym2�/�C/��hXC�����  ���7bT�9zU���[�ȱOu'��ήm�l���!�?UnC�P:5-pT�"��u��?�:8qya�{dy`�ʤ�	��9Y��L��6�����͠Q�y�#��L�Z�Ô!f��0���by��� ,�(צ�S4��>Ӊ�����f�9�#<c��LD5�7
��3MK���h�8�	q,(i^g-:dZ�h5ψ[-��0Cn��<�З��u5���wW�S�l9B��0�]$S?��g�n(�L��ͩPk�vmV���}zE���ܲ*Pc�C�|�2d{T���7?ޢk����c`������(�h�z�r��h� ��>)H�A�S �EEK���с�M[̱ ��N�-xaJLM|�����ǹ#߮E�0�F��]��ϢI��g�����Ə��ynT����P��4��>��7�������|?\���`����WQYL) #]��(ucC���<��M��,����Dwd��F�X0&6�Qb��hT�!o��}�����$��ٯ��_��Z�[�E�I�|v�����¿Xas����{q|��O����g�v�g9����&a�^�F��vUlzkmtz�R5-�Iq�a��:�1%�+<{u�(�ci�F���+(q���K1~g�`���}����5��"3�/�9�a��V��:A��'׬��#�q~���)���;����Wy��e6Epa���+Vw�DK�~;�I�BI�����ǒQ%��Y��4a�k�nu-F��YЈ�Ϗ��A�+'Ñ������M`.,n�7�|�~��73�D$���e�4����|�_Cx+��u�����/QJ�����y���Q��~fxՋ�ȁ�D�`�t/j!2���n�2�Q`n"Lc�U�Y̨x��N�j��'a?�~�X��.����")�;_�E���-C=���@.��/�����$���n�7�H�mF��D�&�+��$C��L���0AYw��*��S���m{��W<Q��3�{8pa�O+O��4*��K+��juׄ���K�2L1Tm�j"A�]5Pu|�|��)� �&�>k'@�����5+�0 jظ��TIr,��Z��YY�afH�fp_eY(����.�G��o�����\ �eJ�j�2A^�l\���u�`ML� Mμ����4��J|<�)y��C�(���qT�Ζ�PRSG���飏�<҉�l�wX[�ܖf"C��oe�L)����!+D��7���2���R-�'J��Kb�����f��<��o���_�h�`�Q*s�x����f�Yʉ��?�%tΧ$w�q3��B<�Rj4ޓ�g��Qk��#ĺ�	FZpN��'t��*3�n}IX&�"�,l��HT7�[�o��gh���>���p�����)��(�{1�.7�
ȡO�3˵�?��x��f�Ǩf/�3N`H� �$ǣ�	u�]�V0�x�?�>ˠfǩx(4t?m$��&7do��OAW���:���X�y���޼�q�a�RxM��K{���C�K��y|��'X�I_�LuVpp�r4�����6K�$!�N@�NjU��S���Հ0���W.�%ME��o>)���R�<3��=I(��̠Y-�y�x,k��L�S-�:�#>��Ʊ� �ak���p�y�[��(������S7�ݨ����q��������LU�b�Ev%S�T�MoN.o�]*��
z�� ވ#�	j�s��!�S���4����"�ō,[e��I�{��"7�K��N�ϻ�����	.%-�,~�v�
,��=��du0�b~�/N*�.��B�8���@�L�-XC�p4�D��*H���J1�F�m�|u�.�yO1L�葲D��Ei�`.�~f�`����Gs�ɉ�������r�)d@@5����%�H � ����_�%
�8Tp�3��XޢƠ�8�}���������n��^�{eGsc�_#�<Ɔ�(�9iS{�����`�jm���#�����3����iQ��<�U������A���1-��51�	��}!�E�6xE}iX�l^[����b���}5`%��M�����*贤�>=DY�Q�}"�r��=�� ��YY��Z����z�>�
d�� �T/�g���>�8	�C���ۛ�b}�wй*�������H�r��g�{��͔e��X���\R`��0��5p./EG!�>�j�%?j�S6�bC��t�&몠M��\{3��'	z*󤴶��5��m"8{0��(%*�&]�,���&J��!{X�w#S\1��
;��v����+O�h���y�7�������A_��O�����d��h�}pu��G�	��g^x��m�I�Ywa���Q�LrF4U �~Fx¤���\�1���xxu�7�E�t@]{����e�kIn�Si�V:(i�C>҅�U�\8�����;�;*�<M��<t������~��]g�&`��f�O��GqR�CIS\3*�qi�Qc�-a!���E��t�#�.���&����'��&:��? jj��н�x���+W4XX�l�.[&T���NM� �cD�g��W!�݌��x��ܮi-��5� T�b5_$
�'��Z��e�B6�<�̐�f�ޟ�B��N3���.h��#��{���e�󬀍���S�1�7�B�V�03��G�?�����Hi�T�d���S=$��� �e1Hᅉ��,8�KT�`�g�%�Ė��B��'b�|��N�{�P��ɡRR~����7g�Z��'�Ʌ~�W�������e�;=��r�zz�T��I�����?���j5�YKZI����;�K�6��4���2-�N���	�Aխ���a�i-��@�2��vn� �#)S��h�㤘6hUu8˄�q��R쵱'��Q}�Vvi�;X��P�6K��Ƅ������O�傣M��^�Ī��!�J�G���-[NV�븝��'+w� �Ŝ���k�����v�ITd���V��R�] �f8�"���lE�{$�?�%[��Λ�_�2�����mc�t����W��Y�+���P庻X����k��1��@@>�8�����)V��`q<RC6�TQt�Oا�HН^bv��,i'�S�(xw�K9�m��<�=<��y���Z��'%�1�����~��`�(��~���7��f��!uGyϙ�:sF����1rO�88��:��F�|��_�l��M%p�g�F"��$�"{&G��
La�� ��n�N�2�d���xD��"�x�ڕ����1�����f 'H�^3�'E�|V����f�ط�i�� lqQ�����T���1��C$ �Y�-,ě���s��=eΥ����Wf���=k���Ii�:����ow�M.X���� �NF�HЛ�I��4(��/�w�j�D�O$��{�"G�وE���-gL��s���E'�CĹ�
��#���.��<�QC���a6�<g)�g��5ݩ69H�����"9ߦ�$/����Kb���֞�ϯG��Jh
}�l%��Q�閸�q��dmt��<8&�|�0��ɍ�f�v��e!��j3eGߴPm��3�B ʉ4��_���$����I���ve�&܏E�V;��mymc�0� Ju�&kҬㅰ�&Y��r)�2K��U*ϗ��9�)/�>�<񛮲�sĥӀ���Ҫޡ�E��/�Q�8�N��W����]���4��Bq�G.���4r����C�t�k�\�����BKBo9�~T0$(P���'�����:������Lj�b���g�V�9�c��W���[dj��TP����>��_:�r*kE�Au��k�5 �R���
2YW��}֟�`H�w(~�.��Q�T�b�r�d%�:\���>`��G��[��T(�~��hJ~��H5�R�!�vQ6I��e�*�e�UQ�b~\�_�hZ1�1Ry��u7v��u�Cξ\:��8�Z8��$ aJ�c��70�_O�Xu������D�ÊX��:*��G�짯��D�z��T��u�^&�����A���z��㒯Z��C����U�?�t����{��8�!˶A۱ʽy�RWm��y"�����7G+��jg('��H�ڶ��+��f]�j?�/�X��21��`?O�ثV�� ��%_�ʌ�궝��P��jkǇUwv[2�.�@�C�Щq��cq6�����L_�]mS�hєJ�#{Oy�9tl|c$�`Ǻ�ߺT�M�1�U �
!S�`{���t���RN�����}Aȫ���q�b����&�����ER�PA�?�?'�.�Ѩ�!I���#JM�ڶ��'��0K��ʎu1M4FG#{�7Ԥ��9����}<mx�^�)3�#��W9���c1��Kx��a�\]d����A��^t;��Ζ�a�j���~Jvҽ�� c��#/f���
U����N,%�;�?52��5�(1���fTD��Mz�v�,�~����r}+{{��$4�7�:�|�ݎfl�0�1�4�Y��ݨA\mY�tIq*����1�|[�hk:���8�w�k0*5Ұ�.A�#��,+��<>�P�g�o�=���^���B��n�cF)ם���#��K��>�o]��b0j�c��۵�6��wʓJi��߱}
J.y�ǎ�A%��}���S��Or�~�)�s�U�2Ǉ��V���-z�1���N�M�w{�[9��h���ދ�z�Z�PW�X�ߗ�������[�S	�����(H��:�3$M�:�n����y~��d�9����C�B1GL�-a���q(�!�h`�t�Y�1��vǧn��n��F����N)>X&����&�֐�����ҝ���Q���~� S�x�Qޣe�]��;�y==����0�w���f��tYȃ�f�N�����0��aD2�O�Q��+p�a��p����J��Ѱ5���9��Ny�+�6��~���o���_�� ���8]��:�4o�E��e�M�����ivIS|�ۉh�T]B���C��(�A˶�U2L�mT����O]Ob>r��,1�s�B$����1B�?�`�~�������.���^�"�LR�Hܷ;d
�T�F��y�UG��IP�.���{P���%��P�e'-�4�v���̍�p�J����#֎r&������iʰ�I c�8cIPQ%���
$�� W����ȸ��=w��7Ժ�X���URF#�6 X[I�#���!~2B��" TIK��5&�����,����c�;�!�a�!��)_�R�ܲ��Z��W�Ǝ�U����eb�\�Ӥ�L�Nݸ���&��_/d`a�R�u=�W�����ܧi�.o��c8a(������I���H � J���2�]�Z���y��h3�ǃ`l�����q��zsgA��K��bV��]�� ��z���W3>t͖5�O�4����[uFF�aJ�8� ��3�żYU���h�uӫ�V�Y�>��3}���j)�K��쪠ˉi��Ѹ��m�ia�O\��p��ܓq7�)r>3�-�ʹl��H�O�)�F�9�v7�X� ��S�L��σ�Uamʨ�,�feJP��8~�ה��`��?e���X,S۷[(N���!WvۊF����F�z*��	_���� eu>ũ����m|����s�E�S6o >�*j]m�$tai�2��"�D0�E/���ks���y�'m��/�?��v+��Xp�n*���K$�[��xi�6w���A%��MAL����)�h2�ߛ@k����g����6 �wr��CĚ�l�V����\7JT�_�+���Įs��[~���	խ�T��%���g�Л�G7��r+�7[mqelddg�pO�h 	�dK�<�"�� J�p�~0�.�e��S
��ˁp���:���wZe��8	��2��|���/�e�G�޺N�����2nC�'E�{�l���o���$�5�4���D̸��L�.8/�VzH�!
A9{���Jr).�4t%q,�f�ځ���Q���͟��^+�]y�޸���q�YR�~[X���M(��3��,����ϴ�,��vǓ(�Ҵ�|	���"�� l�^M�%����+��'���ǖ�;����KD��.��7