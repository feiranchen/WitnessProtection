��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K���.B!xW�����4��P\�T"�8O��y��_�e�d�E�|����X��Nfi�鯸ARx8�\zd6��d��'	s18�Q�nB�l�H�3/�ݔ��ES���ɩ�e��\�h�x�����x�e��L�7�zyG�����G�m]�7��ľJC8	:&b��1�ۃ���$j|� D܌o&�N��XHl��9�M���d����o@�g��*� �ԇ������B),+�	�����SO���h��F,�_�0�k^���$[7�ao�JP��"��̫��EB�(��Jc�D���;S�����"��D5�����3`�?޵�~]$���bJ��\�`��)p��s_lHo�)L��1�ᘮ��d��99.�#e��p�t�:}�.���u/�*�Q�o錿.9�ӆ�H� �vKHk]�J�n	fQR狤��}�X]`E:{>��L�p:� � k��3
q�Z!*�3v�1�`ҋ�.m&W�oF����&�\A�J����'�}�	�(��B�W���XR9wO݅�֚)�29��ΰ~�&9���u��2߁����T�yO�����>��� XdPr�&��̀BO48�DP�arx�På��;־d[ބ�o��nlބ	����7�D��%xߏ���v�����:�f1�Z/�����
94�֨�ͺ�J�V�V�~ld�AC�����q�����L�\L�H�w$ߟ��=$�\R��"&g^����|�|���\����EB�Uw �SE��]�u�7ڬ��y��3������T�)"�gZg�fu�g�D�"�6 ʛ޻�2���e��~�]0�Ӵ�r�Ł�bޅ�p�')��SUT��iA��_��n���z$�Nϱ�,6}�Tݓ����~���15bt�����JQ�d���?�U������i���KU�,]#��\#k��ݐM�bB��u/ )��!�'hQ��؛�;�Z`������c�����O������y�g�tw��J����ɐ��C=�4:�-=O5�1��w6�aLO�>��p�)��y+��p�#t�������Jfִ����*�]��j�㤩7����T��Ο &�D�����2���m�^ ���lJ5��������R�=��]n��������[5C�ח����eʼ|jGom&�IȈ��I/`#=��6�j��v��}4ջ�jJ�r�Pv���>]Ĭ��L�����S%� ��;!�&�I���=��r�3(㓩���_b����?b�MN�~��$�R����ʌX��"��V�1
՜�a�$�0���V���m�v�w�KN)̓籓Y�� �p�E�[u�<�G���u/l�p���SE=�6፠ 姚y7�,�^��Ci�I�K��ڢޑ�?ي�#�V������d[����[t�@�I��Ac�qn���Gӽ6=�ATA������;\���kL���Y��F�F��.���p��Ҍ.���F]_��6���+3�s+,�#�ݪ����7k�� �(��<�^�3`��j�i�C�<ϴ%H���;��V�5�I��F��|VX_H�u��:�n8�[.�K���\��� ��b��R'�G��{��vH�{��ڔDS?0̕��[ �~:0�d���h�#�4�&و�����t޺ ;@l`��CR��*��g� �7f��z�=��*Ę�����������̆�b^2��/w�osKf� M5q�qā6 �����Q��y�l��C��~P^����A�H�lr�d���]o���v�!2`>�ȴ	oD��}���f��Ă9��K�%Z�fH���ɞc)N���ƾ�����-���|��wAg y&��&��&�t�x�(&G�B��{�b�3!<\0����!/�ȾԸŭN:\�e����N�w�X���}*)&:!�W�»-U��Ux m�r�'QD+�E���>29�� u���j�����Q�����j��D�cRx�o��F����x��j}��)�����X���w�Z7��r(8�0�՜	A&�2p[�F} VѴ�A�.�͓�^i)G8u�&�؀~Hk;A�Pĝ�>3�h��֊��E��g�(���ו��Q���q�g��+dd�#�W+��	#���}���OQ��o��p�*�ȹ��Xg#�	5�g���8wT�@<�xRB��N��k0�&��w�:P0�+�	�?��Y�����H&���a��KL���� �}ݐ��%r��b��r-��Ӣ��z�&����� ��h�_���P�;}�9�B*��}�S^+)��*�n�r�ߠN�[���[<�	�_��b� ^T =C�ŚJ���Ǔm �5�e%�l+���_,T�R��b}������I��<�&�U�p磫@Y��r�p(alx	��6�����N��℔�b����~<��i\w���r�:�+4%u�F;J��G�O��E-L^�M�}iA����Yj?W�<�`�Ty�T�@��#��|�6K�W\MJ�<�p��'���W�	<��G�\��x����+u}��vw�W|��.0`!�;��SMՋ}�_/���(o�P��[my�ڃ��7��ʓ��i�ֵx���=~p@�ͨ #)�5����=I�����aHgYh�!����Y������P����v��<ͼ��uZ��N��!�p�Q�W���:��_q��� (�
���Mn�0P�7~���dg���fq�@�e�Y#_��Y����Ҽ-���d�_�����m�h�s�X��VDC���
ÑQ����{h�*�=�gc.�����}�s��Vvϴ�2�F�T�q/z�@��in >^IR�m��wp]��8���Yi�m��O4�?���Yg�%�P�Ƚ ����~LV���qo�D9H�(�Ԩѐ��=�TL)�)5?���'r��Սum8B�[��R���ߑ<'C ���-��`�Z~q�o� �|$�}We%�Yxh��8�j������b�sB1�^yg�7�>����ƞ�;:�	�!u8cZǈ��Xi���V�(ڌ�h^_>ռs[�2�6�$U�h�3��)%�/����w���V��w�?��.k����*E4�e�# L����'l]����*�6Ԧ��\T���򴥘�&�F�����)sT �k�;ȟ��/�����W~Q�����^!���dE\�J�a@T�?���3�y�\X��;�\ dN���~(A���=�,v
�G=��0�DNؓ��.2�=POm��	{v�����Φ����e,����vq�� ��N>��x��l�:e�ic��^��C�#�&̏��u���E����d�el|~�V�OIq��4m���p��S��QR��m���ǆe��nns軑~+K���xu�1�	F�V_B���͑��" ��?�d�(��7��#��]KMmPh!�9x�<���ѱt	�_��x�C��o��U��%O=l2�n�gO��^�^6A������]��c�rN���m��;�k���'�M�]�w�s����f?��d��O���3�N��q�V��?��B���m�!��"Gt���F����y����V����ŌN+VJh��Oa/�R��Q^��s��L�̛�À���u�� k��ީ3#���b���z���9H��\Ñ�s�>��IQ�����)~z���������.�q�,�b;+�x�W�Y6 ��^��mHK��m��ut0QG�����I���A| �
	�m(��Ֆ����<�O�3EP��k]e����1D�J��&��ѕ��b��N�a5;�z}��k��y��ģ�&���V��QH.-�fM�q7WMZ @�J���%�y�g��Y6�'=��y�Ɍ�Q�&�KmÇ[��;ѓ��̈�CiE҅�P�Y��r���̕�9��EM��ī�����`�8ba֝�>�D��_@����N��!�F��S3+�qX�7ߘ[���<��	�ӺTԘ�O-Rے�{�+���~���H"�_?.d�x�ٕ�q����}u�	UD)��I%�^�շ+6�����ʴ�t����`��% V3nK����J2�aaq.�;�@.�b�p�~Y&��r����/P�%ۋ�츇��׿�PO#��y�8�W���wG`��nN`a$@�%�0�m�G�"���ۮ"F��X�Ӊ&�����ߨ$���,�K+�4˷V�^ٞ��.��U>�I�ߑ�{!t*�Cd�ɳ%*��fJӾx?i�ǂ����?�Ӈ���`?�W�`��޷���_�S�!��oZ43�y��R$�7�������k-�Js7KC��_퀛Y��8on�V`��uv�O��5ݷ�&���&Vaw�ABz6�﮿G
��U��&����U�:��^���\�"��i'��E��=����D�*�$�Pt�,&��1����?�����-��}��S���,v�(9���+[o��].������J�k�>ZT���j��}`�7U\6^�g��p�е��s-�h�Gn�/�9w�D��'�!��*���]�C0>q�{�۽����
6m�O�O�-*�[��C���y�;	���~  �1=�wq}���#L�>��o����B.ûK�7$�h[��i�h�a�_gV�YA�-$d�U���y.��1�uAWA��A��C� s�����_N��Qׂ�����܎���T:<5��vЌ��HY3�="�:�8(b�T[^ʾ�ZP/S���>w�:B���8�?��N �X����/��k�L8R�~Nj�����i�#0���v��7�_�Y�����_Y��/�
P����[M�,��7/9&�*B�q�Ŀ�B�`5�c��fW�2'�SL��.8(��/��y���R�:��x7Jl a+�e��gy�FتZ�r�X|�ִ�m�7+J/z�,��151٤���Pi���,�� o�x��ͣY��-�n�'�$��j�V����(As��,��]�ظ�t��bb/�q���p��f�o�T�1�*��%ޘ١�k��Ԛ�_�$/HT����l�ǌP:�t�{�D��Fa�v2[��Y�e\�`#���K`{"�\�1�b!�چ,;J1N�T�-�o�$'�r��&��~~��?[���Pm�Vca���	W�5���O3~�_0hZÜ�1;M�Oˆ���jk�h����yN�D���;�L��̓����O�(�ށ�@�?�����d�?Q�R�`��i�毡��vsԩ��f����q��ɝN$����:%��/�^tzt I�pYJ7��;�ζ�'��{��y6&br$��i=dW*Z��61����*�����	.[�Ơ���L����h}zFT� �9����8A�^M���<���эEnL"�������X�ލ�����:��q�U�7�+��l���-
[F~�/��`d�� &�a��|>W� V�}����%;�����t�7_C�|�K�Y���mO������vQLkB
�W:k�v\�a��%Ҽ>�������9h��Ge�V+���'l2��.���xȅ��D���o�b5<$�5d�D�F����?.�G�(zQ(I�LUfK��ݎҊ���,'��ސ�����|���6�3�˹����s�sS��u����\�V���y��Aaf��;	1>Qd�^VP�D�̦�h�pQSQ"kȃ�t*5 �	�-#e�ul�iToTJg)V��P�ӈ�KZ6�ѰוÿL/N�L��[���3d`��d3d�<�ދշ�l�xs�Wr����oEKj>N$N_�/~$%F� �*V�7�����+�:��ku
��Q�I+�6�r �'m��/��L� ؿ�������1z����Dh]t�w=��Ȍ)#|��}y��ӕ7[��ěb�͖
ӭB,�E�[inP���Q������:']��<F�ƹ������N��ͬ�}Ĩ����@	�Zw>��N�s�֢n�1;{A��>�G�"��hR���ο��O�.4f��	8]�\&:�^�2��[x�6���΍R<�LW�-X��Jw-����v��8�m���p����;��9���*�������ʱ��dRs-|�JAъrE�C��O��(��r]�T���E�01I��'�?��0�O�kqUT�,Ywd�(|�I�/Ԑ�E�	�T�
�K#U6�^���\��;�(Ϻ�ea��¯��Y��Pb�I�?�r���'��Q�".
��_������a}��:ʫ1�����1���m��j�R�	+�^�����>f��O3��*�+u57��\v�����}52�����Z��<�>���Qf�oF׊)��8s'�SPu��:�H�L��(��y_1 	��<�)UjV��m�H�^Y*I#�V�	� k,�Y�.��׬�?���>< �?�o"������K% x�//8�B}���휊���
�)hgg���0V�c5��>�J���P%�`�8&.�^��m\7@���/��f��jԸ�]��$�nY����\��QM+���U����S�F��rp$�$E�)zE��?���$${Z�.�4	I]���#(`-{��y�zH3<�x�ײ70;Y5�'k��Hգ1���� �}��s/3b
.	6.mM1=�~�P�ƍdn�p�48��&��vv�̅�B` Q�U�ڂ�|*�.���؜�0��ӢqZ��ٚ�+,����������XiZt�n�&�rU����u�������> &,o�y�e���&f���>�q��i�7���0m�%��e���f��o�0&Sz�Y��CGn��*Y�	3�Ź{�n��|�1���,�Idȃ~]䂉A�G>�8�qfc�@���y6x��,�H���Ae���{}��}��j��+M��þ�Q>5�?�1��H�%9`֐�M��-��������3�^�Xxڝ�mL�u��5�0;���#I�@(Z�񸤤1�$�=
��Vؠ�{TC�����ϑ�N������ӛC��	v�h�g�Io?�Dh�p4g�̖�AF��'� ;9�H�'>c�<�'ao��e�c?lO<)2ޛ�g���W�pr�r�,A�)(*A�`�^�q��v�,�O<8��7�f���LO�T�g��8���y�19���0�Z�c��>ЬBό3yaב#9e����V���N�R3�� Yt�?(��_@"��*�T�&���=���x�T����W�M�ؼ��d�@�[\��!ڸ�@�a8ުM"�<�ّK���^/�	EC�Kw�ҁ���´�,�[��Lt�Y��I��H'���A����8Yhv2ή�2n�`��?)Hf��4oV�5���NH�H�s= �N�����!���%�d�]�5�D���n�xU�^��f������Y�pO-f��%��[ßq� �[U��X�q�	���_1�c���0ٴ�6���3��� ��[e	��=�F0�1���&9�":s(��,._�/o��Gp�����MMߡ<��s��KDOH�>x@L㍇��,�i�Ca������)��T���B��,o��g��xx�+�/㵎����$	s��Rn��g��e!O3Ս�N��%�����KL�9<�%-KtL��s����bL�y��帠B�fZlM���p�@�� �j}�����PU��"��0�D&�z(7��c'�i�K�������U&rC+X8UM���L�$N[���:53W�^�/$�h�Ȓ�쇱���_6��J#���\)�{�1T^��ˢ�zȭC�����T��h�z�F���7�]/�������������d��u(��l@y�i1� �Ub�m�IX*��(H�^�$e����+zU
B7geŶO8`Sh���*��ow۹t��>�8�B45�-̷��)$;Y��Ԯp[���2����j@��av�u`p,c\����y�1�_��♤�.t�[=X�}KS�f[ٝge#���A?z���\���HD��!)��P�h��E�|��d/�&ÌT�d�&�:Ϟm�I��o�������u�fx���4'X��
�������Z|8V�8ȡK���yx
�9���1�S㏩�%~U(mH�סO��M�st����\R�v��I�jY9�z��F������n�?��V����U��j�/��_S��+��<���Xm:��pk묓�`���gJ黄����֤�y�n�?^xmnr��[v.#��b�r�;.�4?xqZT��a�z���^c�$�Ue+@^��o]��ARR#����e�(r�9����
kv�?��OߗkdEn8ı�Z�f���i<bKѓ"X��������R3Zek\�<��q�;�z6�<7��P�\rA�^�YG��=_��!���0L��O?V�'w$� ���a�ր��3{`W`���:��is�έ����Ao?�ݐ�$���6p��`�K��%�:!�
T����/V�^��sx�;�kD�l��Z�(��@�į��<i��^y��ork�Y:����.N��lO�Xg[{�M�Ř=��x$��}BZ'n.�b"�a��4���X�N=��)�n0��n).O�+_��Q\��5���E]�X��2	Z-����weSW�c��̍`�
08��I�W��8!;�4��j��$	�ֿ&hdHp��E�'"T}��1�2n�:��$�^�eU��a�c�rj�5N00h�M�S�^n��#�X_~��=���l��|5m���Ӵ�a���g�-�޳����o�[��S�Y2$�PR��+�d� Q�8�|�`��tt�㞢ہ*3Ɵ�3P] 
�: �5/���:�	��)/:�Ф�ȼ7Kmn`Q����"Fm%�fu�)X�0�������h��/>e��t�vz������w1Z|��{|0��5��0T�c[y;3�갿���I�25�����wJ�~z[_u�Ck�K���R�ܓ���5���6_��ŢRޜar�Ш"ۋٽ��9�����R�Y�.�8��z�%ad��? ���)R��?=���w�҂�*��߶�JQS��R��A3�=�܅�rsR����|_��_�YPz�.b�o�����k�w�W��Hw.���?7�Y�e��zh�ta�AR��Y9�G�BV�������La�^���$���\��صC�\ŧ6Q��ɬw�a�i�;~-�~����
R7���@l!�^X;a�{����H�W#��j^I��:�C�t�
�0̕�a�ˌ$&*_��IHx�M, 6�9,",Z$��wRAOx�z����}C�h��+�$�����iyK�R B��
�j���;�W���<}^|���Cj*O��LY �l���5�U�-�@���j��4Qz��g�/��>N �9��F��u`{�4�4b��F-rE>lV��2��%I�}���Zng|�oj��s �_�!HXq����3��?��%ZSs�L�&m���6���*#'l����й���uL$�(ܱ�>_��Eؐ�f����]���h��G;S�Z�y!�=Vd�"��*D\XƄ�Jb/_����ؾ$q-�˿��f�2�[:
���2N�Q����.w���I�6[�Ja\�Ӓ68&s �[��GH߾�W��������0d���އ�D;߄�Chp\ﴴŴ���q: ��5�Bf[�~�n ��I�o���H��P�9���K8n������9��b �P�(X�+!�g���${�V@J����&�B1h�Z���	�l0����᭡Si��9u̫UMݫ�8$,�I�l���E���W����/Z��k,ǲ�.�����Y���I*�b�@�E+���r�(��r �*-�.L��d
:�w��A�]RhnTu͗x�y�{R�4��kwk*{6M>R�`�����u1G��_Z�������L̦>�ȑS�F��%9Eǰf���l����:�swڳXQ
-�̰yf�d�a�����0�1���&v�������H��n֘�~��V|i�����F�<�D�.����]���"��-��-�"w�$[�@�=,cn��]����H�̒�w��
�����Q�0�f��
�`��X�A�׬,<�Q�
��A8��Cf�3��� @�}�I�p��d\A
8�!^�����a57aK���6��쯇��O@�<rO� ����a�J�-)�UҙB͚55_PxB�F��*WJ��R�=N+bK�m�m�<�M�N[��������s	Ë�5����'� ��v���}��ɫ&�hJ)~���տ��w���Ȱ� >�;d�WDW頉�1��I�p���%2g���5C��ŕz�3�b�u+���x#���a��yR��2�s�{�8TKk��]�tׇ�_-�_.�����..�R�r�s�p�9�^��(�+h����.��)���o=I�hH|Ј���u�y"�W��0�cA�f}���B����o7yb�w�Խ���$mL!��Y��dt�q�#i�����Gz��Ikn��s�b_�x�m�lb2s��Sgc��z������t����1�!�L���l	i!�ق��z̧4�CVD@��/�ud_��wO�B�+$"�~��'�t\��2
�}�ѳP:�c:�B��C�\N��3�[͖FQc?�V���8�K�P;;�^�6���E�q~��b�
�9m�k��9�5J����V��Rى�Rp6I�0�4�Y�c�����X-ܚ,M7	�=�6��>��yt ��V�I����+bأmV|Mݯ؜F0���*B�-Su�X����i�.�)���Օ7{p|�
�u�C�Qy��`u !��EK��!�4*���!	��%[�\E��[˾��Q�h�p�WⰊ]	/�O~�j�ERa]��L';��l{	Wk���I֠|f&�[�.�xԟ�K�T���Q0H��"�UK��� -�9��J���Q�UQ=�[�Z�k�l�[���m�����]�����n�_2�_�f��^�",ӂv��I�Ȉ�W��1ts"I�3��D��s�I�!�Uæ�d_ngN��lR�\��!L��$�X�l��۸	L��R5�ش�;�0��j�,t����s.��)O������(c̡J_�S*�r�߄DyU��i%���خ��U,���9g\#>5>�b#�i�yk�p����I�� ��{�er	�1f_V��vp�N�;�,�π^[2�5�5��X=�e��/��#%GsW*H�N �C�ߔ��
�z�j�o�I������j.c��*79ݿ����d� ���ڙ��岤�Ū��x���0���eȋ��?�BN�6�o�������SJ��!���=�����e����r/���nVܷ��z��|6���������\�_�z���7w �]j�@GF/g�㉈�F�3u8�v��� �n�m��B6,;�צF/x�9�D^��ܼLS�%&0��Dd����p��6H�?s�h�k��t�J�J3�G��]6㍮��Ws߆m^j�aܗ�k.�{;�@4qK�6<C�ZGb�_�?f��������6e 	��7G�rK��?d��u��8�;rÃ�ARL��jM\������p��+0d��P�K���=��Q�"xgM�Ȅ^�����'���d��y�`ڑ��^p���bM���g�7<���l|�+�/��7w$�1tſ��(��5R U��Cɉ5{�#��$,���dVQ�c�r�n��k�\�op�95�]�k��Vco�~��!8iL))�������.�}0����8��e7�����뻉�JV�C��I��msdl}��l�O����H��\�@��P�T�$�6�Ӫ���yM���d�G�:�N�0�n�����U��x��:8Cf�o�����������᪛��K���������,�����F�q���ݍ�t�%����$�r\l�6���S�n�c���O��}}YX�ߏC=r4,�l�O����v�S��}=��*��6��C@�JX�a�\"�}l�Z[�6[�;���֦�(��r|��߭��E�`��9���#�^��\�'�,��w�z�X���P��kC*�Zf�`�#�~)8���A��!�	bgժ�RjER��E�{��lw��$�;�~��f�������&�i���~�dPT�r��_��ΐ��P��e�xqΎ�X���Qg�k[U�׊��E���2�K6v#�UX�F��G^��I+
VO��ո��>����l�|��w�O�]�2j	��^��rly-X�4���� #�q]��@�Wq��%9I��\L*r7�6>9�?3�*����ŭ�[�|!�4��q�����x����Fd����s;O_��`ER&N6�-�a
D��l�!�a�iE���Q�jZI��т��nr�"\���L����U�ɮ:�/)����"�o2�o)Y�,?�_�n A~v6&伺¼���n��+���9	�}NMKM7=�'uҖO��.���~��h� v\���~a
�XaoS�����غX��V�y-�Q}$�,˿Q�'���W8m�Ta=��=�[0\�#�_U��-
�Y���E[)a33�4��v��l��>D��*���m:�qD��"��0��*��"@C�^��n�0"S�Q1���$�:t8u9�R���*Z�h�ug�B7��G�����fP��g�R�A���D��NZ�G���r�F��@onM�_k��~��d���\��c��ELO�n����:��![/�1]�_�u�b0�l,�O��o��U]G�Ն%5e�qG��3+{@כj7�|nP��v�VdM7�W��By��c�$Q�K�3{��k\��.��f9 �zOY7��gkF��9O��̛0D��?�C�F[����畆��{o�lG�h��Bc=(f�
��؏3LzXm�IP)���G0G����]f�Λ�������W��;�Ɏ�SΖ����d�K[J�:�3a��ʢ�i��	A���ܒ�O���nL��U[�vF?��A!RvQ�O����;2�����_����lp#'.6rK�V���L�z�q�wDc������/��R�+�Q��:���C܈�z�~��B\��=��z=`�X-��n~��
f&r�?�I3�t|��?����������<�a��x�W;�����XE�����������H	L*c�'��~Ҍ��g�\{�����S!?&��,m���RFg�J���q�=E_i5��7�������j(W?n�:����g�%t�CG�b�Q��	Ѭ�2�k�$�l(���w��1�i"p��Z��.�V��S���'�Z��VdD1��� 5�;�'?BA��1�O�d2R"'7�$WS���0k
Ɂ(��bt}���{�������by�����;��35Z]��	�� 9�G	����NH���b;�F�·Y_��,Bߡ����yt�ԩf���2BA�)Y�GC�Ċ�O
2!�:�db���o9�)��Ǜ�B��?�dj9�XX�tjRo&���C�m�����o~�F���](!���:Gf��wdH9�r�^�;�"u�s�YB*�����9$�f�k釿��m?g�L�>�S����2X�fg�s��m�F������F�ɨ����^��k���˯4lgܱ �O=H]H��I�����B���ܿy��>h��IP���h���Ԣ�Ne��^�d���U�������cq#�A*�U#��C���?J_F\ш�
��f(��%�o�,NE�E����E>�Ƣ5N�@�������S�i� W��'��/�`�x�19P�A���om7P�5�V�s�J������e��$��P�?��� ��#��Ή~���?4G[�oY���<B���n]�<#�%ѧpT?Ϭ/2�fU���̥U�����l
�	|���H�X$�&��x���.��~�)l�Тkmq2$�Qn_,Urh���5_dA1��w��_̧i;R�ƈ>~�N/�r�J������Y7��[
)�)��Nܥ��Y�
� &���F�'l�����+�E�07�]/�H�DT�	��)z�H�{/�N	�h�*����� .a���%�p٧��� æ����42�TN�ɔ��E�Rf�m趱�(�by�t�R'��#����C�5�(��$�ֲ�j��~?2))���TEԿagW�S����C C�ge��L�WK������z(hޔf��l�ڻ��ێYF����������Z���e��i�'���d��t�cv/&�ɼ[j{ q>7�{��$9C�Q`����M7xC��_kN>QW@V�-ED��������됴4���?%���{!�B��ɒJ�0��iL��#ϛ������8z[�����՘�OvX�ʒ��<!�;�G_L��:�� t`��~m�-��\� ���^t��S�@~��9/rDbT�N�E����H�����UM�J��,CEr�_��H*Cd�;gG+E~��D�8�
'}�zg$ >��[�����'�r2X��~�7U���|���4Oq?`Wo�٘9[���X&�A���A�ڞb������SlB�B���K�
���8��P�x��U^�8����"�0�o%p29K<�������`D��d�>���
��,4�\C0|J�h�DY���1�L�C�ș��/mt�:ɀ0�����y4�w��K��R�hÐؒ�i��҄goWӬ���������L^�P����2���@�r�C�Ѐ�à8�Ĥ;ڱ����F�ڮ���m�S��-K���֠�6�R��夛�=���s�j��e��>6�
��`_�;w%8�,&LhJB�UR��"N�8��َգ�N����O���}�S}�g�C#r! !���T��;�Ի{ ׏Lg,M���ḱ5�p�2#ց�o�Wk�Ւe= Zd�.h��}/�/L�\���C�͆L*s\5�j�R��)+�$�T�Sq۽MN� ȩ�+�����\�g�:&�_?��Y�R�����j|��vi&�{5 �#��sV ��5���O�=o�����خT�|t�\~I����L5��v5UO�9�F���{���n�G6��1º�b:�æ�!/�G`��iB�(+����@�
�iv��@	'(R�2[}�Ѝ��L�Ϲ�ѿŊ[Kp7��@;��U�p�@�.���B����҉I�L�AG�Z�.L�|;?��I��Lؙ�=��$�|o%�ج�MN�8����ySJ$��� 2��L]"Ip �_�d��]^{�y��r�{��_��@�p������-=r|U�1U��nd<��/���;gZ�9�j����ڸ��*�n��N��D�b�����Uh.��m�-/�<����JM���ƌXg<dNH�:�(�m!c!_�ŋ�sm�S;9�i#8���"��ۥM�N�Q�cbޓx�*��5׺�} �,���P{5�R�X"ԜQ�SI|"���Z8�!�� dK���W��C��>�,쨟������E�S��L�P���f�/~&���2zG�f<E���v��ǃ���k�H�.x�ͭP��7>��K�,�ݝ?<� �*����ot�{�+��p���p�V5��7�a���it�e��I�nW�6B��Q�#>�{��mtK�"�^8���ef�<�A�5�/�b`F�0�)^��Rڱ�=�<_�$���Jow���[�/��Q�IF?�:u�C����i�����s]%s��"��ǰ��PJ���z�K�'�V�����!�ڠ�a܀'�goљ�b	��շ�ZgQZ�l��T�_�2R0.� Q$Q�u��� *ݽ�9�:ܱ�kI�zM�A��6��mz8��r䣱�;
٧��c�I;���z�A�"�1���pp����ٺ��|�����Q��PLM�G������,i4~aHos<����a��D��=��Jo���&�Ԣ���
R�,�T�V&�[m�׹�sK2Ee_����X�Fpf}:D�ʄ��y��gC4}?d��6��m�Iw��v���ֱȹ6)A|�X\5=
��s�	���#[�]������núɘ@�HOӂe��<��t[�<�Cxy0�8c������	��������>f��������{�}�I�>.�g���X�p��m��5��W%�P�J����O?���e��M����� �!����"�eچzVs�t�%�U%�i�[��t�ڌFZ�D����&F'����B�o�ڌd�t;�5v�V��8�f)�HM�����_��l��j�BY8��l�n�K��V�����?9�������D���+��b(l��~�O����du���S���`Q��j�i�ͶM#�ܠ W��ѕwP)@��Z�c��4\C��;�E�A�y��J(L�]WQ���æ�s���V�c[��%:F�1���] 0����)���V9���K��$V2]�v� k�{���2T.����4#i	��%���F�4���Ő�l��"T�.P�Ll)��L$q����q��؁���0:}	�ؗ��Ϧ�=EN��� ���Z�*c�A� 7�ml%_�� 6!(X�zu&�'���uj�c3ɸ�P��f|�"�ԫ3��V�
�T^�xZ��Ut��aP4�\��cdEȱ��
�O��1N�@sJ�/�eP����4R������5��|%d�d�6�T�:�qP�K�ԝ��_�9��A�>ND]�TI �Z�O��'�wG�)?k�x�=d;������Y�,r�_�\Fd�;��~�,C�hGhe��%�!h��ӫ.�	�2�IQ���� ���y���׳e3���K�?��hN��T�-�ֽ��݁����R!�!�^�w�_�2Ka��tw�Y B�%1s��2��R3�&���5���vosY�J"+x��g����iB�#s�W�>$�U~������Yq��#$���iq\��/�9��l+����Bx�V&d�;J�,�6�bfi�s��9FW�S?���.�9Gt9��s��}�?��{{�}�9�m-��wد�z�K�Y$n��J?~�(o��Y3�'5�V���Q�����K�iC�B<�Qߢ���#^"�ʙ!�l�m�G�~^������e,�Y�:�6MU.�e~h&k\C(k��o���UBvYi.�BS� ������ܶBD8q�G��Ue޹P����(�6.�{r�?8�u�x�D�N���A����P+����[5���UU٦|\H����0��P���]�@��4s/
X�I##����4�(?�j�!��F��r���e@�,�a\�rm�6�솘D��{^�<ɗ�l�$�|����|<�������c������#���U� �1�:Q�,ѕ��~�7�HT���<�O��"ep���	hE��?����wd�V����(=�M��t�/�'h�OZ���������Heo�`�m�q13�g��A�(���N^O6C�^n(�0�L|�����{f����g"��5�:>��`�ʣ` �� ֹ׹�� ��~��\�>b:'�a 	�������	m�6<^�2�(kCh��qh�Tn{ǻl�f\3��G��f
���.G����/��X������[��Y6�L���W8�D"8�e�j�{q���� _L���AbZ}���l�ml�P�`�!=ʋ��S��w���zӦ�hw�j��n�k�>
��P_�@5��ѡUc~��-<Rm��>o�Z��CX�G��**8�),��3�fR���$PnN>1��変U�RH�a��0uْ���.�Z�6�3�DD�1sГʯ&��!�:V��{��oA	�*G'�la�k��!��$l�4&�{T�1�3>N�Di -0�=��2�yk^����M@#z�g/���Z/P���@���5����e�y6�c�>��.�"���;�1f������W#�����c���Xl��L���L���0����)�s\�Fʬ;j�HT<����Uhg���X�'�Y�8Y�lȒ�1*o�i;Ii���Q� �7G^��r���?���%�[���;���z�z���j��3��wC��q��hq�w_G.�"-��n��0$�}?f����o�x��F:fx�L�Ky�b���n��q�~�Wx����q�=�@lV�C�̿���$��h�����V5槊F(n`��`|���Jb�3�gۨ��Kd�m9px�������u��c��lv�1�8v�!�Bp'�*��2�tq�sk�����SH����r�P�A�v�~�z�GyJ4c���NVJ�;稦�%�G.�r3K+3��,�	���s#�����õ<���2}ߐg��������iqхd���\1��FU��o�H�p[Kx����' ��~�j-.�K��˘��B�����h�{���ɽ �ɥ��.C�#v���R�TjKܰ;���'mm�j1z���d�BL1�B=Љp�j����fs���{N�S�Ex�h?5���1,LY��� ��M0�8͢jP��䐰�낒����	%��t�� 6h��Zr�S�:��S�Mh!�j:�Q`���/=�$�د3���A����ƏgrQto�z9���M�W���
�{cn��iJˊ�W���.�L��>>�d�r�����H'����fS �^�8�r����'�U�6nZϜ��p	��d�����#r�i��T�7��
�7�4��#�$��5���s	_F���ّE�Z�?G�#�u�
���<��]���	��ΑN�e�+]�U�U��e��6�fI�hC=6��s4����"���Ѿ����
��_����VkP��+�I��)��l��:'�!`a�R�{�!�Sb*��Vx�^��&�S��~�%���
��	��4`�lK�鏡�����`{�zfp�K�;�n��*U����L��~�%�e$�$�;UBz�D�ٕ���@��ozp�H�o�%6�q�]eK!f�?]C��
�~]#;��J��E�1Xɖ�W��g�^�	�C�B��� �pGI\[{ES�ƹ̴]��s%�~���^'�>EH�3��0�|�Y��p������p��o����}j���9��B���o���iT��K�_~�Q�i���+{s�����뻛{aע<�ea�;JЛ�:��������w��W���Є�J���
^�dgŦ��E^-U�͚q�ş�w��J�j���jG�PO+B
�ZVg����^�K2u2G�w2�|�c�v��7�Hm�SΫ4�?��ı 	��J4���4���
�l�����������^���_:�*�[��{ �I�q^��!J��6�_ê��Es�!N4�u����v����R������y(#Ɍ@|��vt����&Uo �J�^:�����V�|���y��ͲY��l6��@���>���	�g�|k�1�q��{{	�Q,m��g5�m�j���Х�Wm��'�	'����rq�,�N��d�fn\����B�k�VA�hӍ�|�S�ѥ$�w"��YMh���b}�UC�j6�0�;;���2��id�:(���ԏ��u�������\MH"�'IYd}I�`8��ǮŘ\ᖚU�V��q?��#����P��Ҟq�p'�e�Ñ1u�[�G!=\��?~T��N�x��P�,�E<~>�:��bє���4��*�؉y�����x��)y��s�PW���D�.1�
�����HX�֓ v]�Ǽ)h5�?�t]�����v Yk�"-��STKC^����)S��%�x����W�xM2U��LQ�e��&~��$+<�d�PU������׎��ԫ��,f�7�SB��;�)��~X#1���o:s*i`1��c��;[�܇-�m����}�V����'��|��B�j�?�PB��ڨ�66�/�`
��Y�"�p�?�SJ^��ϔF�[cX�Z���h⿐�&� �iJ�cx�k��_,�ܥ�t}&z�ݺX5���S	��Al�e@���Z��S;Y=[����<D��#$��s�ܰ'T1��tb��{�N��D��KE}�^^��̓�nmV~�8y�89q*��-��$!�)}�\�Q�
��`v�"ԇť-���3V�B��9I�3>�&|Y>�������KkUuE��E�U�X�F(�Z�|~D�{?��p�u�}8	�.�<*�}���#	�a�A�E�����ޣRw��D(���F����I+Vt��6�C6����-��W��p��i��='�:KB��V���*۹���!|�L��q��)�^�eF�P�f�UR��~���ri�&�/���>S6dp�g�x7Jg���`k]�װ3ǂ�����h&�/�a��ϸ���s��:�`���3�8p�5��l���P�*���	�9�;�Cu��6���z����
���S���"*ِ�?�ݼ3W��驆���.������c%�J�������B�$E�+N}R�'w,��HM+�V��KX5�k��]����x/_̱��}���'q��<U��.�����G��M�_����"�	G��Z/k�7�9.��il��9�䐗�a=m���6��f��܎�Ḻ���NP�|��$/��B%�L�v�X��ikv�
`�������� OCԟ�=���W�\�,B��g�v;J�1i��S���M�:���dS��	B��2H/:�t���[#�΍�#ޣ�57;uT�Y؄ل�9VU��ˇ��4�G�MҊ-Ewc�_#?����^�*��PFR|n}m�Ј6sC�y0��X�	w�0�?k�{9��+!�P�ǀRx:�8Z���L�q�u�x��{�:�U@mG��Z��^NvQa��h�C��ҡQфH�[{?� m�܇��m�^�wa�m˺R`՜<���|,��Lr(ڟ���Ы�X�֦�����1�ChU�2��ۋs������Td�b�\+ʛ�������5S�٩��`Y�d5)�(@����Wټe[:�~]G4PHabQ�sKd_2�+.�g1� �������b��Z��No���b��vh�A�R[U���R�ZN���
��kٺĸ� ����D����'�!��:p_Y Fe���ܸb%�N��A���dx'���Zn�f��ʐ���l�1@%����ԣ"� q����{b�Yx��CfX��S	eъ�
�0;�4BƐ�{,�E͜�7}����I��J=;,��d	̬KKf"f+�{�k��2㱢�+���T������X�̮ewf�h��C�w9&��a>6$���n�=gO���C��;�,+��H��.�$����֝O%�>]�@дN�mE�$<�ELUt�2��3-�k��ܧ_yBQ�-?b�c�X"tI��y:O	-�������jes����2���-�������O����ӊ�"P��<��M�s�K�����l�W���&|�$Ōhա��a�Y{�*����@����5%��D�,U,tO�it��2�vޭ���d+WWZW�0��uՉucC�kK�Y��zn����/�R�����F�\�$��׼n2Nlh���T_ˮ'[NІ`�-��������^�Q��U�[1ɸ	�$�a�6���-K�&�ǲ%�[�}L$���<X,�gؒ�a�`5>/5Hx�#.�P=f,V�b<t�|}�.�l]&���*�YT��%��z%��(�:}P�z���;)R~�¦++~�c˦���J�����s���;k��X.�w�T���\h8���������\I!
��qxG@,�n>��d �l�g��->���?�_�C�ۈ�@T��������J�.��e��^�$���7}�i���g�r�X��� ���{)Ta���m{�ȧ�R���r�z+���.<a��q8��ሺ����#}�뷾a�ҹO4*7pz1�B
���P�1H�q8>�1�
XPC��!���I��(�nmm���w6���טO�+�ӷ����K����O �((��\�+�����(���5�y*�	@�z�L(�"N��,J�.e'V���-�0���WU�=b�500lj��a�F������3���OAa��rL��COs�vg�f�R%B8:3���(���hbnx��� �Y�xF*��&��B�⢞���)�	�ݲ�=$rE9X����8�Pk������ɶ�+��_D �J_�Ֆ�0���"O�io��x�J�ٛ.�.�W�SK�X�]�f�s��u�BpSl�<��z��xl�5��t:���gI��ZQg�</vHi!3l�2<Rw�;t�B$^��!\����Zq[4�2�iّ��U��D	�sop$���d!C��r�O�^M8��<m=�QE�;��'�8w��a��l�tN K��G�� ��6$X� �1v�⹸��uv/=����G�v �4U��@=������3�L�R�f:vƮj��i�|����L�rEPjأcU�,��E��A�JX�R�4�;ކ�G6�C�2I�1 ��h��ś">;�5tЂ���W椝*���?v(�hë෤h���R}��<Ҍbp��+��;�O�r��K��<E������?Y�Rf�iN;�L��u4_�菮gz���$��Z�JlpE�љ�^��V"H-���UF�ji�wDv��߇�S>�UT[(|�v9['�f�mP�ˀ���)�ri�<�/����C���u��̟~3�Ύ����/N�������-�xŰ��d@��Z`��[��k��܇�|6�",���@����Cw �1�Ѯ��=��x��Ԟ�U��i̊P���n��|��+(�8�Ɯ9-x����)�D?:��/�B�9��:�14��Np�QDȗ���L\�\��Ep������b �w�*�\�
�ĖbSF�ۮ[�ǭ�n4e�B�^���4V�W�?��}��C�����<��X��>�;�QȠ���@ ä4Ԓ��b�l�:~�G=�N��Y�{�y�T͘�Y���)GC\��(��Dv�p�n���w�¤l�?�plW�r,!����EN�ٌ�/,��{+�!˒�C=Y�(�B���gTBd���C$��p�#�WλyU�m]���w���`�h����IV�jFEL}2GMݷ��Cu[��u�:���Uf����ov��@����N�
m�ڴ������I�E�G��:�\���9���di�޺�ќ�qa�����)��7Eg
f���c����C�.	�7!�Л�{���к�n�a&O}�7M�Ā�[��w�yS3���U0f�.�������+����5Y���w=w@ń�P��>��7q�L��Q��B��
ĜW�.�}O!�e:!�c[��֨xnmMք��%�ra,tO�-̧Yfð�$;6��f�Q�0������+��v?X�#C���Cu�*;���I�83��2(�Q@bxM��_z��s�1A������"���q��v�T�F?ɰ�7�B�rN\�������מ���{a)_�Zym�����BT�1qw�O�+�I�P^�|K���fV�*'��j��ԁHo8V|����i���* _\^�o����Άƍ±��҇��1z9���E�C�Z��dt��8Ee�m�����m�C���iX*�ջ�U+���8�m���+�-�E5�����گ����Sr�1�2��!�X�.������U|�ܨ����Ԯ ��s�#l����8��~`uP�w��n��)��k{�Q-R����V�kfI
f	�%@��c����iO��5cN���g\���4v��E#fi%�������Oף!��׾&�)p�U��K�h�����"\��Ƚ>IѼ�M�ًy/�%Ss���,��:�>izj熡��}i�3�ƪ�0c���M��C������Ǎ��>K�42�PS��|Z���~���	�� �i*Mkm�H\��-ǁ�i��o��M�Ҿ.���ܣ+ X�Ju<UU	p��`�����|D;Lu�咎��xz���#$��^xz���/�|H{x�ah��x�
nUW5�\�"���	�i����E�c%��(&�9��5��jbu�������t�;��M�@̍p���]�1�K Lo ��������9�C�,D�`\"�T��L)z�Q�BG�4��m~��Z`ի4��MU��H�P1v�١Xkƪ��@g�,��xRv�\&	I��ED쮕���mrI��1j�GXZ^��>�&<|@��{�i��B��� ��\�eDy�����I�-/��W!SۚN�Gw����r�2�>~%s	� �k�*ݎ��S��iK�ˇ��ޒI���	ۑ��$)#��8�G��l|eHX(\pI+I���HV5��+��{`1#t�%��������:A'1����2e.���R����v��D��N9�T�ǥ�Ze���P9�,�(h��%��>�6��>n����D	�p�`��-v�n�FR�¿�����K8Q)��%��n����"�Kj��s��6˛�h9w��VJ������a`�y
���y������+��k}.1S�_NG�����C�ĸ�ʦ{>���M�Ӭ`���R�]56�h����ڠ>n#V�ʾ���!wdb�0>0����t�@�����`����ϴ�e�����*/�=��)�r�!�q�AMF�v3��6^�Z�?z���	��j߭Y=*�K��)�[l9�s���B�d�K��|/���%]�?a�j5�ki�Ru��0�~�W+J.?���c��Ӥ|1u�r�-Oy0;3axh/ڢ����R�O�M��1���
�nG#	L Ԃ����>#Р�T��;+��L: ���B_��C�s��T��,RߺSi��8��&���x}g��q���9��6�m�[ko�π1�E?{6u��Z?2դ~9�P�I�~`�oi�ے��}��	�+���+��E�{�lc�=g;7|�Q�-O��:^�64Ęv���{�n���S1:�9�֓_r-��H8�%��ν��Q"�h�ɫ-vF�e����_F�p/<�^@y�Jo\�2Y(�SC��Wv7f��t�*wͭ&7iX�n��wK"�ݜ�D���@�A��vm��5���؆�É�]�v`�ܝC.�ƣĥ����ƿ�%q1�{0?��e���+��PmGu�
�>�v���ۚư�		v�&����Gq���UV�-zkg#�ػ\�?acW>ce��l�ߕ���4Z���r�׆���<��˄ ���	跒�+��T�~��Ӻ��p{>�o�&L��3(��t4��h���&��5�����#�@b�O�Щ�Bz *�I�R �C�s&V�~�vMT}�ئ��1/V��&`��2ՀunV�;U(�`=i���?���Zİm�[�-�G�e��P�0�"P�>S�"�s(�E�
�2�����f�Pd��u��H�癦���N`/s}�f�M�1�.gFٹ{*Y�I���˅5?�,�~<�7%}~�pM���DVs�V�GR�ל8I���[_[�\U���mO���{쩔������mgC:ߑ|���c��=+�帉s膱��[Z�H�L �-���}C
l�+��$&"x���?�0��V�g�Z����<Mp��oJ�i�	��D�s�C@�w�����Y�2_�q�"1�Sݗ�ઞD��1d��Xx
=�o���l�Tџ)W��7F���x���)=m���4�@\���'ha�����nb�F��Y!��0�{v�kG�G�E��F�<Dg��7(NB
)�\�,%���yg�\RY�b�W]R9���a$	�i��{\6�A��s���נ]n2i�� �Y�"m���Ҥ:zq�-�Շ��*=�7�c�ǰ��RW�R�h�������Ln �@�],|9��rw�|+#=��@;g��x@���C_�M<�$�z3<	4X|��(338�S|�e����=0��p1�rW��k[�����tm�`���m�P�4������j�����x�RI�x�~�ka��k8�����	C����u3-5��p�D��Ɂ��%��,��~��7��fX��VC�`�'/fR�A�tnsΨ�1��K���¾f�֖9="Ƌ�g�6��eY⾜q*�LЭ%�'`F� �B+��(����Z�����a��>������X"�v�K���V�0�7:��S�(`�4H3z?$�q��b�	�k�`��¼;�R�*c�,��KVG�3l�6�/d�|�fjp�<�(�n�����:��:�*+^gjz�[�J@#+����M"U�@<B���&���F�p�j�#�BEH�&e���8j�!�X���u��+�Fޞe[AmIxn��栖^���ȼyk>^r��������IMï���e�U�-T����
��$���i�ޒ��wi5N�<[���@����<"-�I^����$B��cu�v�>�����C���׫�5�����"�{css�2��>؞B`�.>�k�є�S���O�S�v�'���U�G�c&l�(�G����ɤ?a�ZIn:�0m���D���w��B��V�4Y�wqȀ7��:<��z��J��jْ),�g�e�9�^�+��i���U�B��P��ÜeU��n)$0�H�[���40�j��+�L�d�d� �0�Ug<���RDe��ʾ:��i`sHҐIg �zjVx���1-�C�px��L���<YP�q�V�W$(���R��� ���S���P�=~I��V��/1����~���i�)KmM �8�}d)ΔƁ�Y;v��V�y�2���d��Rh��]���9���:j/�����R7z#UI��Cp�jH���k��Np��z�|U�˛/�dr��8�l=����1����ru"-,����W��6�wgtE�G:J���"�t�Wd�>_��|]]Ѝc�eH�(��j�;Ʈ=UbЭ���3��KK}K���D�Op4 Ϝ����3� в����U�.�]�b?4^'׽d74/��\_��Gtܠ��_�D���99����>?�c�6)Ed�-i��>>�$|��%�&̓�(�d��ۻ�θ?��g���'SU�b��?�t�WV>ڀ��vn/��]���-/�������F�W�f
� r�OZy)R/ѤV�-��Pڹ��,���Fw=�7߁Ԋ�Jf^�zRa���P�)���I��_v6�n�1�(Ӄ�B��sJ��U���O���r@�"Ǣi�x���I���)M�B�yc��+��/�����69�Q1YJ[�(��0ƠI�pL�b����(��פ��S*�	O�E���ʝ]�D0����/�ϲ�UV�.��,G�z���g�?���k�kvT�<3���ݶ����Q�/L ]�Ѻ��^�,�r��G�n��J�"<V[����Ղ�V��������~\��Rǔd��gmC�\��d���$Y�����P�ƪ��.�	��N/��W�,������HT������O�O�K�	p���*�MƂ�<�!���?ٓ��L3o���|dz�{u�Gt�O5�R�������z/�NV��#8���n*m���K;9�m�3���łܪ1��a�]c��#��k��][�<ɟ�E."K�V ����`T4e��$�	�n��ʗ�bS*s҆�>n7�8�nt�cD�5�/�zhE�M�zvQy�$i�I������q� �ڬ��跍%��!�{���Gna��:�~��8ҋ�S��2�喟_����z(8�7�e�d���oZsdN��������nY�:��Nr����om<��R8\�_%��q%x	�Q��v鏟�h6�d�
�����W��,gF�z�AW�j5�N�C�����%S4*�3�*{�h�J��@�
��R=i��'iUQ�H��E�����'��i|���ή��K-�V4�rƘE}���gX҂1p��N��
E9�u�u��;��Z'�����̢�(>h��kU2�b��R:zv�����ߒK!p#�:4�v�I�5�]���mGU,l[ѵ��0����cyy[�Ow�^4b�$�y�4y�F��4�'x5hL?;�� 4��U[����3��m��
Œ�XmX�>g8A�`VI[<qp��+�C�OU]>�`]-P�P��ZM)T抟�/O���]I�>7��
��!?�.a[�2��� 7H [�őn�=Z����Ӑ��u�[j�d����WDҒ]X�ψD��uɺ+���q�ŸK2�i;��dt�؀�N|�gP�����H�f��:�pM��o~9�Q�_�M��(�Ӟ1g�2�g�0a����DX4�jOD�(5q��L�$1��`>����0���U���r$�������^�{�R��&��(�$D]x� �2ڢMhm��֝��b:}�H<fQˇy����9͈	H��Z�H0b&fե%���lO��N靌�rX��y��e�`:	���h���$׬X���<~ND!s����m�B��G������I�ZD99��'�Hd8�Qڰ+�~?G�J�J뤗���1\���]��@5��\$� ���t=��!�)��]��rej��t����XK�A�i�A4���?:��ቈ� ��N;���Q9��T�T|M��CB��F�-��*b�s���J�Ǫ6"�u�V�h��M�9mUD��A���R>�����%|,M�y��ф��*o��B��~�vU��ߢ�*b���+���W�y�n��R
�x~���;���&+o�9h%/q�+zm%Q@"����MI��s�Z�U�f���P9�{��D��}E~̠�R�`���W!�b�����w 	 ��GJ�X})h3D�� -���H����ߗgK-4i)�Z�j6�a�:�7��tNڰ̥�P��`�s��p�fÑ� Iu��a$�~�fw��<L�	��0�Du<�p
��>����:�9-R�ߙp[��b��xy5f6r9sH��vm榱`�xâ�'��|�k�
�D�l�r�Rz��n���q�)�BV����=��Ɓ�,(u����a�������J�#F��C���Yx�%�g��B
��e$��l$��4����^ޭLQh��k�4�6U��)C� d�E��z�>ae³�6��hi��.:�ƫ������d$-�z�1\�\�(��m�wh��LyA�9EÂ~�4��ѹ�$�e�F�HKЫቑ&@03�6:뀾�u����Bz/J�lU��[�n���n{E������Y��*�1x��P�A����l� ��o�sށ��!�!��dîH�p�,����
#�O+��X�����aɭQ/�%3����fA�W��G�Y�4�
�x���c��LkV3������}���M���]�%)K��e�z��[ՠB
���k ,#�h��v%�?m����c//r�7�5��Iڂ&�IQ�}�G����{�3�	pXߞ/��~���<�ݴ����2
���ֵ,+\��eL$R�z#��G��U�Rƶ: A���2`Z�߹q�If��c��9?��W�Qt�͍��Z^��,�S��y!�vϖ����J�g��*�Chľ�ص݅��=`�J<�[K ���E M��4��.؃+`�T�4ZD��+}����x�<M�c�Ne�ꂼ�SF�*M^0��<;K����:L���O��5�m$��7��	��'��}KE�)�E����[���)�{�)��ԣ���$ ?�`ɑ���c`�7oK�&S�J8�xȲH�Q@�P��ͳ�Iy�#�򤴅�V��E�t�����SNAJ��8��\}z^�O!�WB� �T:��q��/Q`Ua�9D�]dOVT��<���L��S�-1���.nE��x2T`��c��;L8ؽ��<sBM�j���@Qε���Jw�t��Cc,����.�f��oeЭd�Og���+���fh�r=k3x��k����E�Bls9�����xk��UҐ��9Aݶ<�TȌqQ�Z��;�� {yL�s�ͮ��az�
�n�2���5�R�m��تeX����24��&YЃa�G66�ӀN��kȶ���V�q9J���P��H���rBȹ�1s�;��S1�]oU�NqG�Me�r댵��cQ/�ّ���JR5�EP�n`�HV5�q��xȌ�����dyI�5q�
�M-j��<5�t�ԭ��wƼ�b��F�9��tU���R��j�Y1H�����s$������"\ɾ�k�rn�~���~��)�K|�q}Y�+�����)������ͽ��A��12���T��38/4���h���9�g�8���?�G�z�=�^���ԫ��Y�f�;��rg�OE���hM}E�: O�M����r�����,���'�s��'��t�t������������{�\�0�<��@���"�z="��ց���ds���K���oB�2<���4K����y������o1�O�!��$	��VY�l��Sv"�K����p�{�Eב�E�S�S��!ٯZ����4���E�78�k�S������|�LC����M�Ϟ�E�Y߰E��J(	=�}!�V?o�<�pp�5 ;��%��ݮ���,�N�.6ձj�aX(�Jں���Tf}�����+SKj�$��@�I��:���qb�$B��Z�]/�@���H�,_�A�`<2FΧo>�*;�zYϟ��;���N�K?���63˅N����V�]!��{@�Yf�|?w�	�wm\�{�ޓê�WA���oN��#���FEU8D��K�N1S�[EΤ��r[1m��X���-1��ֿ���������� l�'v�����=9[�#�뢎!�M_%+�����+VN���o��j���K�Bc�]�����y��K��L|�D|�T/	���[ʩ�>�\c�Ӳ��p�b���͸���t����6�Y���<C?�c� �-���Ļ���*�J���T�j_�l��su5�s�H����a]�p�h��/Y����eq�����}���	 Q�D=����׺j���1Hj�����y��W2o!��np�̱��;+��oU��4J��tq/F��,����"���m{� o��	Q� Q�U�od�֭��\|[H�(�U�w��|Gb���Z1�����Py5�9|����h���@{���j8���}���QG�9��#?�8�cil(T)�#-��%+�:cn��g`�����)�!eW���ޓ�5��FZT،�F�d�jګ<o������H�O�f��ϳ��)�@���69�:��8g��0T�be���j�cb�̀�^�.(@�w~�]���S�4��t|/��K
j_+9:�;�\�z]J$V~�]�yα�.�6�)��LTmE%ű����*���k��c�.x�[nu�z�6�S�2����gNw���-���Ќ� �c�����l�e�]�ۜؖp�$������:�{��A�S��gt؊�+���[��T����+��>��"2��#]�krotӍ\#��K�I�H���b�`��GԬs�ܨPM�:���ˊ��J��ŏ��;`�d���i*�����l�����`7��<�f�8��H0�&����B����IZ9\�5yĻ��>O��y�M.��u��i	ś�VnZ�L+S�IWZ��f�J3�[q�}k�^���SD�HИ�&��,�5��D� 1�Qc�����FJ��� sI��O���J&F�YÛ�+�g� aׄ��K���K��f���.l@:Q��W�����J���r�3�0�
&@��� �%�D��U�|	���V/���.����F�a�k�/�t`FO�FF����s%�2���7G�8WmZ�#.��m�X�U��!���k�aE�)j�1:�/7	�_(<^�����A��=j/���L��#�dp����g<p���� P�!pJ[�=����<�,�fJ#6*��0�H��/�ޓ(M�,����@�fSz��Gѣ˴���-��L ���uRr<- �m<����Jc��k�6�Tb��� ��9ŷ�ޣ�.MA�2���A(.�ď���fH�-4���h��>z���Z��m��{Jt�c.�P���Xfh.���#�O{l�����u��pH�W�"�����<*���uI�lsp��>��D�$[-��0�����%y���e�����gn�2#P���)3�RM�/OW;�Ρ���4fE�`b�=|Z(b8��v�T$f��˭��iy/�� 5���qLa�]R�$t����ү����;_��|4�
����������D֓��GOZjn*�[S���/�'"�DK�>����N[�يbF$���pu��:
*��������Hw�O�3AX��C��/����5"0J�N���3T���|nE̀3�CJ�53����\ 1�� �t]�{F����`"iJ,��>�e6����Q8�7A-�����dz�uv��%����ђ�<�TO�|���E"ƽ,�&�)m���2m�C�1ٺD�L]�(����"�� H�rFs�_��[���Dʊ)�ֺ�sr��k�A
�Tdo~�C?��p��o�9g�b�������-����tl-ez�ů��ϸIB8E�1�l��&	�)���"U�2n���^"i^r������&�i���>���%�miא{7<UA�
�k����|�#�?s!�As�[�a������in*�׼��O���H��7t�J��Ni�����
{zL�H��#�*�� رNۘ�tP���LD�X~��9A�x�h��ϭ����=G�At�o��{ҥ�|Mo��؊Cu�0�LT2?Q"?`#��Pqg��6��G�"��n�&����3~;�IQ�0Qˆ�$���ZC�Ǝ]a�編���ʎ��$�m�`�ہ����+�>��!o�����{Or��^I����IV`9��y�{1���\��GA���ޘ8	�����ɫx6`��+ɹ.!c�J��_i��;�o��2��C/�p8�]-�SOS��!>H���R}�by����f�׽��H>d5����5}����T�Uηv�D>���|��(�\J3[���!�UWu��*uM�)���<t����Lʀ���$֊FK�x$A �(wG�l����,�T$R���e�QS]s��L@R+-���Hi�<�6�S��a"�.���!_�����9�`e`ji��u���N�Z?4�E1�Bz� �B�Ą朥$�S�-E��R_����1|�� /�jHDW�0eh����6�E����I�.i�V"t?���㘛����f$u��߅�{,�g*���63��|2��md*��_H;���U�\�b?�M��ds`�NIǏ������ۿuT��Y|):��l��)If�S{U?�*��g-)�>���>�8�j����p�fC�A1�!'���,OW.��\��
l/�9��/zL�m͑�w�=f�N�nC'5�x��ػ��㻋�㜸���w��؍w��x�}3ܽzk�Up`Ԍ��3���OP��a�qI�����S/*қp���rʏ)�\�����N�*�{�2���zb)x�|�07vL1����0���V�N��'��t�J�U�U���U���`����4����ON�q�21����v\�yT5c.j帎&/k��H8�u7�e��W�z�"�9�i�8J��.�9����#Υ%�����TX���'y��Ch"����o�)�@ǎ�?��Vn���1`J�&��u�o�H�!�pu�π�r.ə ��*��ҨU�`K���XNI
9ֱh���.qݮCu�ف�D����ܾ�jq�����J�Y��%�+��-�C��G>IZb-�Jl�kZu)���x�pl�?�s���t��睝��86%%�W�T�c6,�b)O@�3u����H)ţ�`�.������ޛ�ه􇏮v�{"���-��KU��V�b�3����2eX,��
Qo���d���n?Aq��fY�g��A�cRI�cp�/����6�����N��V�����L�d���|��{?��-i%���oB>�r\�Ι�m��:�3������X��q�>~�L3����f�w'��Q�3K��gC1s):�O[�z��R;�hQ�~��娹RY�N�/�ݫ�_�H?o�Q<��U�3� a9r��2�D�O/*�����
`�;�6\c��&ڙ�7�l,���f��b��Fh�n�%5�EM"�Z�]�����$��o̬{D|���.C����"�*�E��c���ch�����t��>
 �y���������|�$	�J�i>�+O�w(b��Z�
��y����/�|�O��)�Tw��uto��/9%���N#��@�
�A�MH(���V���K�*�0��`��Pl���ǟ�W����پ?4�]'�-6N����z�|*J�z�G\�'�&�줉BC+�k���å)x�!���|�lŷ�8s��k+���n� ���߄� �:3-�%JD�3F?r�Z�c�	�*�����@�B��J�&��5�M��<Lrg����8��p�_�d趩։���#�� |U�~l��� ����`h��ȗO����<�yM�lL�ə#E�<��-�m;sAx}��5��?rm~��$�m�w�J��w5�_.E7SN��V�(:�6�O���,�5.�-�r��:��w���r'�]�B}�y��l|��C����E�q�JUQ�T�)Ul��jAv&$��u�e+�bHU�V�J5d�と�؝�=\��l���4�͓V�|ê��%&�����3�`rsQxarNL��¢���o����z���[���G%��vw^���AC����(��H��_F:�J0�����; ��ȭ���k������N�xС����+qn-z��X�>m����r���Aȁj�Ö��~+��3MJT�Z��WSۄ	ٺuKA'�}��?p����գ�/i`��~v����͚��
���P�z�)��!�#S�`l���n�yS��Uъ�9�s�t�tMD�
P�ΰ��,�A�cLs��'1Ę��o�X7��5��SiQ�¤o��)�H�D�o��,(�-#W��!=#�ۤ�B��F��N�|\����ôLb���4��'}��4Թ]/�|$y$����u�gؔ�ae� �q�|#�Pؼ⭤N@��S\�l����J���	Hj�V��e������P����2 �߭tw����$��C�c>���9�2��S�
{d!����$�2�8|{,TGɑ]BJl��*�R�]p!/	@KoM��L�Kd�������<IRF���_?�P�n��[пv��k���uo-�z�lk�;;�Wޒm�a��M��j{�?V5�U��EN�*?(g�H'iF��q���YD�)S�P,e�2��|�����u�e\i���s^�2^�ê��-~�)���ε��1��HT��m�ݴ0�F�~����9���}�5��3;����+���(�t��y����_�OIJ�n��+|����T1���)�M~�1iTC��g✩��O0p�j��k8H���r��3悅�u�3q� ������a�Z<���I�Џ��`n�A%��M?�i��r�!X�'��qj��9)E�B�rb�9�Hnn��{�>(�ql]8���kHGL��C2���� �-��A���L���^s֛�q���\����m�;�tƙd���ߐ���G`����������
�,�r�3pb}�HjK���;a�c�sa�t�or(�����T�kq�Gh �(nc�0O[:��,���Ezi=���2�qJ��ӧ�l�Nzap�j�돎0�X� �D)�n73Ӡ7��4J�~[Sq�Shԓn�:%� v|H~5�s���e�{z��E�((;�_�ZmVfz�_!�I�Ѿ�3�8��^n�F�o�>I�9Di%r�p7T$����E'ز8�h�E������A�0�T�D�|���A!�/��A�O�R9:�nS�v���L{FTe�_3�92-���I��v�C��F��#��t����~��ޢb��}����wa�[�
��F���*U
q\��|�Rc6Ɛ#A�����+�겱�pG���6����,�y�jhޫѡ��!qX�f����Ԏ7ǒL����(̔!⭲Z3
�,֫��������;F�6u��cj�c�V�I�|z��E�Y��l��b�4ѐq�
wf�R�Kk;������
��C�a�{+�R<�~��?��Gy5�T���(�R�T'��D{(BdŶ�7��tم�RUu`98�"�f�ըљ�e�R�[������� V��G{"�"U��"R��Oq�	�ɶw��-���oVR!���i8!�ᦌ:�<�D�%NYl̴3��
��xٍ��4�����j�J��X�a���AZu������ŗ!`AF~�F����ޘc�C,n�s��6�L�����D�.e��$��2��:��]U�%u���%CՃ��=�䥣��m����	����]�ּ���C?��5��A�&�rH������m�.7:gOsSd�,!&1��b7��g��q� ���ڴ(n]� u�ç����ߜ	����҈�I�s�0 ��M��2	��>�~�%Yp�>�r2�nl�;���r�(*�.k�w�LUj_L��v[8�=jVRy�&����T;�3{��E��e�#�3z.��b�iK�����3�f�PP���9��{e��u�~�N|ea�*W��"������D�$�D=W#@�=U����}��+�Mr��D߹m����-[�r��P�෰b~(�{u[�\���z������
s��ɱ��=�`i�SA��Sb������'��[�ܠ�E��TH��9�jpS�@�C�2�Qm��X|��q,V���]�\�c'qi:К� 8��	�z���VnL�����'ez}ej*5��hP��t��o��W�,ɡ�3�sR����ñ������@�K(U��f@ҙ��1��'�˥J�(�ɳ�����ZGw��d��	q�ٸ�`^Gm��>X@����l�[X1�|c��!许����1���u)�Vi��2G^��)׭Q㿿E���r���R\t�5up¡M���m�nj�r�(S����`��U�s�Vpt�N�1����_팤�\����e��`!�Pp9\1q���R���(}��dQtgh2S��W���ocDW/��'�^�HN��=�_�g��`�x&�[N���)�ُ	����5�R��|~gFt�>a9��y@���J,���$�'��_SXz���@jqa�&��R����)����\.�w� C��W/~�e<��H����=
Z�O\���M���i�#��B�*iv�c�~��hUO�N��l}�7��2n��T�}�\�K�涢'`$r@�%������U�A�E欠Z�dN��� �8�Z���Y^��z9���b��__�74l>�������I��5��K/�t��sj!{��|1F���tԷ-W2�/��)u���He�>讹�Á˖~?_[[�s�t����居�sx���{��'��!o���k}:N�!L� �����l*s��D��n�X�3m�쇀&l��yR���P?R�̓E�ܐװ���d��� �����ֈ`��k�PIe��i5V��z�LfH۵Q<��q|J+7qԧ��;:7�܀���/�ʖ@���e�ro�oh�C����X�z���[��w@]#.�گ����N����H���_�������$��'H��G�Z>~E��N�7����J�.�MB*�EE��jbU���
1��ȳ����m�RR����qZ�}]���@5�O�TqC�Ѭ��@�75fIC-9�IJ��k��V���~?��񋛨��6�Ϩq��Nl|��Äԕ$��	�\~���q�MS�"(�X{�S
��r1��`���ɛ��c�hX/4>��c���N<���,F��rH��0uZp�3����5u�PU)p�q��"v`2���ܶZ���l�Zk���DzLr.�F��'ɪ'�vx!�u���(� �.�*j��O�}��@��z�P�N�����5�{h�Q�ņ�B�x=�uV�4-IJ�����u�F�4
�e�H���赪���pa���#�5624�y�x�9n���Ɠ��x;��w�J@�;��@��X�*�1��fx'5�|�`Г-���e|(GG�*
˕���l㖎�k��?z6\���ЫT��V9�
�.��.�\�و8�.̷WՒ�e�f��������D�1Ҩ�7\uAaU���|ɵ�<e��|�����vp���&�D�����r�*ܲ���*#�9���a �O�?:�.n "�#��}?T���EAF�$�v�����%�k��j��Q̱�ah~4��v<�e
�L�[��?I/2g���Q�+B9t&�^Q��яy�H2��F�lAӏc����(�I<���_qt�?߷�E�Ի>�g��� C�����C���u�398��E}��i�z���t[�(3�{�
�1�A2�
2�f�T��&��G���ӥI�{Z��
�v	�nI7�:=�b�l�}H.��~��"sV���^����|�>֏)R~2��ɖP�4N��U��c7�N�8Vb�S��r��O�v�,��j��p��b�ه�X�f&ڥ�qZ\1�|ڏ�]֦�9^|�ۖ���k{��!�|�_}�^�W�4 �;��n���f�LV�=$ҝ���JF�-�1�`>b��w�j)�܋�D��9=)ܩ�Uc����p�g��$H���a�r^'�(/
�<��c����>My2ś����/�[yj-���:��j\�ʆ=�tRw]DK'~���������a�/�ڂ�P��<Xu��"���,��N�q�������V$~��E1�$��g'M�LC^��[+�~!f&|Z�J���-��*���4_�]���l�g����5���K�k�
��k�q$X��ˏ��|�z_RZo��Ÿ�&�)�e��`�o�����%Q��I�����Lū0��Ŋ��q����D�����jY�2��~\�4��kp�L>�2+'	�-�_;���L,�֮�sG5�H��rk��[.��~�ET=H�,�����E����W��kA����f0:2����1i�����*@�����QZ���e�+��{��X�0ˀ��L�8��0�����g,{��p���S�:��Z�<��@إ�LJk��8Qͼl�i�'"�U���=cT��>VV����r��W��ƵI�0�Y��jA 8�l8�.�z�F�JG5�'�Р�[B^��N����1�!�@�|�X�VL/z�*�j&�cg���*�p�XL�1��(���҅�\���z�"���YjN`���j�kЋ�N��BO���'hV�T��DH��xb��^<��@�4;�j¬Ԭ ώ:/x�V�B�f��������sלH�8E���!�xGXu��ԃk���}���p���@���si҄TB݊�hCt2�]��$��3���%$��@`��)#�r(
]5���Yw�"�D��3#E��������p�����x|sA��S����_3��VP�n�.^#|�9�o��Q���+����L�������"��s�����ܩ�Hy{�6�FY�Í�9k�|AcN��7[�)T�/��f/hbnW =�������n+�5>�K9Q��,�w����W���!gqU�In��W���e������@��R�*�	T�{�h���� Z�����Lg�ܘL	Bz_�<"��WBy\����]7�G��H6D�Lǌ��9���`7b�Y��y4�aD����h¹ǒ5۵F�d��ke��<����Y�Qw�o<���������x� �J�k`���4�ժ��~^��z�MS�Q�&/Z�c��>��կ\��d��wƂ�G����y+�2"a����S�������z�t�+������g��m;��{�\�2����2�u�~&��G(ըu�n��.B֢�ކ���v�w��1<
�+$de�Y���W��r�'��x��
(7w�O��l��F�45��PW�f.t��2��+ �#����T�<b^��(*go2�0L��.��;�l��a8N{�=Ո�+n�_����Fi�e�fL�푐_�/d/
7�K16�-Y�K
Mر?S!�������`�s��������f�v�Y6"�h%@TOͺjL�/et�h��Ԇz��r��[ ��J-���˻�li���j����A�ʖ��y[�R~{��p=�g��k���>�":��.��J�ǎ�B	L�a���!�/TG
��P�l�dV������5�#@c6����މ&'������3��G�{(|�$#�Ll��{nM�GZv 0�|eC������d�1���"��$�3�rR����Y��"z
д �@'6�/HK�r{�������N���#v�Ur�pB}�� �x�(V� P-�ŉQ�Ct��,H�/7	Q*���AӒ�;��h[3拏������wmN�厝|�|��O�w�Oʽ񬗤*vN �Kr�յ��R'���2��t0�[��ut;�@��I/�+���{�wn�zu�ݣ!4!a�ʷ��b����5��;A����!�1�	�Ӭ䟯�fˊ@�Y�@uN�wH���م'�-d��x|��@�I"+���kݤԭ�:#��ñ�C�\������ ����:�X���~B�sbO����D�`�l[&���ڎ�i/�Cn����A��7���`���ͷ�7��fUc[I��*��@4���	��iq�!�u@�S VjZ��7i	Q:p�R��Z�c�$(���|^%��Ay����:���տ]���a�" ӗT#��db4v%��X?���s�$��q�e�8��L�/=Ժ�7d���m�D��E��"��zp2�}>��a�+�-Ls+���{�,J����ע�邾���B�bS `��y(�ҷ|��;�/0!ɟI���޵I鲳WЗ��<���?�n����.R��=�4:�?�@����ny� �H�aժ�H�<�=�r��}�8uh	As�L����)U��F�Ֆ����F���1������a&(�Q\�t?c44�	I���_�\�~S���i{�9�J����U��01X �!Zю���G�-�R6�2��d�Xg��==�[,��f i���o��
l�w8�d�O����L?��V�6�y��1(e��`�8;��d)#7����ԉ+�|�@��W,�&�? ܫr��ʚv��r�C�[����7y{+�'%��v8�����6ì�@ڳ��b�Z'{�Ga�\��eHV�"������,'`^NVREy�i�f��s�O����S	v�q�?�'������?�tm�I<�=^w��#�r�VT(u.p��Ձ�~������T�`
;����T�=�"�1K���A�E���|�����L;���zg(!�zSK �*F�Fh����ܗ���2bנ�'��>���l^���|d�����s=g�2�Y-<P8M�,@����!.$s����j�t#E��50�Bh���ز��t�(�X��\`U�:o?R�w[��,�e!�&>+n/h!�S��MSL�_�)��{$�䟻�KF�����8���ѪV��|ReR~�)?.֬���eҬ8�P��̀���O[�0C7�o��1������p��3}�(�����uū~=�6��8	*q'DC�,�w�4!/u�ư��}�3���<>�h��za��e� ��&9�ϭ��/%=�Ov͐�1���k�DM���'��r'�izf�2X2����5�%���kW��<$@mf�� "���!ЫtI0hQc.�$G`�/x���N�/�/���yu^&�W�cn� �3�rw�ղ����Ň��e竢�W"x�do "j+����VbVcQ��� Ȇ���.���*�ܸ�TtB6)|�2Ӄ
{�Q�c��O6*�G>j�A�����&���]��U��LH�'v��h�>���9[	�����1C��nz����B��h�� Q=��.���j	��ׯ���?�+����P�Vz�0J�ހ} Y��rF�l�W����fRҮi1��ݎWS�Q�ͤ���8���׾gi���P��}/3�x�ȝX���_)����t�,�b�b�Q��%��*U[��X���8:;4`|D|a�z�d��e+�x�"����{�ٽ��y��3Y�����36=	�o���w
�W>�Q����lk�tW�P��7l����3��M��G�k��x���Xr�����oq��HiwG��2����f ߈o�e�}[L9�U!�`JP��Cfu�X#�d58ހ~��a&��4�LaW���P��ƺG�����q�J�X�5e`�[_�6`�������h����o<<���!<en(�K#��!�$r�J��Pi%xp�;��yK~d�F���9�KM�%{��lrg�wC�x䩧R���n˪�P��f}]�%��&�CD��G #���y�8w�:,�Spc;�~�w��/Lw�	(��D&�gXρ!���ŊS9K��b� �|!Zc'�/\��v�~��cM��٣���bY@"������Rz�6� ����}��8�"IU����څ<\�_\��!�W���$�?rxG�Yj�w8� f���̮;�j&��T7�R�Q�חTpL�>��㓝�	�X.�وʔӔq�s4��Z�V2iK� --�78X�s�:P�藪�e V˲����1�^�Q���d�����ͭ���`�kJ<(Ў�g����R��P���k���B�
�7�l������b�T��u�E��r����ŵ��
����F�4���P;
ݪ|�?"A���Q�Bo�:�i*[F��U��4_M���٠-��m����[���g�_h�¦a�P���+e�c������Y�C��B�-pO�� 1�[0ɴЦ�N���� p�rd��bݚ(����{�O!��p��XR|���G�Xڙ����c�}�ѳF&F���&�(L�yt�G�W��	�Y�yp2�/��N��,���'1:��=�uгpT@��#���L���CLE�ݷ<�j�}��nTy1.ʺ-���]?�v��)>m�r?�T������>�?cS�'Ov�>R2�-�������S|r<J�����fe�ݻ�L��%@fFSΏQ�;�����.�l�e�{z���xjV��x
�k�Z3-�"�Wt�Q�]�s��-[�!	09�T[7q���ڦ�xw���Xm�U݈���ﭗ�I��F�= n��o�Ȁ^�z)r�p^qg2+�������?��� �YE���B�aN`� ���.A�5����%�\��i��k�|�T�8��Y�g�!���=�}u���l���C�_�L��{'���q (׆զ��r:G��N>�H:�hE؈`֛�40�׻a ��#_�\������D@��L�	��_٬j���d/��t�+N`rpt�����AG��Ȇu{d�0���O��}o�k+�]�ؙ�.V�[4q`���4p��Br��m��9~� k�_�ՂY^��ٳ��Vx�ӄ*i�sWw:��#F5!/�X\�{�r�*# �^3�y�U**�Q�"0c����3zQo]�;����F
��l7?:�Ҋ�a�)����X�@&�: r�N߿��j^[�5�`�|��.��z|Z���i+�BD���⛪�$��v>�g='0G�5�/s�m�	�l�8��Y޴,�T��!<��ت�WO-�Q�6E����"ٖ�Я�x6��V�������/]�I�P��Y���o��=��������qq�����o�uu�|��HYNS_
�G���3ds��h�t���F>�����z�y����� K'��/�pS�B��@������;�o5�P�Q���_��E�o=��d>��,��	O` �囪$}B�;V4R���T�=�M?A)N���y�F���剦�iy�V��f�[j����v��A���+�q�DM�1i�6���8 (`�8�)�ܑ�	6���:���C�.��j����f���h~��-J��' �#.%�f���F|u
Ջ��n�գ��Jc ��Ā	H����z�]hO�yҾMI'NG�ݣ\�)���u�����~��.3Fs�D��Q'-T�y�'�T�����*�R4e�����H�V��4�hA�~��VCN��k��$��hM.9)$�7���#�*��|7���&��y}��+2e �eV���#�{n�bN0���j\ߑ�.�?�R(1�نa�.û��Ibl�.��:��9�2�x� ��;�5} Hr�쌎�
�D�V��n:Uu	ڸ�pU�$�����/���S�8��!��0y�����<y�3�6���a��*��eW�{VT�+�kt|+�wLǱI��2����*���,�)�q��a��H|J��ȥq����{�8�+�l���3��T�:.�;�Kɏ4��~�\�˧ڝH�Ն074����q��ڪ�F�Z�%��u�� �KC'#�'�ivK�I$�rSi��k��Gl,1��k�@}9�$��x���Z"�m�ȃ���^��嚷D�&7_���ܔ�MB�m'R)�M��޾S���0�&�X�NŊ��>�+l��fH�Κb�,�Su�4�d�Ҥ�k��u=�"2{�v�E�6Yx!�K��!�.�����g�ʴWW]3�i�"Lll�D#V>�M�_�ٙ�͏�ݥ|7���'[��Ax��M���Q��� �5�"[n�[D)y��h��3�ԏ!�L�
z��'��������d_F�x��	P��av��a `�,���d_�/,n��d��3ld�C�F��pǐ�Q��K�'�}���9�/�;ɇ��ږ|e��t�寭lb��E/��T��!�o�^�y�ҖK,��z�/�v>�m?�&*�N[����}�AVR�����#b�����A��J�>P�6
��U�p��N꘤-	C����Sx9to���1^3��,^��*��4#x<�Ǉ���G�hg�-��:�e����|<E��3��li������"os<ÀݳOjD��sw�q���)vj$m!��l���I������xQ���o���TVB�~\�� B@��D�?h6u��
��G�~����҃i���r𽈡]��+������%�۳�uU4y�d�����\:V)k���%��W��G�$��ϖ��b�~���/P�;Wҕ cη!tHL�1QWU�Ч���:[���������:�6��!Ca~sR� ����~ct�Ǭ�H}��z┋,50�����,a�d�o�� 3�>MY���u���'�M�����(L �U�_ǭ	ul9�T����ԕ ���U
���2�IZ��>�Z��v$� �~�u�ls�H���|�:�osՠ��.]n���(��<PB��H��5 �$��o����������l��	L���X���dp�2������6�6;o_��ߟ��w��/�X��꾓ؿ^&&4H����pA�a��8ù>L�y�>�v1$�Hr�fI$%��=�/٧�Bvk �#c�A1���, ���4mz<ǷY�����p��f!G�6���S���ek�ߢ0iP?�G֦2��	►��a��_��=
��2�xK.��&��-8a0ߜk;��26u��W�M~�v��{u}���)����9����l���0��v�S�
�SxZ~W�����ꦿ[s�^g���Y>�V6�`E4�-�z�P%���S��[&�4��}�n��u�;3Ԟ��ʖw
�g���5�go3[�?^/����V~�TG�O;��)�Q�!���hk����i�̃�[���u����²X6���
O�Hj��5?�e�\���jrzBj��������B�`T'9��g�7B~+��O��x$���C��1�ӭf'd~���#E-�5���������ᤝ��[�6r��Q�&��	aR�n��\�ʼ"ꘒ���kN�����}�xZL�S���w�)��z
u����+�ٗQ�P�jk�_��N�I�̈́���|���''���9'�$�y��'�M6B:�I0c���a�nQ��qp-牖zsf�2�+~�G�4W`��霎 �&�ds��;x5�h���m�F"SZ�)x��|�Q	��-����VG�c�>�qҀ0}Ր�Ǒ�@[��v��G�����R�`
�~��B"D�����(-��~��H�;��$�5�U���\���W&��g�	V��S�q�ň(4��������(�4ݳ����f�>��@t�m��{�O����k��H�e.�Cy����+�ͫ+�V�ؐ��,lD��e�8��ğ�Y��!�-}^����7�ydr��f	�����ݦ��AB_��E��!�)��!�7�.�{�jw�)�G���0���~����f+�q��ɓ#�,��1���?5̸�ztG�;t� 6��K� %����k��f�5�,��AL�E�E0��*���x��Z���Qȋ��p���^�H���O���mX%;IX�P�7L�~�7HQ�^m�h��m���r�C�e�Bj/-ҽ��� )O1��g�˰x�Cۂ�Ӯ�Q����#> ��
i���l~�����b]���Ò0���pBD�P!,�:�
�݈���5;����x�M��_��*���=<J�y�L��� t��6i��K��d�*v�:�
�!�����ȁ-�&.�P�T�FJ����=���B
�����u0�5[M�?���M��g蠛.Ӎ1�F���X��B&z]?V|]��h�����AY��"��������z�O���[P��»Pۭ��J�nnR�f���ί�6
��������T����"I�C�r��������b�v8����Y��4���f|V7�/��8�5��N�P�ZU�2�JbX�z��E�E��4K��"�O�L�N%p~|�OI���h�pe�e\����o܌���W ���V����7L���Ѿl��ǏPζ�fŇrW(�k�]���Sl�ua����q0MSɪ��1�Nf,�g�8����t�c���Sޘ����ޏlD��D�1X�L+�� ���2���;Ҧ|���S}���fm�Y��3?�(����̞�oy?T�V�ǚ0zA�E�!�0�-&��|�v�'ZVc}J��Ȫ�M�
��V�A�d���#�������k���/؂��Q�"�̱��`M��m�"&Ers�%*��P(W�K`��x�:��*��nq��,�M�:d�:����Ê�o{O��0B��"ϳ��Qַ:�
\5� ��:�Կ����)G���"�Hх�= ���.8���l�0���'7-�3�h����)���f���1ni��wE�~���.������ *h���R7�F�<�8�V5T�&�Z����:�b�o�k����S8G�5��y N�9 ���pu�>ҋ�k�Eݶ,����ym�A^��͊,��d������0���b�Y$usB�'�a,V��iNH	���W���������l���^��Y57���쌪|����yi�vÅ����m l;#
#�z�yА���ә8����F��.�jĘܩ�TF~�CvNs�Q�zCR荫���W"�d���DHG�gb�,��^�NU��U�v�Cd8*��I�J�8U����WVP-�K�j�r��N�ν�"+�A�Ui�=�$0��G��H���F]x~�K 2�'2���t3H�PYh��[�ϯ:GƟ�v/E�l�_�V?և,Ӡ�E�Թ�gݔ�Q��-E�R<�,�����C�E������8SGFd���\�$;�A��,���F�D����Jk��	�����[X������
F�~i���~��0%�F{I��E:8�[���@R���i�W�z Ձ
t�|xXJ�J�@���)k�-�8�2��g9D2F�Kk��V�P0��m�,\���R�@Q̩؇�.���Kиy[�Š�֝���M^�M2����cw�0�0~����o��{"i*�|G/���L��׫@c҇�Rdma�n�#�.�)���X�(`�0��粏����^3�c����z�R��� �T�L�jU�r����2s�>� i��:�w�X;�u��n	��!=�V����f�x�*a2���oέJ�&�?�R�����e�	�i�a[�ܪE���s`��¥��+�m�5� u�8G���#B2���jc7"����AU�OY;e��=���	��g�$s]�]?�n�o�������*Ӱ��
Ѫ'R�3�	����E�o?�<���Ρ�'BA�D'uh�v��T���&=�|�v!P�Х�]n]Y�����Ts�R����=1���|��,2��8% ��@�w>����c|��dV��f��}��xb�������z��n\kZ�&�5�n!	�0���̝n��ؔ�@ �-��{Ы�p9���.���0b�y�,�P>�b����d!�}����rE���ظk|�*��d>1ldg�'���+�MgE�}�Q�q����%Wl�1
H�5�U^�����MN�������FG��MMI�~�8Oq�8n�xW�����x���]馤�CU���a�<v�>���R��|���L��N��/�#�t
~��N����E1~x�ˍ$|�$��Q��}ϣ�0�5��C�Y�
�#�^~�����k%�n���y.�]�bL��%+�4���ͣ���r�Jn�M�/g$h���>DJ��''���nr��O�y7a�J��1��F������ �A���|o�b�;IJ�>R%�ܨ�9 �h�:B�#ϸ��&�:���o��(���x��R��xj��n��*lt���$ #�6� ��Ǳ�v�a��,#�]��FV�~嚘��%�vj@{��fo��菧��~C�N���kۏ���'���~W�B�Nʭ�*K��
Z�
�/cg�v�T?��v�����F{�C>��`&᳇���#��
LP�s6�,,����}�S��n�2�y�f�>�T�Q�t�:&ǒ����VN!�W�<�xjq9\:���諊�/6ĕ-�٣�t!��R��V�f!����)�3�1K�S������p����W�0w۔=^�k�"�3K��$o�plk�o�rekd�+%�?�+/�ES�h�Ǻ�C�r��ě��Q3����C�G@CD���.΂���Oe����+��JG���ϙV��eQ/��v��n�K��չ�.<�=*��p/^�I�سG�'A�o%���1��+HF�[|�Lx�|�]#8�I�y~V7��*LcƜ�3��Qѻ|��_q��P��:������+�6k�7M��ef�6��°�B�UA�UI'�~��'�*Z�J hU|4��z���$�Kx���_���L��ך�N��D��������d,6�HHp�f�&��L�� 9[��TI��i��p~hh\��dRZ����D���z7%j�Ot6Lw I��sS��&��<��ƚ���U�@sn��Ʌ��Q��|��AF+�������UVڂ����H����Ś�Z�{:FE*s�pwI������[���a\n���AZ�����$X\%�"WtlLz_ >k{>'�͆��\��hW���4�8.��p����23�!�-/[�P�@"Vq�X�6D�a���óG���B��"\ԏ�~��5~U/�_�V\5�M��\�Iw�Rf0{�{zg�!��ˮ��6ީ�-}��)��z�:~�{�1G�|`�~��Ȭ�?j����XKp=�~�Gfa�)z�V�fq�
='�;��me�,�.����O��/U��L��d�c&��s^���y%}&Y�/����R�-2UU%�ߓ�M!�~�RCyc�֣�I@rH	��y��(�ې"�a��T�d��'�i�-��\��4����ec?Q;7��2������.��"�ɀ3橀Y'ex�\��媙���G��0����kiAG�︑L�NwB����G���$�54MO���骿Bbn'������I��谓Q��r!�G;Pśd��0��4����}�y��5������-�B�F���e���@�@�9����#�ZP��nkk�A�Ð`�wzLR�H�74^)�o=:{��iRL��r.N�L��ĕ�Ϗ��D�̶����G˨�Q�R��Z���.N��d{���O�K!Z����e�VK��@sZ.e8Ӓ��$2z�v�tG�6}a��&ӊl�PH������#(z��D�P�X)
ԫv'��f��R����Z���?�$��_��k���-L�P>7g�"֔.N���[�����E�l�-[i4�uq��_��+b
j)iKC�?�������Q��E�hF��=F�8~������l�-�{�Wy�I�������i��X����W��!�L�DѡY�χ�`����5�_M���0�&>f�eJ05��	�f����l���>��'�P�v�MA���nPg��h��|?�-��TaX���3'���<k����V�X'��E�Z�35d�d�o��� B�T���}S��ٱ)�:#�}�]�A���¤{}�u�����ie#i4y�ȝ7d��B�����A�~�#�aG{\�GV��s�\���*T���8����R�<�����:k#:�持8x�'�3������Px�p�{������z��+J$��tg��e�u�+|��G�f�}ns=�p�?�w���sڈb�6�HE�1y��Qw~Ѵ�o�����H� ��.'�����oY�E�l;�~]7���i�~~���em�o9K��s�6�;�)�x�9"q��OT�8"�9�ݧ5�bgU�������~���vۅ���`���aG��Y#FB����Đ��-��v��ڣ�����4*n/��Q�l�s�Z=�c�b�5I�P�+ �:���(w��n�G�Ó�q夃�g4Pc�j�w��w3z�H>Q��_q���2q�+V}|G�;�@R�"�~W�p�s/<��^א��J�V�/X=cSr4�~�% �f�Yt���zr���K��E9� A�1G��� 欼i�VY}�ÖI_������/zf�W�@���)�����s�;�UJ���l)7�3g~�pۛEli��\2�9P�7�ν��T�bOWgPEIi
:��P�9�Y�.�>���?r�5���O]3n\=���R�W�5�����iΜ ��a�bY����Vb8���f�r�� ��v��d%ü�d�P@^D)�%v����.��&�0�_�(<���U�=����b--��zqJ�z��T�����BFv(�,e鐵��O5e��20�%�p A}`?��+��;$��X#�k��O)�3q��k��EW�̺��&>+�'$~��j�G�*9/�0���n)Q|�/�f����r�U�WSz4��7����re��'[h�ؽ�$��\	꡼�RZyzr����z���7Z�b�I/6f6����3sä���G  *]���X)X� �1́�;w�~����-1����_�^�!�<Rr�ޱ�V�)w�0kk���*a�*\n����<�g��{��P�r���,T��a}ǿ�G_����\G/:���3݋�6<����㶪�GC��7�?� �#��V��\O��]{bU�Wʯ&t���Őck��@��^�5ۘsOy��[r����(#_p�����u��eK]�f��ynZ���/Ĳ�؍��B��=�I-��'-E!Z�K���½y��!A��&���B�i��?2#�Z��ʲVy#4<!��A��6�j��Z�W�A��X������]}A�GlK�q�nv������7w���6h�FUgźH���ɦ��W�C�>�rO�й|@?�+���=����9��	T��.��UQ��`�-�Y� n�5e�H�9PH�@"˥����g>{(+�!'TǠ�&��-"�}!���O-�Vj�j�b�t4=��.�Իkkb����L�_�����c�;��k9,���T�h �cNR����+M��NX�\b���-�kޮɏi}��" ����	w����<���4�+�"�ê5�>H���<;�m��dS����7�uʊ`����#��ȑ}���_Hm����6ʍ͉kc$�y,�' ����e�|��F�=#�id�R"x�/L����zЋ��I-�XU1���5�%n�*"��ш�S�i?a����s���Jv��@��0�L�xj�!��������ݬ$�$�[zU�𠾢6��e�s3�D�(�W�kTH�ѥ(�TĘ9�v�I�P.���i���U�8Ǳ�����Ԯ�ץc����`k�f)��(��~���}F�Qב{����+BG\>mb����i�L��/z�R✬�AO#�(�\޼�S�s��2?��#�]��=N�����5.5�[lyW�`�������M��Edi�$�K��wg͉7$n�|�\g_��T���k]Z4�C`�s@��|��fOS�M�3 (�p6�i��n��>0!Ea6ʁ ͌��^��d���[E���9�,�����Hh�揞���������C&�s�莔��>	����1*ԞT݇��%u�Ey�׽"��?�L� hޭl|�+�W�U�1�3��!���r� &��� }2o@un"�N�|�q����Z���%%~�+�$�H DOi�)�W^`j��rh�(M���I����2���ҹ8 ��x�L�.qA��6�B����&����)q]���.���w	Ź���q5�����1�g�h,���{�<�*IIl���T�����e��b ��T2	Z�s{Eam���8m.�>���E@b������	)i��ê��i`��U��Y��m�@t��6=۱Pxݧ8P���;)RL�<��?�����P��M�����_��r</�{�۝�_��(��ףI�Ϋ��KD�^��J7-�:�
xc�ǻ�@��J]͊^˻i��Y(ѯ��.�:pN��r&I���+[b�ie�qO��_߷�mGA"� 
��T�?hd[�8;��d�I��U]*�{��9�Q���JL��#�a"
J#Y_�Es�S�e�E�*�y`���R�r�����P!����C�9p�?~��ˍ���Ll#x�HL2��J�uޥ��L��1��0�~yO���]7=j�pݐ�~.��h1�p�W�wl�U�͖1Zyoo{^�1����豬s�@ ?(k����k�s=�gh�# �b5�k��;�ť�[cV}�y�@A��qI�?�C.l��)xr�������5�ӫ�n�d�7�&C�����.�>g�FS�D�����r�DJ'_�<\�h�xT�U}W���-�E'�	��3$?�h�NP�p���΄D #1a>M'R�p�*���? �u;V"�Α���q�ƠO�|ݸ�7�Os"����Σ�6n���¡���,]�-�{BSb���� _R�|2��*����<���4�� [���7��C�#�ҿb�(5�EE�������4e�>�.�Ϩв��?r2�p��^��;�4��L_�ƛFy����|��NOATj�/q�N��ޤ��
v5&݀o�w�'� @~LJ�t�����(\u�q��9���3�ج��_��֑G�ũ^��c�l���^5X�4zB0%���{�1�O��h�V�����aY�}$��x����Ja)b!wQ��`���L��W(� ����,�&�apk��~Q�(X�.e��3��=��A�V���2��ixޚM�_x_m.�0� 7@�� ����k��`w`;ӌ+�k<3=�"e-�o,�u6�<�H`j����\�_�m%6�|9����r�Sq��S)���� ���S����0O�p����g��đ��!�;<�ޕ<�|���@��}|慹��\�d��U�o'��[�f.�
���[B��F�+���䃼P�n��=��� b�i��*q��*e�����2L� ��M+��l19f�"MFt3��<����t�[�-��A'���sLn"��{-��A���jҠ��NbU�|k!U�r\,N���~M�nZ��t�5O�֞����D�]d��TF� 1v3�9���;J>�`q����u�*qe��.sǳ��1��U�>9��f-膞0��	ǤX3����D��F,ߞ�f��"���(������B�(}�A�Hk�.�R�"PN�A�3@�.'����N/�?��hgjw��d%Soץ8G�dX<<T��K���YVFbر�Y'v�<��9K�}p�l�2�X���ɢ0�_���,�u[@~���a��P�@wۧE�?W�rՒE�$ͩፕ���G����
��,�kׯ�S.ԛ�߈�:44����'O���$��4�Vd4稸�u��'?��T������T�_�d ���&��� 0>���"@�ǔk5�w!`��ڪ���U֌75@����-!���~�y}C��f� :s�-[Ua.���ؘD�[�฽�RpB<��J^��Z����@��3xu�?۬����a��x�v�êP� ��""}<�e��`�Fy�]g=[��yl��<a��67�8ɟ���,g��1	bV#L<@-�&��<��jpy+f
�:���)���<d��O'�R>���+�Р�-�� u�O�Z��WZ{8��������n�J*��B)��뷌$�ķeS�ܜ���V�U�FX� (2��>\�� 8�9�=�����"1;3��� ����0kX�=E'��=��fgX��|x̱{��%!8]h<��t%�"
�M�b��0����]�����Qn�{�,M㉭�-�q���wK��'?��Y!}�57m�e,{�.�]��D6��m�2r���� �#��M�e#tx�A�PM�@��x����ܯ��𨖎�`����Q*_�g�R�gN�ڪEa���g~����#�i�Ye�,�#t{�7ξ:�����~���ٷ-�d6��H���O)V�2*��0*j��y�z3�u�j����a�4�
�d�MK�h��,l��x�HOTA� C�m��Ouo�,Ô?�@�N%��*�U3�ڙo�魞����۞�4}F?�Ez���8���V��n�mBD`�8Nox�.TE�\��|��4,���u�3�%��*��l+UЭ��߯��<�9�@� ��j��\̊�zTrh���C���a�D���z04);�  {��'�!�"������ᅏ�Jز�">���3��`�.��}׭O%ҍ	 ��z� �dS���r����oX�]{]���ךn�՟�� ^|�{�����P�7�1>����H���O����j���>�o�[/�i΋�ᘆ}L�ى�d֢�b]��$2���s��FH�dx�5�!�U����#x���e���'B�P̉%d��R���~��rN�F��2���ѣ[,��mB��gK)�����	��K�A��bU/o� <�&:��-��Z}tz.(�Vf\�2�ަ��W�C^�8y��x˸��17�ƅg�0;�k����6��Q��,w�}��w~�,����;�Z ����R�CK��ɚ��q�j��,,Jd�Ce�D��Hd��.=���~Y���*��Ɏb5��[tȦUǻ����TK�,jSƩ�4L��T��l|JA��{b�wԷ%#ݐPA�_�.�SA�\�l2��9='���4�N���щ<?���p������`�3��tBW��j-�l�b{_j�l�!�����$�<�	(��TZ�퍙v�A\33��+��8p^��=��	XI�2�����Kٝn��\:�(����J���kkk4 ���#D�[�QY־�o��dLri1"�����°�A�q^D��,V|�e^�9S}��?~?�ޔ��3���0y3��vb:�f%��S�G� E?V��u�7 �e���0�N�r���}�uzvp;�d�f�~!`�J#`a�\'V�w�����L�5�Z�xQ��*�0�<���*���yG=�bC�`��l�<l�!�4
,�̠�_�2�o�葞 ����WY��󛡛8��n�En�̄+4H)Fe�?��<�xnU�A��l�* y�Wt%��Oݪ ��Hf7��*��mF�[����C�P�C�r��k��af��A3#Z�k���l��7������%��|F׿Q�wLR�ף�Ў7)����T�֩�o��mׄ��ק8��toջu�W���������J����UAۅ߫��k��;A�����73��x4�ɪ$�'�	�f����\Zv+�8O�|>���0i�9e+��w&�2�{�@�:\Q^�W�[Z���٧)�t���f���Խ�4%1nK��?V�5)پ��U*������Dq��>ɲȟW���~4�6�l�"����Uj��3�LJQ1�ƙ
μj���jЂl4�8Zr��:��*)}+�����͙��Y�-�oOe��r�������̢^	���WBƠ�Qb���S����K��T�{5��-�6�-G)���� c�8t*�󌠥 ^� 1�5.�
����";}����)�7��x��Ҏ�p�c�Q�fW�.Cլ�i��$s�Q&�ˊ����E���-�!�"��̔��n	[bN-M�O� wXZ6>-�e.�wB�֤�.1�x����Lv?x�xr�&e2����Hg����6�k;5]�wD�D��.�S�(VI6��7�D���b6�j���An�Ȣ�>Ί��h��8AE�L� �����$�X	 ����/@�!��^����ۧ��i���~����v����w�ޫ�Z�u��tį������D��3��x�9����ׇ�t�sF�;�LF�f<��F���'kh�E�\�VY,�����
VX�c&���Ch�w�Nc5E�罹�E� t�l�T�����R�1���t���ı�~���?8����Jg��`��	7ْM^r�J�V|��DQ���G/���@�z�� n"�\/�w�~G��u:V�h���/��2��ey4��yjݑ�2!�}{�<P�s���DHg�<&��n�6=d=��9���bja��<�;�I	�W �0�v��ܮ�'������z��n�ZC(�Y���չ�Hc�����:U�[7�*����@h��8����v��4j��19��C)�%ʝ}���؅1qɪ�/�[��$�:h��n�6Ad��ܚ���w
?�c��t��8"Z��'���ҩ.����2x<�X~�d�����
N.��]���a
��u�#�]G�r��1h�OhD"Iy���~`�N�7h�/"���H�z���Y���zڰ�`�`J�=1�Ћۀ�l!y�>+�aQu#�@疮�?�!�xUR��5�!�)��&���_�Y�J���T)�:�?b!�����t�>pgg�#㑧�=��2m+h��a�n�2����Xqo��-�F�&�	���4�n�U{Ea$beQh@���3���5�NQ�i4��m����>�@�ܰ�x��}p~�p�v����.#���?m�����E�T�m���Ĥ�R[�*I���8�>�R�j���&��ulO���ҍ�`!e�F���#�n~o�c髿Ô�B��{��sQF w���T�>�*_ˀ� ��P%��5��BB�t�b';��ۀ��O�q9�������;���%�u-M�ì�X�(�U����wKb�����3�z���t��	+��M8�Z��پ6��3�⋠��0�_����=DrhV������[�����ط}�:��A��}�u��ӑ��dB��	��WFc�^�kݩ%�y~�(�d�r�ƽ
5Y��XV��#�u��DhGE�|<;�*�bۢ��D<��6��h#B��'�� � a(��ua�t�[y��q����U�z�+��Bh�9]�m�g4/E⧫�dN��I�h�*3����:d����R���ʃ��@E���ʰ�e��F��g��[*)
?%�,�_���k�t�w�-n�AF���SDU��lH��������i�r���Y�WIT��[��i�o�5�lD�37�L��58�יU��I�Z=��y�'v���{FD���z�ϱ����7~��V+`5��\7 9F�۔�/m�KBr�C�bۃX�+�3۷�Λ�F�y�~=b3Y!O��F"�<�wL��x�*���@��t����"n:� ��~��\ޯ���`��Ui�{��?g~L����:����X����`b�7�
"�(M�UdѪ��R�B�p"A�e��	2����7�o�i:�/�&c��$_��Y���-ݓ�H��Js/���嵲��Q�¥�X3��~T6��C,�ƹ=(`�[+�������ڿ�k��J ��KJ�h�ݨ��e��{E���U�.ɹM���=p	�q�|̷����F�W���4B�j�g��o�T�U��g�K8u'�@�,F��Ve̔�΂b��Ӈd����Ȱl�m�He����w[�6�J�Ԧ�Sb
E-i����e��QN���:U�X�!l'mN�k�>������}�v��r�}�UW�gvTV:!J�vŐ3��Z�=,�3�N�w�NH�,!�D��;�5�5Z�i� �;���L����?6�b� ����3�0����r��^_�C��^i2�F ?뗑0-
]}�q��Jl�쪧��;�xD���v��n�t f��9��L^DR��u!i���wĎVʻ�����_F`�D"]1L��W�(�o�U��
�������6��7��5�6Z�f���{��j �4�Y�F���z��A�^|{mâf苩D��Rח�"V����o�U�3�_O�;=�&a�?�v{r��@�b��:�N��+}��4�U��k��\��4+��["�c����e��(s仼@$Z5s�u�"���p�����Ӑ���Z�,�uݷ#UT���	�6.n�m��-��3����g�%�hd�|k
#nwJd��]���ÝǢk�A��-�Hb��:��3��j������ҥ��lE�ne�{���,2�?�},���6HO�V~��O"d[ /n��9O�u��VB��]$��D�B����G`�_S�rlڛ�s��f���,Y�o�%%� i-�7��4��q%��<L.]x^��I����4�*֟�Je����1w�p�	K����?�n�o��{Op����Z!�W�}�aH*�Hp=n+Va��(	���x#�����5`O�r9�_���U-f"v�B�k�|���ʖW���}��^� �`�[�����K����q��F
���;��i���?�6HdX�'> yA)Z��	�Q�� 	K�:C�`�(���P=a�^��=O�����r�E��_}RĆ��΀� 2\��@��s*O��,f�:�	�?
�+�S���٩q�l1�jS@{�'�+�cB? �����ٮ�N۹=~b�Yy�u�=&�/1��/Wa.�����Ā&r^+�;n̼`��@6Kys���l��Z�����e���\�0����6��8�k�p� ow��#�W��j�(���DZ#�����Y-x��~����`Тܩ��	�����A/s�y�My�[:��F��^:B�8I��<�yo��$P�;��uk`�l>����5��oM$���_�ܬVCĉ�W9͠�9�آ�p!UȘ I �O+�N%ߎ�Rӣ|���Fb��ځR����笉3b�7-�v�v�~����B�����k\$l�B:������.���B,�_��n��`����@�$'�� T̅v��(}2��0���#��$��@�J�&$�볜GEn�T�nn叡�F�D�����Zޛ�\���d9A��J��9��G����Վ��(�^�:�5��O�i?��>� @喀`G�q�L�͂��`}��=�N��Ҭ
��a�sL*^��k��'W��G��J����f	49�i8�"��c��N�k��Uߙ]e(��3p+�v�s�e��1��6-��Gf���'9������]!�l���-*���RD>� w(IT������V%4�Tճ���w�4�z4I"9K((�+~����hߧ��"p�;���(��������9�TB�
��-�c���RG������yI�}A*O�����iQ?���n��@J��Qh��*d�1Eՙ��H�����2�Z �lG'f���v.H�g]<e�Ǭ�y�%u!KP	 !�a������Ba{�HOƜ�e{}z�\���3�WB$o�V,���՝-F���>��a�Xq�	���~�ah4�g��:44��0>p�+	G�K���Z��a�xz:��me��ы���T"tKNƔ�ϒϠ�,�*��^��|��
�_빠"%���e,��]賰0-�����-���ʹ����^w���=���$6?��&�q�rIAF47�_�H�~q�>s���F�����^���8�S��l�ν���rjA�ˋ�Y���ái��r��
�x͈��}��]u7��bjw>�݈�a��jOYy�j�߭$S���Q�V��~��b���Z��*����u��Tv�$�d�A�ڟ�v�Mr��-WC/�_&iD�L�0�z���o��G%_Z{�
┖����,��~�+g78zv�BGc�"|Q����)�#�����s��q��A�r�e�2Fʍ�4�!%I��I�o]��W��С?�C�B�y��)��3�UA+aŰ��`t�n���<��>�f�<ô�j`�4(M�vS�/�W�$BW��|������<����`C�
��b4��H�_`�ȱ �|D�C�~�nd��. QV�eGB�%F*7��$>m��x�_2��;��ܨ��Z��z�<o"�O~�I	'6��=�8��:�?ֹ�Ztpҕ��T�/^
%�Y�	�F�S,��x��"��nc��5�lL���Ĝ�f	/�R����x�Ú=����_K�@ �Zq����E�Yw�l'��ky��R"uf�����_�u}���	��_�z՚߭v������ӳڤ����Uһ�s u�l��
���^N΋cH��������9d�V�����M�Ģ�U}L���^�!R̷]oi�PIӼ"�`��Iށ�^9�Dn�M�M��Գ�g{ƪ�]|7(3���:�B#���sH/f�����)��l��%�Ѣv1��]�"<Ļ�I�K���iV���N��7�?8����� ��m�5�ەY�(�֒�/�KT$Ԇ0�n4bj��u���ѡ�0f����u��A�JO�%=�T����5�D�`�P��E!��0Y0&��7�BBc�(�4^_90��DK��%�I"}sLf�:��Ѕ��*{���t/����w<��]9����i��_
��S�kH2r+��Kf�'���x�g�0��_s��>xM�������+��B}�b�0��ޞF�����5�@�,n���}��_+�j�9' ��`ƤW�����唃跁�{P���@b^� �ln~�p3\�~�y���Mk�e��+D�1��XY���i��,9'J��Y�7��_��]�R�@^Ԉ���b�TH_Q��D�4Ka���AK=5x%$��'��Ϊ�Պ�\)�/�ְ4��+�]2]��8\d��0���J�"6?�'�< Q�S�ࣨz��=ZB65î:M�ј�(j<����C? ߛh�r� �u�Z�/��.�s
�uӅd�\��r!�2� ��yx����&��JB����m8<�X��lq�,D����'�Q�3�p���~X���������㎣KF��dǫ�q����|S>�lӷ4��Z�[?V��u�V#g�*�?���[t��br^�J�$6+�|��X���j2�G48���<.U�?����jC�f�Q��B�0f��^�t��I.&V%a�t���x�k�:��avy��c��DՆqtN�e�K�i��at!)��s����.nӎ ђ _���Om|h����/����	����6������){�f�x.���(��-r9��u��Obr/{�Hf�-_�q��mW������a��j��(ؼeJ��T[�&�:�	�( v)c$����4�KP�7�k�͟9�3�n�x��3<[kR���J����W7Y��[��'Y _��	$8��}6BB���N�e��S�zI�4Vm�����߈Eh�(���|��w��\�J��eN�E}��vT3�ϧ���(�?�M�������]:6�A��U���A��Ol�����Ա�F������r����jA{���)'ց��aU�@��aa�Φ�!���v����O���8�ػ[�۟�� 2��(>�Z�- �Z�[Uv�^�:��;e���G�!,�lm�9��
t��n �hz(������(b������I��mY>�*�8�q.j�)D~�(簠�����3�'__7U|��j���WS�n���;h�u�w�k=q=���F�T{aŧ�V�^C������]���lժi
����I�G3�f�t .:�xҋ��x��|�����t�r�r�2Ew��5�O�k����"k��gλx��f)�=�9Z�t�>��g|$%�L����z�� 7�1����Z���2�����VKsq�l������W�Po����S���D���Y�ͻ�_�W�\M{�L�{���q���ISv�~�M_�y����8���AZ��q(a�uX��A���>{Z+L�b�
�uތ��q�/��x_��Ʒ�q���ni� _���� �@�U6�8�j\ߎ�4[���}ԟ�d-�R=�X�~Up%.�)�{�����P�y��J���Cd�8�+��_%�a��q�KH��E��|S`A�hp��xa<�,�􌏾�m��f�N�6PX?��u�-���\�na+/|1�n|�kC�i�9�;�Ν2�/+p5]�m������0���)㱔�PF��zj���X��������L���b�㰵��)K�p�۔�?����JCvO�Y�wE�jg8�ʹ!3�����d�m���c��7�~�K$�t�g�0��L�:u��k.\7}:Q��d�y
�$��`�<��6�B&�y?�(r�8�UP���ae�q����r���M�T�q����-�Z��6 pA�-��5P%m$Ў���QJd�o6��[�����������̪]~Aa�����g& ��CZW�j�h�1;q!����Y��a5���6��K4��ݖ+.�!0_�.��4��}����?#��K�78�Mn�'���E�<���g��
�#�x4��(��kZ]��g_V�I��Ij�ﻊy�d7\V����jG��X73v����E����wz6	u�}I[�`����8�it��?��N65�^��+�bN�)ǁ B���h��NV	��	� ���"W�7��萼���`2�� �?�Z�K	�nF�nPK�:�u+J��<J���u���>4|Ж�ѐ�4����������MjgH�Q��=B���.������U����9�n�^�Dְ؃)|P�(����p&+�k�r��^F�_-`�����	��Zѓ]F�$ѰՇ��ѱ�_(��X�7ς*�t}���T�3o�)�V:D�d'�Ɂ�]��ާ�a=r�̬Ϊ�P�E�(����k�*�	`'�z՚n@�2�#l�m�x|�M�9F�3N�`'xU���rA ����J���|6�>�A�h��/�Y�h(]��uGK)y�k��d?>�a-�k�)��r�Y�Qt���'�i���4��N�n�9�Ǽ}�f�lC8Eh�V�Vw�Qn@Z;孺ڜ ^�C��B }g�w��{����]�3�@�Xa�v�D>&1�L��FI�^��[������ŷR����_0���%X� '���'�lF2�V=��L��(��K.u^�D���y�֠�.���V������?�(��~��ɬ��Å���h�"I[RLs�Q��H�MȺ��x/����ʍ��T5�D0��-��\�G�I隘ύ�m�sg�o�����C����T�����~8����g)m��i�f)���4��X�p�{�B�`�
���P�WW�F���d��]޾�m��Ј�l(�=���6��&�ʖ����M��&��3�^�q`K}��=p34Z�΅�����g`�|�7�C�b��z��pme�T�|ɏ���WUxz!�X�14y�
7�v�r�ׁ�����m��Ũ֕�wD\+�#W�D�?*(ŋK(Z'f �W�˭p�%.$$����;2x5�s����L����q��T-PkMى��?��5+l���c�g�o�8ڗ�fu�g�Gֵ`#7u�˧k
Db�P�˅��`�LM�o��K�m*.�!�CsU�L��g�[*�Ț���+�2a0=����z�y��P�������Rp���H���xR��R.}�����K}�0=_{��~fc�$	z|�[���ֱ��ӆD��^IA�& �c�ґ�h+�16����VB`ᮉW��AĎ��l����lC�d�7��������mj4y59�K�|���.Ҁ��h&�b��-N�r�ge\/��k���]p�P�P�u�C��ǮK$DWQǊ���g=����]RP�*�B��������FQF���I3�t5`����lh9�5�$C���;��zLfI��8a\��,@6<�ix��RqZ1ܖ�,�����#Ɏ�aE����o�˂�2�tI�4�}K��uɁAyɀ��W�S��V:�K���tc�^�/��HH�3A��я���n����k�e��Rh��'e8�[�0��$)��B���HSAf	h6_i�9�>g��mo|��5����dp���}�1/%4q��'���'�g��m9��۰6����A�2��I���9U��������5>��8�w:a�Q��ʇ ��8�W����T�[󛕻
W)��C6?A��s����(O(�Iƺ�H�O�\��_ʈ�q�=��D)E�,<j��r	&����ԩ�H�U��G�y}����{���#D4�jQx��+Z�N7yE0)&��[O��ʚ��gV��ؙ���P��xd��(�מ����ޕ�T�%p���xin%���j5���%b@�$:v�����7
��t��K��o�o3:hB��8}��������$�-��ջ3/Y�z��V�� ���W����2m����XC�6b|�๎�n�Ye=ȱԹ���f�ơ�VJɵ`bh�����GQy�k��`�ejy�R�B��
VҤ�� �̺ow���*�r�>�c��C Wa1��
�B^�����}<���`�c#'ZY�Ϡ�sԐ�hﯷ�XږlO����O�S�v��f��@���~d'��\����O������>���%�r�0kſ��Ɲ�]R�<�׸���u	Rn���B�P4�ȼ;���f���LFy�,�����GI�]�&��S��ʢ=�T@1�L���`�������dS/�@��S��7��yC���>��M7+�Z�à3-O�������yj���9.���?:H<Mu��K�f��*�p
y	�Uk9��vUf1˜g[�F�0���/��Ǎ8�P�BߔΞ�I`�чk�@����N	:.�v�0��W�.BU)�$����07�#���DC2���'�]��{X<�k��^���w��Q�m��O#<$�![�Y��\��$��o������X����i�X\�N�ӛt]���ԛ�w�s��`�  �֨����/iPI}���.[�}1"�!,���9�ޠ^�� t����r;��YҔUz�q%�^gE���@Ď;l��=��KC24 �P�`&�K�(\�W�3٠b�ߨ�6g�eDi���Ic�ryCU�Z�|R�ۭ���*ަkK��/T�֏I���;��V�\��]�;*f�ݜ��lDl�쫖QƲ�UYL����IO�Ҏ��X�*����85k��bĿ[�d_~�kv~�"
����&յYb,���1/%�R�`'�au`Z]y1K%A*���`�3c0��CELE~u�:�':���/�He��Z�y��L��Xh:����[w���D
�������<������+$A�S����R�ɰƍC��1cQ
���n�4bǠ`����.T��IB���?rEʛ����2l۴��<\��[��p��",3 �����8v��럅�#߳}۾d0
T&�\�B*��ͳ�
��]�X�Z���,�K�E�b���+\㹴����iu���/τ������������}߁��0�YHڀH@ a뎂��Aa��!��fN�#���,C��|]�|�^�_+���>m�{?�,�1�����%�-������l}��1E�L�Qb�'����M���Z�ۡ��"0<�*��u*�i��-���(��M��9�))_l)��J���4�Z[��b�zY(��󘩦�F�K�>z�1�h�m���NX��=Ą(�E�`��\�@�K���_g6��^������*�X�>>��0�-7�J�߶%����*T�����gs��~4Q3H�K��!�7,�����`Ђ
5���CJ���QW@�_����I�&��'(���D�`���:�%Wh�h��T�(���k���O�T�x�ߘxL��j���m*\�H�.Xd�`���8>u��ޭ�&c���3W��&�=TX�^H]A��!CP꣔�.��Jnku�-tb�M����5���G%@���vY�\��S`��;T�� ��=������Uul���tx��]sg����\G]�ԃ�	����!����;�SR^���5��ּ��iN���"lue)w����TΏ!�G���7�[�%#��\�� ��}K ꂦ97�#X��S	x
ϖ�)����tr|Л`t�}�wӇcܶ��4g���(8Hk��\��4�%��p�H�Ns�&/�6P;"��6q������PW�y愬E��հ���r�Y�������a��Z�LbfL� �����<.8�L�j��RN)`l/�?���y3�k^��`�%x�3�!��˰��:��
�/^��Y�P�Tw��˓za6�K�����(ǜ��+] i,��v1� ����,�@Z����
BZ��z��'5��	�G����ur�퓇�&c�|הQ�ßv�j��h�$����v^:��x��M3N>^��uu��G���B�4B0��1�(G���I/�G��_���hy ���&�X]�9#�G���;d\Qi(Ǧ��-wS�{��Q� "�ۣ�a'�5���S�����Zg֥��>0�fx��=ѫ|_�W������d�8B3�K���+�|y���03�1�T�T|x���LNpb�#߻?[����#1��.���d��.+�Ki�E)
��2	�iD�x:�tUNM�)o���"/&�I����L���̤�6]q�7㇎f蹳R�	�(w�A�	���H�7�(��M��'�N��.]���#2��T9o�iy/K�ʁ�)����F"��E���2#V�K����	9ȫ����¹Ӎjџ��&\0p����1id�5c]7����%�ky��:�u��A����!��Ⱥ��R*F����d�.v)�x��o���.�S�!Je(�bi�w릗Qׄ��`����*MIϩ�)�*/���&"k�%�m�U:$���ρ��%�i�o'4;� )dQ�k��~I{���.G���cb�/�l�9�E�c�����N�6��d�*3���� �^�^���[�3�36� ����~D��9h���bL>�ʚS�y��wq�R�DS��H�U�\��
�K�M#"���p�ı ;6��ڹ�dsX=����Eo�7^��F>�Q� Ǉa@W	"�5�"�D	s2�۴�k�y|�{���+�����2�;O�;��hv@��9�>�[ד��!�10�+�v׸�*?��#5��r��eu�<>�@n"X�8���< d��8;�䭜e~�d���d���OC n������Y�C�Bm#�jֹ\E��t1�L��g��V���7�pB�&+�H5�v�<zm��>��/�P�~��� ��uT7��[���*�p�q*���Z=�0l���-��F���G�i)��Ql��>Mi��1$��:U��K��SG~� R�&��z���Z�	9����d��n�4U &�l��*A��s�]C�?fC���GWi����L��E9_�ί޶�����%n.AQ֞<�e��m)o1������ۈ�<�iR�����՞��s�-p���K���Ę�sj@��^���a�)����o%'~��X[Qa����ɱ�$�{�k�ϳ3�DB�|�i���$�i�аZ�e%��c���@��a��c�@0{�B�
a��I�(ן�}�K���#�׼�;
����8��e![Δ�k�9.{�]���*��Օ���4%S�=m�zFrb�h#�Mymq��;���T�I��*!�e�Q�5�F�B	�>`T��}^�<m*���mr>�rU���?W�X�<�{?}/����.����Ũ����(Dy��O�[�(�nUk�hH	k#�o��/j��-P�f����Ր�e{9�a�ڲw�=~3V��p���4M�5��O�:�'v|U��pe����|ΓaI�/Lh�B�(W�_E-φv� �%�d�T�q����d�ɮG���^z6i���0�����R�fiPgM��K�t	h��}u��!g���h���\m��2�Ur���vH����dt��<,�l(
G�w��)�}�ҫ��\Vix7�aNb��A�w~ɜR����mN�Pe��f�$nbO��I�~]�����Ϯ��ߊ�S��O�h\��^T�	G�K����7<�s�~A)�O-EE9�����C�:��D��.�Y\T���s��QI@/����+�e����A)(��ț��{�Z�4��>�36���k� P�^�|���y��o�����W�-b|y��.�i��>��x��u��ޣ\��؆�2ez�J��Oe�0�:-?52KT ���:�J������hţ��:�1���5jcЫ�1��b0��q�|�T�
�;�y{H��1�h������}��uphJ����c+����&����rW;�ǥ(�J�Q�˳�>^���[9A-��hq�0fvl�ûh�
���F�i+<�=���1�I�z�sP&:���t�_��O��\��M/Z$�C�.�D��-e9ͯ�7��蕄(W��m QD�"���-ݘ�Ųv�ȟ������qN��dQ�VIBU���Y��mG�ؾP���Ak~��H��Xj<i��=$2������A�(��2�dm᳘��$�����tA�8N�W��rQ���c]K� �3.
������)51�Ǣ���<V��7���m=����N�[�Z�
�{�%�cQx\�H��HC�T1>�tEr��u�ۿ�f�F����K��$�l ;-�&i�{L��Z���N������bOS�MT	������ �����8���w��V�"�IRu���TB�� 5�`��ƃR8���� ���oPE|�xl�~ڏ�B�6~ޙ�9���{�K ߨa2�|���i�#T�K7��HO�֥��y�.b�Y /���P�
����O�����7�?�lk{�ǇD��U�ʞs�Y�;�ҀF�˾Z<S��(�����&���[ȴ��)����+Ve��ta�|9�.Q�ɏ�d#B�X�{N���v�ZP��b��i�F��֧����o����B2{�`�F�%E��VZ}�����-=e{�Ԏ����e�Ii-��� �P$W�YsV����C����Ѵ�wuP��!
D�-�	�5[+���7�D% ���$��y�r���QI�S��D�̳x�!����cz~��� '����x"��h��zG&���W~����eC�(�� G��aG�:]��Ӽ(P&�,ٲ�Ã�SFg��Nߜ5~\ <6�Q�yO��	�^)���O7	���b�(����%�*|�zɉ�5��l1��ʆ�wi/0��&6�&�_#{��;����!S;b�x� �z�����=A�\0�����Q�����(/�d����;��/�Zm�/f��@b,_e��R�<Шy����=a��T�O�0�� ��w�ḷs~�[��@� ��^�I��!���G	�-#����~̻�O	��I˻$$a�m=L�PEB�%����h�4�\H~��aNj�Q���jd�$
4K��Ú@o.-V���s��R�E��N���~��'s*?doW�1j�4�j9�@�~�_ 6�=�'s$a�P�LR�2eb��c�	\\2�k�W3u/�M@�X��) \Q�N�%�r�7��ۧ�f�jr;�<$[�[��l�����bv>�"��<"��NR�K���
����W�5>� C�3��0�
]c:/HZm��t6?y�%��R+EC�>�]V%��r�Sj���Jz�M�Ȇi5Z�"�.l�5N@ *9,;�Y����
�\WA3l��9�1m�{��$v#�!��ӫJ�jo��f�>�d�Q>�A�5�Q;u��Iac���G5B���$�{z:~�D'� 9(���O񦻣��Jo��ݺM����TS��x\�ɣ��%Z��LeA�$���b!ohp�4���@�Pa�����W��9ކ����I@J�]�bR���v����nWMWcL�N�,>��)�X����wE7�와.G�~V`bYH�|."�(����[��Dl-N�NA�����ezε�c�u~���jGn�%�q��]Ə�h:4"�R�ٟG��i]��Ё�ێ�M!��o�vs���J����(�_����wͧP�*d�5v��dD����M�9ȧ{��N�Z�k%N�L(���u���\__�ߣRf���$:����%��v��7g[��ԍ�v g�������=�������Һ����ͺ�.'����Ok���,�F�.&��$��Rna��MVa�7�d�0�\��[}Ȯʬ���|z\��[{�f�#����T�i�xGّ5K�ߑ�C����&��De��قz[}��fڿm?�)P�����X��l���F+	���p4�$�{k�������s��Y���Hv�Q}������������^����}��ڭǴ>����1Sv��,���M�WTCg;�W���j�Ϝ)rO�4 ��87�dL;�V��S�x[��f��"'ֶ��l�����ߤ������u4N���I5�<��D��~�5��K0WFh����k�$L=G���ћ}�Mxi��C�)��U8)?���e�x����f��昧6>�2hB��o梊���a��W�0�����Z��7����"S:�H6&>�ߌK�ON���s���W0="�Q��V�K���C�0�u:P��1��#}��Қ�~��[k dg����l*��
���z�T����1+�Ȁ"7��fd�m��l��^�vE�/3p�e�Q$~�M��܇D�w/E�3E��cx�m/XLmU�S\'����`���%�Ͷ�fu
B��0��]�3�5�>Z��b�1g�!\�eg�+@�Ǽ�å�P5h?�LY����[M{������E��뮋�^��g�:��%�뼕6�ibL�|�b�(���K�h`H�!Vq诖��� ���F`>`s|�sҞ�@R��W����Rν��R���k��:��{��Y\�L��R�pz|���su�JK���L�[,( X��<H��<k�G�$;e�jzQ��I����Y��\)�g=4�́���yR�A�p���ܲҀ#RN�4J�>��MV\WsBR�C1��yC�QU!���-����'7�Pnb��(�q�">LD�c�Wt���{�5����%���AH��qP��T64����њU=�Ǣ9� ��K�74�1_ә�6UՇI��w,t�<3��=�B=b�,�i-���(�H�Y������@	j�!D�
I�"�\?�S�ͯ�GF�ræ!|=�j�~�XxF���N}��N-oxǆJRɆ����q�� �`��߮ķT=�H���ٿ��v�S	�d�wRI��)�HD��3��T�Cbª��0p��w�M\�q��g����:�M5~c�R���8�������ފ�QE�l�'��t���JW��R���d^�2��L��U���=�:�E"G�{߃h����{��Ykҙ"B⍜�ԙtU�7u�!���uŕ�P�sir6A�T���KZȇ�˶O�wL�7����kY�"�p%�������Q��X-O��^����{~	���R��\�R�aʓC��>�����qɲ{����iT�dTu����p�t}Y�g�������5w�$�e��vzJ(��^�F��ω��CG��Ȋj��� Q�<@��v�/���c���&H�^pzF�L����xS�Z��GJ
dZ��8�k�����V3��h��3c�A�'=�+D���sY���A\�c�x���<���4�*�#!�����o\�7��|���nFxyN�P�������ߣs���]`�8�����G�ƕ���:ԥ�"���c��|�w����ǔ^/�Q�iY=�G�6uól��:؟@n��u&��a�������u�b?��I�|K�G4O|y�> ����V�_\{\��M^����Ѻ�4稈�m`M���
�xD+�G`2�e�%l�o��z�&���J_�ۇ.��7
Q3��SK�A��O����n_?$�Q�Ң/�}�ќ y��*�Xb1�R)}$��H7�F?�j7���}���fT	�d;�x[���㓘V�5��=@��k��wQ=����7�T��xl䁉�,�98���F��j��M2C����4�(U��S�V�gƷYu��J���;�T���ܞe=^c�
&uJ;I+���U������3]�S�N�������Q�����
{]���HǬ���s�61��$q֍b�q��8GSS�����<B����)�Q7��<��,>I$`���%(n�ƚ�&w���CYgZ�=!�R�1+��
�gܰo䨿<��� ��#)�yѿ�ֺM��_g��4�x߇�����?���?�}w]	g���g�j{�$�q;IM�*���B�����ߗ�`N�m�Q�����m�tI�r��"�{�Ȯ��g�MZ(�gVr%��k\�ma�ԝ O&��<&^�\��%?���������]{�5��^����0>ÚP%�������S����F�a_��Cu+L(e_��#�&.Q�b<y��|�t�٩�&X��	���~1WVd�S�g��U�a��6bl���	/�����e�&��ްؕ�ұě��vX'�>sſ
�z?�$�_n�d�8��pQ��b��!�F���x���e晦�|N\!Z����`҅�S�lվ*'"��{x?�-k*�Ę���t�� y�`�TG*�j7=AP�X��j$|pn{`��e��K�}ht�̝&J��n��-W���_PK��2�Q�0:�H�T��ZeI����y�W+���͈�S�P�\´�Y�f�.=7DY7n��Q&&��<���c�4g�Q�P��xZI�W@����b��Ӣ[�O��}���^^CQ^0M��~t�Y=]mF���M>[ýM?�Vޠ�pO>p�y0�3�@z@���hE}m�d��hql��
D@v��3c�ml�\yE..��{.�o���ۑ�A��/�}5��S�,��-��Ӝ�Ȳ+#Vf��A�UҔ���r��}#J����l�����!O�O�<�j!w���<Ě0����r�'^)��+Y��F���di��}܀�qf�a<Q���]���;E}��/�f�N�ݣ�Бq@1���R��W㿧�7� 9���t�������h�}�1@��xl�Q7��1�D�՞���8��O�!�L��2��P�q���ȕ
y+k�|u6��}�i~/]���4��9O�`�E]�)�o�M[h��@4U/Z��b��>a����]��$\�?Z��A*��JЍL���Jo:��Y֍�RI�7� ����=���,��=N5�A��9&�[?�+�o�������w��@K�+�e��W�w�^�&�d:oq��33���?\��ڙ���7I�N.H�r2�+�����Zc���?�wЗi��1�04D�f�ҩ��P��%��~�V�|��[Z�r�P��� �ήc7����ڃzK����E�C(�_�j�}��o+�mT`(B�prhd�f(pN�izx�D��Kz�ᨰX��OԻlk��8�j;��9�*X-*.�]��.�7ǹ(C�ȉ���<�F/�4���ß�v�=��$�*A):E��-�S�ON��>&&�8��4����w~oi���`U	v�F�־�#�9���"�M�X �L�1���W@����0B[ƃ��@p[���p���zI���^��!�lXC���)��heT�6�F
�#VSk'�l��>q�0���S��E���(��]]˼�!�i�!�����f�J\ޔ�\�{V7��!BP�Y�P����>�#o��JG�H@!y	��E��=����^õӷ�*��آ�x��?�������w�Q圲�WD�jl�A��n[^W��K���SK����'��\}42��)l ޣgk�+g��[�S��E��׿�
�Ǖ2���p+���08÷�T l��8Z��}V��+�2�(D��z���n6�!O�Չ"�<k\��UTۏ@-�!�+ �'T��lk��T�[6�-J�vKP��ԍ�RF�q4�<�w��Pꌫ�ð.@��W>�1�r���H�6\|��E3(�^ @ �S4���C�vls?�n����`FN?����qw g[�z�C��q�a�;}�%�\V|@�\��E���c񄄚K��x�ZA%
$����8Ct×��A4�GPU- ;�Q��SD؉|̇�t��^�@���� ��X�F�g~\�ϭ*�}�l���Y*�/��ȿL�Vzc$�0��w�?;�"6%����s�64�e����J�C՘Lᚎ�֫��������ħ�h��Ϯ����/�aNi
�_&-�lRp]V�Ծ�\Hb��B��"RL�vE����oy;���b6�NR�'��!1�5�'���GpV��Ɔ�pZԐ�L�?��S����9�V.EH���������x|�=6����*�d��??�4e���%�=[c�ň�ˑO���VF�n�Ij�v�o��u^�x�}��p����+���c��?FZ�e�̔��\g�1t���Zl��3�C	|�����Oip����P���t�k#!0�ǆY%A�Hf��}���Q!l0�����ņ�|q��R�L��Z�� u�$�v��c�m^9�`����j+�b�" ���#��qU��~��Dӣ�o�x�W����J�ܷ��,l�%�L%��F��շ���؁���!}5��X�Y�N>��a�3Q�n�B,I�/᪰Ue������@vUV��jQm��xe�3�1ӄ�C�uc��ƓG��1�S�e�������%KޙT���� Ra���(��|�'�Y7G	��c]!�Y�{�%�f3�����,�I�����K��)���;+�s��?ǑD��	�j`{��I��Up,�Ko�������䄚�9�~�w���6�����BXu[�v[�:���bc՛,�;J9ԗ�Rߋ�[��T`��*�>�&~�
/:֑c	����	���(;�_��b��z�A�x��r`�W��E�޹ކvs�$�Q� ~�j�Wv)�󯱡�B}�F�r�̟�Sq�j�ǚ�����=?���M�E�I�4,�Q=՝��G���g���Ӹ�@��Gi(k��/��$�jڊ%��ܤY�Mҁ�9���0�(�Ќ�ʟ��ρ9i��>:է�ƕ�9*�X���	O\^9[���N�d#����=.������Y��|;�+�DG%�g��t�h5��r�@�$�۩k� �U�����l趞ث��3�S����oZ�֟�p���`����" �%�����L����V$��@�v�FW��Wȍ����O��L	��?��7��[����4����f�M��n}�P����񥊪��Jf����sp�'�����|��)'ax���E���:����P�����s�?k7K�>-./����0��J�0E�ͨ�6��7Q����<Ղ4dl���*���	Iǀ7E!�g_bnl���x=�߂p~���b�b1�gdP�u��NӘJ�4�lli��E<<��������"�LV���kqET�KV��	��}D��/-%�)�_Y_=����h�Z