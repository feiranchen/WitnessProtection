��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f���*�x���!�֡*����G�J�K(�T�haCﰦ�4�af��5�_tA8�QO`wqM��0@o?�M�+-����8%zF���@M�$��-4��s����$��sp�-���*����z��2d�t8$g���YE��;)X�<1�?[�(_�{��ǉJ�oG�g�����v7AC�O��I�h� ����`�.���;58�%����÷��G��adt��_N�6��<aFg��ь����Q2�����C῭ن��%�i\R�H��c9�LdZ1^F9�Ia�Nx� ]V��&%OU�{YSy<d3��!fH�ArWr�A����?��)��"���vbV�f6��#���P��c����Q_i���*��'�A�Q���Qp�h%:?H�4`�Bo�x�9�_ ������^�dS�9L8dF���Yy��{�с�<����'i��-�\,�{�{���/J,�u��D��d%h|s-�3���i��b��+���|�q�bO�!���]+���^5��"�u����q�w
P����2s�Y�j���܂�\}�LA�ʅ�:~I�u������@R�x�EN����$��3�uN�xnO�ۭh��9�����cy(���3�R�.�2����l�����6� >������`����y��׸<�nJSO�������~B�x��.TR������]�Q�Z�@}sRz@ Z�
K��yA���'?Zw�k$����,��V�[�_D�~��t�{�Z�?�W���*��n�A�3�;Q>,��w������.b��W��b�E/�Q�~2}y]G����I���2��4)=��+����z��:27$^@����h���8���n6E���!w�.8���$Et#��Y��.����5�p�� ����HQ�@��f�9c���+"^�T�;�GD�*�F����(�Lj/�hV�~�j�7�#����b�6��d�uR1�O���,��{�����Κ�N~��氒�j�Wc�S���I�� ����;��QPL`�Ie��@��1����	K�=��X����lw�w�����v�ټ��Gc-Q[���Ż۾B��5�'Z�y �-�ր�t~��  SBx�'�WCd��*X�ʧϦ̢f�>��D�d2N�6.��;����AS͆������=���"ݨ���#.6�V%N�j@y�3�7CL`H�k�nB����x�q+���jh��kq�Mg�_I���jգ�|���(�Q)�3����ɻ���C�x�J�?a7@�=m�B�����Y��7[u�|�ޞ·��F�ڕ��>��%�y�բW�E���q��g�T����X���˴��}be���m���O��L P��]i��#$U!���G��1�4���ih�sNv��'����X�<2�bY��ߡR{��#����������b �m��(�l��D]>�})!��hp������g�=)!X�&��b�1=�#��iK�2�]	U֣v���WWhL;���n��Y����ʩ��+��0:{�C��b~�;%��
�LaK�3���h���x�)�}J°=R
!\�ot`َkcO��}u�|�?��ag.#���靗�Еb-k�֮�wp�~�:��a�ۍ"����E�+�f�}�ѾI2o[���iq�V]t;�_W_1�v�nB�z�s���X��s�Ɂ���*�������Bf�bFH����&�q��V<�b�+m�ò1�(�NS	�c���F��t8Y���?�$d�B���`�GL��Ht3@!�ău���Q~�!~��I�B���O#�򽦺�k{��S"(�m���Dz� uɺ�-~�y��i��u��,�	vޏˮ3=��ǳ�U��������3�֒������iK�Cg!/�_bÕw�����~C��h���{-��]�+g�� m�@0�Kf�#V���� ,.K�}�FFr��y���Y݌�d����[��zC�;��c�p��0��U��!���"�j��>�U�Ӷ�R�/1�")� ǜɤOJl�H3�b��5�ޑ_�v�k�.��������&5ȉ�H2w�c�8S-gL�Sd�Fˎ�o���=�I���Eayڽm.(�8�S{�����d& ��q��9�D�ώx'3A5١��_��b9��L's	i��[���@	�����7΍m�%s�W7������S��Y�����_R�t��KL�!^����<�ݦ6�E��~�����UiH
�)?�v��o͘�g���U��z��" �/��'_�23%�_�#�����9�)�<b�{�=Ya�G%\�h?�S��7<���z^�_�8J0�L������X���(��cq�9��K�%G�oˍ��r�9v>�r�V2,�Ff�DGKS�q�s2TX݌.��X*K��l�KzQ�7{�,�hn ���y�c�ف`��OSfkY�gL�Y-c�T�~i8��~�V8Q/=�f����*�;8.�'��@��$t��'�x���H���;=�Je��W��k@qg�.�Gv��M8^X�*��X���O�h����u�^���C^��;:���1~�T�,Wy�Wh�Lf���7��ԩ�d/���X���fc���#Hb;B�1#��Ι�=��K��Rc�g�W)���5�&׃���ǵ�/E">:S��ѧ�yC��89w=d�J9((g�u���Z�u�c}�l��3���Ŀ���ښDM�S�<a=q�g!v{W�_�j��
_�����N�?�1�u�N2����|KJ���L?�k"�,�vV�&��N��a�`Q8r����֍R|��`/��8�	�	Qe��ɡm����kI|�M���%f��f�]q�8`�c��R ��|F5��VHk,�Ko���'ز�ʘ��AOj?Oc�6ȩ�=g������*w���lDԹ�П|��o��c�lYf2�2-I�3�>f ����ZƗ�aEnv��¢췪A7A�]������I`�K2��6[%&�3����I��Т�AV�W0:ݣ�f�@|�(��>(ꋋ=��K0K�2�K�S͛�F�-BQ8�!��8����j�5`71���$��9c�>\ĦZ�0�O�Ev@Űgs�gm����m�^�����kK��M�Rz�:l>ھ���iW�ϹW���������E��B۽M��e��R��R�,%}-=6��Gަ�m��N��pB+�Ɠ�w~��/>�|S�g-ETk0r<�_˲��g7&���Fw��*�㎩�"���\y ={�T6<�z.'��u�H��?L��C}����>�q�A�n�'�pɿ��(v{�D�h1Cg�치����f��K& c_�^x�Կڟ�i��-�� ��䅬���/J� �Ǵ1%� "\>tª>��x�'F&�c�ǸW��:�ST���$e�������<���m��p�ӽG���m$�'�t�[�4B��u.�t�(FV��Ҡ��Lu��鍶]�� =`���㈾�/`�ˑicO3>N��M�(����C�M"�4??� �8z��<�"�n���f��e��ܮt�ջ���g��s,�cg������ț��:�3К�(�/�����VиW��{�6����.���u�C����q[�v��O�}I1EB*�xzZ�/�����mlUoFO�H�;C�VA��OVH��3�ӧ�(��o�,3x�,�|��4,��$G�*E������z�ݙQPU�}k`�^@d9�!��Ǟt+�q�x�ΟzΊ4�jb�j���W.ew�2$�j��}�O�i�������5o=ϦԨ��,�Lc}��-��͠��A�l��Y*%�o�|�
�� qVV�K��&uiSwr��P"c���%v��-5j�}܅�>c�D"L��s���I����>���U�ibK��5kT
E
��;�f��P27�>-��^�����ZX�����ѵ=�)����q����ҦH�S�1#�p;�%?����rW�/���)���͸M�fٖ�on�5(��"�Pi����[�������^Ғ*����EK��B�H�p�tқ��}���O���>!T.�h�.8��K(�X3�#6"�~�O|:P�L���X�����7�AT#M�c�=�ƗG	�����>:�Y���qz8Y�š�!�~z?�)���Ŷ|j�jeJ!���%�[��K|�M��ge\��AQ-��1���($����Ê ��E_���h�c��,���xW�)L�+��W֔��GB{��8�%L\���<a�;tY�� RkA˵?�l��8a����������8Zv�X ۙ?H�į�����N��@�QT��8I`(2��1��O��՜O�`xzs"��bF���o�A���eG����;�m�I.T��ķ�����f�B��_���р�G.���(��'킇���=�q�]]O~�k��� �&����!�����N�DI������hW�7�u��A,9�p�k0!������k�<>���8/�j���7p��?��
��N���Eov��s���lw�X� lˌ7@�+�7
)S*cPI��̙�/|g�WLƀډ��B(���L�Z+	�����&G_U
���=k���ȼL-��=���I�65�C����:3h,��R-���\�����8.�uq%�ɵ������/%��
3&��뢙.-���2�:-A� �RY`�ý5�����?b_;���B+-�>/sYy3;'�i�u�D�m�sc<������	�!��B�mW�t�
1E�A�X6l��\���uL�V̲�5*g�� �V�uIs��^�豄�dl��]��)�4o,�V �Fe;��p�D}~$�V�`x6Dr\��v�W��ϰ,�ö������q�!W:��������};��oím�9���)����Tbt���Ƞ��0=& �a'ĆZ�Ռ	��1�s�8�yK�6��T������\/2��R.^��x�[WS��p��\��%��%�_:+�;x��O����c�R�87�pZ�lQ���w�K}�-�H�^�Z���jm!��$�H����/MD���q�_�E�=I�8��g�/X����e�$�c��������fM= ���x���%�o�<旟W�Q�n����y�`��ߟ����	!��� QŭEr�T�xj������i"^3b�s���.d^+�d���n����;���+,�:�L�u*�a>�o�,���d�/�Ip�O>s3�r_��c��M2OT���uK��A 3����ƕ�ٹ4?2�9��7�O�����{]"Q���iYƬ���.���ˊ�W��th���^�\���Y�\���Y1�V���.F�t{��?T�������Nq#�4W{Z�[�m����x�<|Uo�T�9Ğ��_5޹��ސ�7�o��=2�������gfn����0��֨�ء�̅��+��IX@,�Nm���5VĮ��c�ś�H/L�������l)/W�7�z���A�� �j'[��M}�\JQ�Ϣl�b�lF��m0�0ܠH��\mq�1��O[r�g�Y;Q�<��+l��WƃH�]b���k�!���&�p��cZ�Z��w��M)�{s,:I�O�oBʥ��lJ0��.�l�q 7s��}M���]���
Vu�ւX�w0��X�*�"��Q�� ",+h���uJ�+!�Rw�c�JNd��RE��a���
ƶ%2J������gDm�A�O����W���n��k�����%�m�8�l����[~��U^�0��������z�D��T4�!�?L+���Bܲ �c]�Σ���Q��:�$J�C4�e�f:�:p�m�r��h�djb�g��I��4��o0r���d^�2��U/;��`��9�v��ͳ������_Q�!k� X���g**O���^��B쑯(<�4� �/��� ����w�x�pE�3~TH'V�W ���{�������`���{l<��X_�k�=��y�~���o�@�� i�F2�H�r���t
mۓ*e7<���(�C){Z^4�}�"O�!t) %��}�	T�C���$�.��Y�E��	h<�jީ}䞽�Q��$\�)je���Z\*�R:�i��l�/̥־2ד�M�ر����sx��qL ���r�%r�Ԫ����jI�H=���BV,cq���\~7��Tێw��(Y�g/�V�.��Z�Ѽʕ�pNr셹]1c�x}�_K9M�����l.��q�`���+�u)Qܺqr��j=�7��h�����F���\���Iׯ� @��N6;)�>h���>�*�AY���M=��s��stR�@�Q&�5�Ü.62��^�	�o;���*����E~!r�~���H�-� �↟t�,����%�q�O|��.F$[,��4�&������x�.�Ρ^�m���Yf���J�e�V�aD����5ΜmZ+����bp��E�%��I�b�����8�-&�����@WԔh�.u���u���r/YU�S��Œ�=3j<�*�kJ7�rUm�PT�#�!# �-s-��+,8�����#��G����|�����VcSi�|���Mg<��c9z�^��4����0k�&BH�M7�cI�x�7b��)�����&rd�E��p���vё�?g�9����\S����c3]��;s�;���R��X�m����
�(�����xNN0�&��%9���á}K��U�e�ΎAD�?7��$��p?ӽ؛Kp����l��-��Vh�a nF�-g	E�~q�L�ksa�ɮC�jk94f�e�ժ'~�O��Ҙ��j�єv%yboS�����k>�BK;�;%D t�<���Ŗ��X�̞Mi�X�9�?�*�g?1�|WE{Gt0nv���K�u���I����O�{�a�#ϥ�X�k{�i��3[_�2��wTNm�m$j���ET�ۖ֜{���M$���` �wJ>���շ <�o��ɉ�R�ŠE�C���d�	���O��>� p2�ĆJ5��,����C�{�Z�EivEsQ̓���y�:��Z��"!����\����JV��*p<ޫ���3qb�yrz�+��a�3�'�vQ��m8��ϲй_g|��q���ԛ/Ҳ�������-���d㲥;|��>��