��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T�K�b�;�m0�!����׼���	śCqe��R/��z�z�$rf�����y��7��e�h��Q�Td)��+mx�GB�H'S��{x�Q$��!�b��5W]�,OSo��zA`YB���!٘�p�HL87?s.����,�����/�a��m�^Rһp48�.�/�-����b�u�g^�\���Cf�uV���7l�H~#Ʊi2��8#[pU� �m�S��o�
�D~f:���X����z�� �L^��^�$��	�q�	(wV�L�I���!����%�hl)/��K׀��-�Y	�%��^u
����|��� 1=,s�ࣵ�$q+$9U��5o(��	Q\�ަsq�*XKqᰢ|�W@�ߎ(e2�	�<&UXy��X�<qj��6Z鉲�x���n��q ���Q��k;֏ R��p%��>X���57�,C)�$��-��2e��t��!�h���#�֓i>@1<58�;PP��u���O�ݮ�����k�D$�#��3�Jy��3������Wzgef0x�0��,��ig|1��!E��7*b̳Ͻ����HXFb����Zl���J\U�ᗳ Z�F�F�K$��|�;��������|{(�}Q�J����2s_�J��i�z�#>j��ļ�/v�iEDb�%�#1w�Z���1���,�o���&�L�74�C�t�v�nk˄��j�M`I�@�[E]'�1��>S��\�SȥB@֝���"�'���f^71��\tx}�\u���DT�'_��!`�ߖ� �b"��v)m��X��iQ\	ƚj��mJ�b��髠�<3[n���j+͢l�~�=�%=_G��mW� ġm����5{��Ӥ�N8b�ٷM~P��u�!0ؒ)o�>���_�\�W^�,�Q-h^�b�z����7GTs�&�ǒ� L�x��-���
]e_5�}m�iѐߢu2���8"������YԊet���7*����q����ѝ$�(�;�qFJxd��q#@��I:��$}g���-bď��p�ܝk"�&BϹ���j_@��z�����Dr�o������+,p�^���^�Y�� P6�Q�2!,��7�$��E�����e��8�
�ݓ�Hר�q �Kaѕ��d�k���ٯ�*;��CU�p2`��_�����H0"�U1w	���6�MTI��!aUO@l���Mn���!�V�C��ϥ�*�,�j5�%��3ߖ4K\�h�)N�Ű1�U{�p9'�L=uõ�HȤp�m^�P��.a��-��1�-�_�w��'�]a^��G��{��N(!��`T����m�&�@� c��wYZ�G�p�H���6�o�qklc��?S��*��m���/Ն��@;٦|h!��_�I0��m.�y`����F`��n��:Mc{E��e���$�8 S=P�=x��yo���v|�c�;w8����� �%E}�_	*	ͬS�o��e��HD�{ݪ4c`E�䖙b�$!���L���}q��'��`�U�t����l�]���N����As�v}l�f7�tމUf�=�T#h��x��G1)2V����=@N�fM���ő$������9��NS͗���r�����<Ƒ���M��_�������B�
��|���\hBbX�3�$�Dl�aq�e�i��Mr;�DI���:M��@4�[�΀��������w���мѼ��z�ɐZ����LQ�\�����~ ���˃�WL3�t�5�d+k �Guyu����dVa��~=Q��V�ŵ4�5GE-�}m
�d�����qL6X������;�ft}��q?��4�uŝ���%�������}�
��DU�gc<2;�,/���GIa�����!��tC#eS�9����%��pw;�6<�͉�"�g愻��h�r�o�䚏Ԍ��-�!J!Ʒ�C���=�>��O���KjF�3�����ⷕ�x�u�?3]�'"�'�g���(��=zf7P��ŏ��0�TsY�Lm��ϱ@������Y�P�8���_���y�C��3��\�IyHL���}��T��?rHe�>J� ��[��K0�O�fh">��8�{(�=T��!Ő����Cq�t�Y�Y��u��\���k��=�j=�=ң�^;�.�&��a�Б��%w����Þm��Q�"�1���t$c������I����	�E�b*�sݴ;]��w��]��:[�;����$!6�o3�=�Mי�1�"z֎JOv=���*>�k�}��!�M��ݔ}�\dΑ��s�C�N.Á00a�)����㶞E)��U4��Q���{~)��1��4��!F�;nExug�V��̧gj��������گ�{pSN$k�?���t�΢讠�!�s�)H��R t�T\�xDCO~��+��D1��;ODfv�K&���2G�^�h��� 5���{!�:5�p����7ۑ+������{���g2e��P���v۸�vi�ȹ �M�&�!�<�	ژշ?���s�*b�>T�-"��J��O@�7|�
��uJ$ L7�FY�)Z�%�WE0��j�{w��0�z�}�%�Uy[��2{����w{?���9�������0S�p㋨p�8�v�d(Tmgś�KI���C�/J�}�]>V;�X&g�'qm4�Juk�kܳ�����?6��S��Q
��p����R<8Vz?�����OIQ�e���N���0�`n���J|�[�{�pVT��4�~�{��Y��R�q���q�(��%�I ��w�pWy%����TK�b%8��VS�A�.E��b��!G�C�_v�0�|C;�ʛ'	9��?���[�"�!�t�64�����B�4�
���*~�_�3�0��W�<�ЌR�B����~~n��a��	R��㥛W:��k#A��ΆG���������V��C�F|�]򵔋5��6��Y�/��k��m�{&f[�m�w��^+�+����[+?��>݊O�}�Ĉ����R߻q�'ԂۜX?w�̼e4�!�sˑup��ݖ����6(E�p{�ip��C���h�=���/e4�ˢ*���

�EFs���ż�9�����38����e�_�M�}_��d�Q%Ƶ��Ĺ2v�f�a%$2̞�^[��X_Ew5U`'L,y��a N1��Q2�,�N~�@����_���gǝ=�y�(�?h:��A�uD8���jM�O���!���-��-S���	A%q��0ܶ�@��$��ZM��	ՙ��V��Z�_�� d	�%n������	�/�J��W7�5�eB9y,U�M'w�[���9��MAa{�Oй����ac��e��&���s�~Gw6���c���J"!��(�����j?�ࡐ�^�N���,��M��E��Ѕ	�ӏY�4Ğ���v_�w�<�!-�ٍ])�l�~����
�t.��+�Ez�zfB܂\}����_�L'��m-М����+�
|��$Գ�e2*���H������9ް>���e��S�]G䭯�_�u*�3��u̒8z��> ��5Y�
��p;v�����+,�Y�`����I)��%�ф#�Jn�f��	|���eo��(���^�)���n��ux��!z������O����T� U�YJ�_�H����I��ɍ�!E���
�ҳ����8��D�ޕ�\@���B��Kc�M�Bl�o����rsثFl�U���4mk�I������W����A54�1�j}1�3��<�i��c��=��m�]�u�Ĝ����I�C�GY�(S 6���ދ
hŰ5�
�0�M?��p���i���!܏��M"g�.q�^��_�Ĥ�oH�.Λ��~�A�;�x��y�@����2p}�.h�UP����\Za�K�x��k��/8"�c��N�
Z1ɧ��	<mjg�w��4��S�	iD����������?*r��_��<�y���!~6=�qp�	���bS���vsRA��L���<nل��"GŹd6����K��a����lۮ#r���]�q�ŏZ�O���Zˏ)+��a<�*�����#��P��?K�`��mR<���pYT�q|ؘ��� �',�'�\��=_:é[�kʍ�|�GDB��������{^��l\��$I���kA΋+�7ԇPgA�;���i�1�o�LVT�H��AT)t��P��J�������[��enN�Og¯�z��3IK9���ǅy���c��zf��4�I�1�=ߊ��ÜI�~���g��y|���Qۤ�c`5��*D:�����.d�_l(:�9���N'�}��9��3=^��N �,���S�W,{3|p�f�O?G��~߫��Y��O�^�Yb)li�������:1?X�'kӯ�SB�~xݠ�YC*�s�jQ��OiV�#���n�eF��#M�X��83�m|�V��1QY�p"z:Nd�.%&���?Z���=S�npDn+�(��Xhl��m?��L�."�@2�V	��#=�P(|�O*����w<g��9䙊7w����c��������^��Ν�?��o��ؾ��[*���͖Z��Fiǋ��)�hs!^^����մ D)�̀Z��=��m�܀d��V���C������M�F�c?������(qV��K]��Q�o���'�������N�:vU�vV��&�>K�/NKjp���©y���?0�-``��3��I��l�7Z�U�f$�7Tґt7���3T�?H�;�g����b����eM@#D^b�b܂l��鎼sh~���3�^�,T��o���D�8��ĩ�k:h���F&LҎ�D�a s�����1�3�eӥ�o�� 饯�pZ錞��O�d$y	���_�^�M�/��ίa�)g[��T���YwR&���U�R�g�
)鸑檧�$W�~gx'w��fJ�d9��,�I ����U=|#�#;�"3YW�R-��xL��o1���8d��d8�?�r5��Jzu�s=1����c���TX��:(�I�u�R����_��f��h�-VC�N�A���ƻ5V~8�p��)
��oz��A������ɿ��!DRKV/}�L%-�D���������<ws���+�c* ���+��& ��J�����9�=��l��,9dhk�8� b�6H��>�3�y�]��q(\��(�p�ӗ[��t��CT�7��_����c�K��L�$u�ыw��K-#UlS�|E�}=l�"�>P�&(�t�{5ҷH��Y�sn��q6��Kk�'Kh�K~��<�N�	�E��O@��h&Rn�F1��T�6���8ֶl8x���ɡ�F�����3$�[45`��K�"��v-H3���/׬l��Hs�0u��oOh V���}���Zi��\c."a̶84wgܲ�2�B;�rm���L�[�����������j����;���މ���[��Ltdx*^]��!�f�4
��wZW��ԝ���L�%@A��ܾS����P�X���)J�����$�j�}<|RE�7C6��m�ta�ji�m5YW��ַ����.��4�NS���W�p��1gj��x92T�O�$�g^��R��M��tI
 ��?"?��2X/�o/�vڲ��0rD
=�B�^L����ٕ`�c\P�y5��RL��~F�<{2M�-�5Y�V�OU���$�b���}��j"e�[��6�\�Nf��8��g�ŸF9н����S� �3M�?-N�LV�駷d�I	�e����F�� I�����1ʖ�J�/ �/��׿�iAA<��Z67� Ȕ�K�؂"
��T�� S"
���\R��/�7�����i����
����&X��BTݥ`ŅH??0�&�t����1΀J���.��J��W��"��� `���8Qբ*�oK��\Γ�@�����_��#��	�.�	3�/�h?��r��-_����)+)��
0T�r�j��2`��}��5ٝ�(����i'a^Hy�C�nw@���P�SSᛴN�%�7�;�{���BF�$����N*�c��� �����>=��Z�N�V`�Y ���M~�u��p��<��E�bc%������I��<<S58љJ0N+CT �?rT�,壾���_��gK�z��${�'H��������)�j���"w��������,����n��~���|:�Q��������P��{�"�{����_	Y(�&�}����L�p����3^,p��ĉ��1�俽����'8�[��*2�(�[v@�W:��_bG����;z�Ύ3�B��=U6��	�Y_*Q�o��z�V{�t�trg}�]a�yBQk���^�I�"�\��Iq+���.�<& [���,�n�p�-UL�Ň�
6�fAG� �� ����m��A�	�s�0t ��C�@� 3�5���*�*�yE�C?�5Eh�	��X����%Xʶht6�Y���hN���[F�2��*797��WXVtN�8��	��R�#�dN��9~�HH�B�ST��q�?u�w�-�qQ �o���El!��G� j�.N��<*A�5��	�w��[�S���y��֟�����Y���K�l��n|Ė}Rh�|�~�AY�	����:�L����6�Ī�:��O:^���u��^��՚���dEr/�m�@������Z;?�%V�wd�?�m�O4������G}+nT�̀��oP�@�<A�`�+��{4��=�Y���iX����*2�@�\Hg������3w�T'8\��X�������eл���+�S��w.ϑWj#w��L:Ӣ	a?~ib7��B�J6�����Mk�Ɨճ�w�;���� �N�����B�CI��@g`5�&�"�����FM�R�`Y砨�����w�h/q��V�nt�0>�������'�B؆��:��^*��)�