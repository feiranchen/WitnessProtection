��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ訯.$W�7)�v��_��F%/���٨���)��?_CіP�XEmҪ?��������[VpQq��H�#�)jo�A;^7"s �5�_��R�_��d�&�՝ELu�|R_��u�D ��B�(������VI�nW����Ы�MT�I��\��@��S>]I�K�:�E�a׵תQ0Mچs��T��Yl2�Ջ�:�?��w��X,g����޿��0���n��1߷�{�����|��I�r���WOX�PE;b�0�PHr:��"�h%�='�*�ǺSR�A�h�q��F�B"����7��Qf��!��z�5G��bEdn
fy�Lx�·��`��E�Y����V�G�d�tQޓW9�oͪ����KbU���E 6j��G��訒<v�|�te�%���02�ߋD�q���V�7���C�VrHb� Mn�d����(�L�1�a��鏁��*H1��R��dN���"��:�9e�7�*�P<��	.���������YQd ����:t)ﳡ��"omy��4�P�NA��V���2��y(F���n'���ř�ðW�f��GP�����Ѿ���}�8����Y�E�`q}U��G{5����eM�F1���OaAюd����=����,Q׉�����:���J��X����oΥ�P��g��wv�&�K�>����ZH7ύP���-����s��l;"��m�.='��i�zViʰ,�p��gK�g�s2�*� OqO�Mۭ�ltQ���l4���.E�wpES��*�~C�F�ޠ�;�ٌbN��"�ŽSY�o�W��M�$�(��J�3���/MT�H�T��W<��D59cܔW�Sl�,G�'?~2�����:��X�tŏ�@��v�EG��VL�jԌ]���_�����Z^(f�7�f�N���D�K"]�����Y���p.g�o{YD��~`�qM83��db棭�Q�g����M����HO�������M�m�/�G���N�k�yu ��Aib�^���`��q�!�����q�؂^]M�UY�M��.1"F
RFϣ�QO�10�{�hq�w;�`Ƽ<�����"�У�y.}�H,��G�;�%�qZ����9@���6ͅ�Q�U���zb��z�ak�=��$V��%g�a�.��Cr��K�'k	7 ��kR�l�H;�;W����^�����T�hW;��0�<u�g��G���J�&+H��!���x�$Q��Lq	�J=Y0��ץ�3���i�<��>��B�3;:(W,�x�w��XSY����|�f��/G�#^�(��8w)�9��i�S*	Pb�ˊڋg�Q�ML�R�I[^?b4�p�w`����&��{T�|�!�yyCh�FaP����FK��)c�3)
���W�V�D�.��3cx=���d��s}&ƙ>�L�p4�j��(vE�ь�a��mS���)(l�Eބ>�VR�wi<tN�İGo����wݲ[f�4��<�*9H����m����Q�HtQ�XW�"��.���i��)�hD�'�N�,2��X�#�F\�'jE4��ɑe��1���K������T��9�9Ѳ��z��RX��W�D�`c���� IY�N1�6�sS�>�g"2Y�t$#qs�ۙH�8vW3?3��%��h)�逐{��ܦ��P�^GIdk��
�p����gك
̠�ɖ��n����Q�b�S�g�)�Ռ�wCc)���)>�X쫕͉��7u��K3n˪�b�޲�FZ9GM0�k��S��|��l���ݷ���_��K�nB�A{sB����CзI'��}�#���ʓ��(ۊ�wzQ����z${=�=̢�O��*Bq�h��(C��]'8{	�����'w>����:&p�Ux,RJR09UϿ�P��\j|�x��Ǒ��Q\�U쟋���:H���������-� Y�蒑��h��]뢛z֟���$w��*[��Iw��Nu���#�ջ s��ghB.g��$0�U�,��㶼x���1o��$�]�|�k��l��0o��6n0@S
���`��4MS��sP��̪H��
�=bMp_Q����b��[u�kd)Hp32.���F ��ͪy�D��׾Yo�w�d�N4�-}p���6�t�~w�V�<��\m�FV�/MN1.55�A���� �E~@w�K�?�W��%��!�Za��PC$�xpx�����e���S�)E�03�fF���=" ��)�.lŇ[�'��8O[�(#B�(�k��&y�Y�t�Z,�q��hM';KT�>��E�b�#������5V��"-����2��T�y��(9
�Ƭ�Y�-.�@A�*oK/���Z��5TU�W�]ո2��K�KuMO�I�stv�8�dD~e�'.I���>��wױZf$�1A��G�M��D!��>��M��-����,�Ko-�����w�Q�e̺8�ԥ4��އ6��ݎGB�cT����`�h|F���ł��B�(��{vò}eꃚL�qqܗ̇�[����`��J�@OkHlI�o�o�rA^$�e�����$� �K�v���	��!�yy�?�h�e�-����Y_��V��k�RL�>��1,���{ԭl�
�%EU��'�unS��7/E��6r����o[�p����Dƚ���n�� ���#ښ���Y{
��G�� 7\@جE���SA�p����!����Ԕ,>qN��=+r��D�Tf� �)W�`��ԋĆ��9����za�G�mQ'"�L#��ȫjǤo�G}��p�uW�!1�	UoN�Y�2�E��<x�� ���&������h��wdE�IE�/�Yo4�T�2�?�M�f�(�m;���^7\5�GqLyB�`yO�B�$�	��N�>�V�>���W��ir-��(>�{�w[�:�Ѱ��8g��;y@� M'!�N7�f�Q|d�P�_w�;���X%k�c���	�ߜ�oېa��`��)�!�[���2�Ob^S2C���h�s���NViB��&�h��)꫍���aߝ�۳U�	�&>�@䑜 �3���]rbƩg��,�|���׆2����r������YQ�77tT��設:��]/���@��E�Er>t�� �G�
�"U�aKu:vc�#�p�ק�|DfS�#U+�>�P+��pO#���w+���~��@������������9���-Z
$��_&a<O��{^+Ι�KIiɊ7�b�ͯ�*��PtH�
���o���҄�b\d$jO�M� ;9�����=p�C!����1"��i�`Do��P73%:�=$�:>��v�;0��I�h�uG�zʦ�U<�;>ղ,v�i��B��q���<�7�7b���K�j�D`�k,}7QqM�h�
��v��s�;�K��`�;���$����rϻT�MX�|�B�cc�j��$�!>BQh%�Ǫ��1�_��6�[���Vt����k�D��Ǉ�.Ó��m
�:����:+�� y�������u�ӣ��;Ħ߃����F���U,C��R���'8\.��f�2j�W�K!��ޠM�~I���0��HIj	 ���iP$c���܂-F.�YyVERJ�FiG1
��`���,y.��>krx5�\�jө��S�c~�n�픥��>θV� T�ۛ��X��h����$����l(bF��~�6�b���$�=lQ��Cd�hi��Z_�y�,w� �c ���
̤��������J['iC��.H/�om6Z7&4�1q�ƽ�d�2�.��׳�Z�pڅ���5e��"��>���(m�)�v�g��9O�Q{� ������Sߞ?wմ��o�MP���k�dY�U�,Lfk���ڎ�`��w�kۘ�X�K$K��m��<E�fk �D:��R]K�\Y�Y�+�w�!�z��MOK�A��x��ԧ#�]h�# F��C9w�Ҵ�E	�©�#1"�5�fi�zT�N:���>�y�@U�Ĩ��94m�O�2�z�^�MKT���� �I4m��=�!JI�nt�j�2l�9:D~���~Ld�T���_l�Bl�`{C�<~{���q��!�3Q��@��}8dګ�[8J��m�p���p���.��2�"T@'���$����h�#0����V���!�g��� �:D�i�[.�\l	T֮�r-��?5����P�Kݚ~�^M���当��2�����u��X:�� 9�0�*� 5d�����MT��{��:x�$����{je�XOv��鞾�ɓxNĽ~��	�˳�b��5/r����y�F�ǹ7&�t
</5�⣲�Rr�>�}U|��j=�cf� |��j�X�W�+N�7����D�CW���.u�j%��x)vE!3�6�p�ת%�a`��o�,F;,rd˜��&�e]	Ql I��V�6�My�2=y�72փ$w�q��}Ȯ+�`�����m�a�E��8�eF�+qc�Ul%�ᡚ�* "����,K��W�*���cHܿ�����
DICI��+cD���HM�/_o�]��xp�v��_��F�bQW�@��VU��_d`e��W�w�=ۖv�����P���
�7H�:c�)��k��Veu-�;�m��.��F>�{�5���@@\�kօ@S��e�seu�1"�Su2�k)8��"A斀�:pd�"Wk=��,r5yuR$�q���\�[0ÃS� ���y���Y� �{�|
��b7끢 O��(�M��.�������� ^;�מ�[��?���;-��\�M}��c �̚�mΊ��2b`|�B�\�䄰kz�O���aq��㛭`0
��O�����J�����*��Hdҝ��R���7������KLd���b�9jS�H��&B�y!^���ڂ`�^�8�6*��Eܿ�1P���.Cg���Hl͖�L%Č��F$����gEjz/�)p� f�I���(��z��`��<! �0�$��1 Ðv�M���%�ěU]�3:{�bl�f��9jG3�j���oUa0i���3��v��#�Ȳ�㣙9�t��W�J�������G� ��c��8���}_�4��p�3�	�(H��z7y���U�'&��S�C'�?��@d���.M��K���P(O�"�Q���0
 a�����t�rS��%�m��^� �d�������@j�{�����_�k%Gpțo7n(��i:�JF��/��q�r�[+L!O�6���Ԙ��o�JJ�қ�uIH�FS��j�<%� �Q����_n}Tľ�3-
2Ã�/�V���oE��4��,����"����m��x5hX��*C���$雏Z߮-�J&-�7;mX_��l�gt���ѧ���A��u��i�2�������-�sEr�� ^.$���G�9Bў}n&ɓ�A�ab��i�U��$s]:�QJ��"B�c
f�E�6r~5�g�w�]���( #}j^�p�L �J�lV�%��?ͬ�py�T�꫇�n��;��
��^)1������=9���冀Ұ�t+\O�AyDk���I��\�K���3,R�#���z1qE��Yf��1���@�[k&��U��<�ȉ�0�*��|V�G���3d�M��,S��?n���1�8	t��]Ǳ���;ٻ�:=�$=F�����p���U��K�?�����m������N�Ќ�%�LC#�G`��X_���b����n�yW	��[{[��K��$5�,X���	NIH�]��E��K�'���dj$>��]���Q�==&y�����R1qbA0>��!5H����)�I��SjJ�q%���M��≽�W���r�c}X����3d���@4�r��̠��(֗V�![	���B�RoW�Ѓz�'H��z����P~AВ�h+�'��č�� q��6���}�|*�3���Oz9(-`�ǄM����(�69h��O���r�ⵕ�nr���a�@E�2?�]�O2Bx���u2��z�VM8l�"�>���/u_��U�Fá?%&`N��f��'�W	iH@l^k��G�D��k}b['ӭ�0D�.�|�ay�P@m
�����څ�L�e@�sy^v�����,&���4�`m�
l-c���!Y|��E�]���G_d�7C[}�yN�-:�k��HjU��{�D\�,Fۀ��b�%�0Z����M��?��^o���-�F	!���ɶ��ک߉�͈��w迃{�'�4~����1��Iע��g��ǋ��E!��hi�߳(uE=�~��䨲L�;]��B�E��.�1PU������݇ �'��7��	7�Ŋ{]�sl�/T���ó^n?�|����{����,�FR�>�+���V��DT!Y:�y)8(ђھE��3��.��.<�S��F��7��+�k�zN��u��5U�iLDz�5��d?8I����V[�U�"�5�#W��
k3 R.{ū(���j�<�:�3���l6ܔo���d�.����G���@�N�GRRd)J�E�Zz0;n��>߉8����kG�����L㽏S��Ƥy�e�d�g��}Hq!n����,ya�K]M���Q.�ǹ�c��E3 X����}��t�PX�X��2���M���yZ�fݨ�r'�Q���W9Tz��7�-Q��m��9�r�����uN��G�����{eYo7]r��r��X�t��o�t��2��8�CҶ���빢r$ڣ�����j.�R0�ă�d�#8[�� �u�Oc��t����a�s[H4`���+@��i���v��~���sw��]���������e���oXܗ��K�(ɏ�3�jV��qz��|`��,�֫a�k�C�r�T�v��H.&�7@�L�R'�UF� L#.!��������|�v��)�Nԛ��]�3�8ֳ��+����5�3h����(_)S'b�i@%��cL�(�?ns;"vEN��2;Z �Ɋh�b�Ӏ��-Yk^~2�W���QwI �~�6�Ҷ>� G z/e��I{�U�Rs�j���\��bg_ �F\�>��-)a�B�)%MI���PPa�,����i���M��p�^�6���{���w�ePn.�o�q���=^��cr�T����4eG�!��a�9���U@FV���>	�"���Aɭ�	���H�3ch���јOu�S�W��v�9��R��p{X �X�]���#�?E�(y���j�x����0���%�(��ָCI�i��g1��x�;6JA��h��?wi������O 6��Q�qe�-��־IM�� �D�Aۿ�*�x�.��K,���;s�W�U�	��f�H�Ɗ�z�O@�I�v`�n�[�'�k�چ�x&�?����k�t�/�f#&E�A��<Is�y:F WM�,o+�.�)��A؞nS������QA�ƹ�]����|%[Nd*E�}��3��S���qR�� 9i���5�|�!,����Y�%�Q�QȀ*-�!�S�jb[�W!��ϴ&�+�ވ'W1'��#gԨ;S�a(:R�ʶ��A�|�9��<�QJ�cW�=B�Ү`�S�[W���tXiFA՜G��&V���L��L��)cM�FF���U9���!ˁ���mT��/o��Y����L���{�f�u�뽄��5���x[Tt-B%v�j���)WGX�֕����̷�'$�>&���w�<X�2����Cl�|� � \V\�h�L��k�
�4K��{�ho�$�<����?Z�+.�g_����=9���y@p�s�6�^9�J}�"M��p,���Bn�p��E�.  z��ʚ�#�Ɛ�o9c�C�R��}�K�|5G�?��w4�clE;��J��Ja;�h�!\���'��1ه%����D���uY7;x֥����s��:2�S�����Ն�q}B�e�KYG�Z�x��M���g��H��ʀ%M�=X��G��`o�$��gCU�`d���1��Ԟf�!:��,�Xj�]��9��g{K-{d�Q��R8�\L�$�E��h*i��ʬ���e H"�F��G`��r�6�L���hOc���XvL��_>07�^�֘z�_SE���]�L�Z/�T��Gn#@C�x���̓�{��=N>]��`)2
�?��]���,G��(�qd2����1��,1��	��a1A��-(��Ϣ�������!�tiM_�d�`�y�<�b{W���*K�	C��;��ۣ��N�n�~&�F����v4V?�l�����;|�$8`kf�;�؈j��7�s�+a-Ē��ď߆��'��ﳀ4t6aK\���5��gn\!�҄@�R$��B��;�P}��}�4O*��T[4�$�bBD�0�<�3G���4��!y��E��]���e9ؤ���{Y���>S��"��V�cԒZMxi��٠�R�Ws��Q�`)��Q��u������Pb�}
pm(�� ��y��$�ګA��#�=�����\� a��Ft-�ùw��j�X�e����I9.����l�}��a�2�T+�U�$Rs��`xD�m���9^���E��+���x��=
8�:�����5����7���f3_��|�y�ǘ�ۿ�!���MMRg��:�ö�vA'���!s�I�����t%������hMd�
r&6�"��ֿ������#%VxR޹ao>Ǭӂ��y�6j�V���%v&��t������Rm�u5��K����jR�%@˄���W�P�D*��Dw^�]Gm^"i7���l8�H�]	�+S�>�ۗ=߄y�R�{ø Aքܨt+{�;p�̜��r*�*�j�C��l��ci�6���gR+��36<�_��8�,s�	��Y Ό�$G�3X�Q_O*�0�x"������q@'߂�q��l��{J~yu�M
h ��_��M�K2g�d��ߩ�CȮa�Q�r��W�m/�g:=ȍ檩Q,���Ds��af[4���.FT�&*�E}��Q%U]�#����6c �Kw�CB)�g�?~N8S�Fߤ�S�]\��u��sLq'fh���k�i#XAq�j��$��N�J��ǕØ���¬~����^��)��8�u`H	G���8Pp�d쬜&��=*$��܆J^"��nӄ6H]O��6���> ��/u� S�9?�6i�)�Q^
%�zǩ��>0�=�{!q'�n�C��Wǣ���`8of�}����=�EHƾ	wX������a�&j�ć`PI	�"��$$�IUF?�\��5J��RPh4��M���,h^�<�EM+@n��B^�)��F�ʋG��Z'(Z����@�:�����C�z6�C��;XHʖ�L{��'��2GY欏������:I�n�a��ᳲ#z���8o\?S�b�~�'�&�h� ���>X�k�jc�6�,��@U���̸�<R�����*k� ����O$+�*�1���ig+�v�X��,�JK���$L�P'�h����y��x��!��'q-�H�|6���bk����R�s�o�H$h�Ywd'i�zp	��耈��&s^X���5�f�t熇�Y��WOy�J2��6�ϴ��Ղ�O���r<"I.�P�+'��$� ө2e�\4گ�N�)��{o3���;<�4�!��/����u
(���І3��ֳ~���$zu�Jl���c�	�v@�I�0���)�7c<�zLG}�d�3_���y�ʼ���W�l� �y#̏%�Q#�y>B��F.ڟ3=��\�'TU�ʔnl)q�v�O�3��*j1q��Z=�+JxN�7(�2j��k��Ş�n@�8���I�A(�Oٿ�e���2<	���nV]|����R����<�}��
W$��41Y�X��	��A�8��>A�BU�3���ꃤoT����Y�ָP��K{G)~�u�8���5���D����� ����bԉ���"�+�9.|�D{*a$�
�.w��fN��E/��V��hB��U�*�퐻�i�&���2q[� �Q��G��{\���j��cȮa`�����K��:�"����>"}�H���G�N���t7�S�5FoY%�8��������'�hT�߬Ǒ���G����k���v��$����q�O���(�4ء��R�J��O�|]W���T�k�f"g�(��[�'������>�dgv��u>8(i��0��Ab��_oЃ�l�� �5-��x��.������J�r+&�h�$��D�(���޵�"%E](m����C�s����j�_Y���ivb���������s�dХ�k�Cv��?�y&���Shc���ŀԽ[~�\�m l��>7���:��:�УA���Pzފ�FP���Ĕ����v�Q%����D0O��{DBih�#����2R^l�e]3coH6N��
��|�>��g��8\�T���T�?@8��$O׍5�$,u��`��%��{uk�����:�F��d��[1_�{VG<޴[WH;Ӗ�73w�.B�7ւP
=�A�h �Q}r��K�O"�+���)��ݹ�9h��!�-y��KS���u:v�Zf��wCaeB�1D�͔�қa�Xk��f	�G;����X�m�l��7�I��'����eS�U��$�w;.��ʶJ�@���J������F��omfc��n+R��rD�4"XL�����T�"P��8��q6�ry�����J�M�Н!�x�)�咕1Kf�t&'��4�?��	�ğ.ż���}�[���|��s$���'(E�K�}JH�{sO��y.U�W���`/��O匭��ѡ훝�T��ϡ���Л�7����;�ηĤ�h�m �xɶ����@�R�p������s�F�xN��lD*�>Nsl�>9��߈&��䷬�Z+'"�Pk�d{/ވ!���p͉�[q�wr{@�S<HK�E��m��;�k jã-��=pO�^p�pz�߅�W������ ��!KCѠ�ln��i(:��D��2�F^qІ�d�3�~,/M�?"�׊3%	���*ڻ8�Z]��1�0R�ZH��:J���i���[,/����'���ڮ�Lgt��Sn_�~���G�d>I�f8�%_�u�L�0�@h+eI��\0���:�+]��S]�)8�+5���B��.�1^qD1����μ3�%Ճ��SF��*�;���l~Y�S�xI�}���A&�f��d�vlм���<