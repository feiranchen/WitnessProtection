��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*���o�!��=e��O�	BIλ������sI4l��N��z~��������bW���v^���Z<R\=r�R�(�Ԩ��i*�VD7��A�����#0ٴg{��]��z�Rx� >��%[�Q���J�&��u7W��7��LP�NΏ����Y��D ֤˗�2����3WX�"�V[Ĕ��|��0g ~ ��?%�9�B̫��TY�q�eybz��&���*ʢ9|a���*���{5fdXj>�56t�Yrj�L�O����
�Ak^�描���>`SˠQ����N��ǽ��<P7�]2�nȆ6��m�� ��}IQ"�j�( �~\D�N�TQl���R`�.���i#{��KW&��q�CS��	J\��̙є�Ņ��]�[���&�&	�5�D�r��=rg����t���iM� ��|��dS���,&�����OK�Mą޵
�#	��p6�8�����U�ل���8�(c�C���O�H�����XUbg�nT���/�z���$*�Ǜp�훙h0f�?>���Q�D��\��)�����Bu�[e���L�ҽk�;��Ȧۈ�m�}���g�f�_Z�,:>aK	T0��*V�Xd��̨o���| �g���%/2�g��"��]�㖱�z^��	w:1��j!լ_�JPΑ�A���
g�S�L��#_�3�<��Y�˨��D�:7`� A���g�O�9
ƘN���V9n��(���[$�D
U~���{u�����lk���$���A/�hCK5�W�����H&Xrm*h��+�<�~�m�s�(;؃5L�ӽE]�����n�N�R���p�����D�o�h���(.�Ć�Y�L��<@���H�}�����fJ+��,�	-�%�%�vjڗ����jq��M�2h�L��i'��w8h���{�`�~�O�=C�>�o��h�Qb��7'@�%�a2�E��	�yW�`0�D��'��=�
������	����V�1˿1ě��۟o�.��@
�D�Se�+��ɲ7XLOvv�>ƺBUB�cn���p/��3����#�DֶPgd�kv9�9m��/�V��Kb!��l���.έ�+�˭����n��2��N�����W~���Ĳ�˃'��}�|55o'ѮF��w<��̿�@E�Gc7�{�c�]ƾ����)����7�u�d��%��	��\S�EW�R�+�䵉n�ɲ��iҖ�%U��װ8Y��+:/�mn\�Uv�{鿚�S�n�U�
��Wb��p ��H��g*�RU���%.l�X��5%����FR��݂�I�"�{���8?�K�P� G���,�f�#R���ȷכ�)�������|M4���������lT�	�,�Mb�Z���1e��f�Agv��=0-_��d"��+O��\���L�jr60t�.[ɩ�ҡ�;�6�M[x�H��`�p�1��6敇����8$fz([c���f�}�� p�F����d?��9�v����P�E������3b;��Hrj��L��A�=�B�1�.�x��˨����	��S�$GI����~�N"YZ��4�"k���y�9��Z�(���e����P؁ߓ�y������D�W��u($�$�{����r���
���[�'d�RݎA��5�Uڀ����q�]�[�k��v��Ձ�t��|�I�O�#s����Y���l+X�G0]���ςfv��O�;�1���?�
�_N��T�꫌�Ś��6�Z ��BF�3����k�X���H%�	kf�D��kKr�W���I�}$yqH�7���S��ط�jC�{u]V�ɱwyh���n�����uh�R���{��� ����o[`�����u��(s6�������ӎ�v8��v[�F �~T�'�<R��D���^B�	��B��&w�NVv�]D�1 ���r�$�Iѐʔ����
3[S��`��O(�bc�6p�՚y2���.H`_�� �ܫH�A�����4��%�_-+��hP�ﰧ�
A�M��&ݛ�����)��6j�L����8��<Q��P�40��.U'.p��EA�I����;��(�@��6Xu���|���3�`m��5�Iys��  �#�1�#�4�T���'	�����35�(o�.9�rH�r1-P��|��5X��j6ѸjQPFq��c�|uY�PF��7� v���ZC��Y�Ek9"�1-OF��9�4~��Xi��SL���5`DcQ�[��N�e���{�AE�R��B�^.aV>Lqރ��"1ƥ�����X69��zE�	�U#�<!��+�y?��:W'�sx������ P�f��tD'�dxQ {ƿe2�{1ֈ�ǂ-+�z�A5z�Z#W�BP��W2�tߡz��T>�ڎ�F �G}RD���IpH���V??��S��"�3�Ν�oD�g��0��n뱾�yb���S�$��W���wt�!7pqpm��*���;q5l�OvN�cB^k7O<�R�w�fH�3�w����k�R2-Z!��Vhr�e�¬�Y9A��W��P�~��]��Do@�.��x����\���&�~6C@�1�pH���*��!�p�`�-`�`��%e<�$�s�0a r�`��a(�9�I�8LIB!I��	*c.B9��7�w��}�2J�ߝ�h��Q����ٵ��2����wp��f_�BfG��RY֘�e����+����vպ����2Z������ɑs;ܭ��q�v��y(GD�P&�н{z�΅ovc���&�ŃښWި
�<���Xc@%�74 Y���~������{Y��i�1�i�r��ytyE v4���m���1�����b��?�n6�9d=�z�z��!�%-@��D��-�\}w���HS��f�/:����:&�F�!�Mi�=��y�,P��y����X�U��qSIJ����be�;��?��*1����'��o_��3�ÛK�4��#)p7�,Bɿ�	_RV����6�;���R�Ǻ5ƭ��U�il�r� �U����`��n�x�$�20,;�u�[��t�O�h?ݝ�R$�dI*� J\�<��u�/r���M���KVJ������V-�%A��x>���� ^�ÄD�D�i-^��l5=�ޥ��JՃ�+���Z�X���Z|�
s��	s�o.� r3������ωQԠf�ms���.�=���]��$����Z.�7m�cu
@���ì�����m�@���:��1����Y�$!0 ����|����h�k��)��N����8aG�ϼ�h�>k_z�)���H��5b.h�Ƨ�9?�F#�0c��öY(�$��^V;���p����fh,�����6�V_�����&��Vl��PU�3�}��D�A/�P����ӫي��26v��z��$�)b��[4pؘ1�93L#�
��j[��d̬iB�^�A�±��I���N�� ��F�A���eĠ�g^E%�� w�a�����]�,��I���a��8M�X�-�@���G����D���G_�3�`�'�a.Z���<�lf�&��J�)�3�P
~�/����`Mp_I� �e���l��KgI�)���T����.\i��d��F{<x~�$i����:5V"|��v�Z��=�08��0&.k߰�
���KY#�[����Q�&�F�|&��,� u]�7["��au{�?�R�F*B�g6ŉ{9�K��Aq	T�X\��A�l*��n��t�%�ԇ#��d̶A�wa�HL0u��!^�h��-jtLK����͊3�x(�bq�+:��Q��Q/�]N*�*W�Q���6�GIMD���G��w�N����[�bo���$���������6;e��@���ݑ������X��]24�ZM�.�bZCw������BA/��$D+B�Lw�RD��nqL�Y^X���K�LhJ������+��F�KA�>/o��Ί	�4�Jjc��A���[Bw=M�Ŋ�WoL��ϰ ��d\�Jk���'FU��B,�7�?�K�������Nu��r��xZlۂG1�R�P (��*� �/�o�Д=��Ǘ��d�kb��7.�i�ê�j>J�
�� ��W�MY�>�݄H������7*��A����Wð"՛�8����%]F�Nu����3i�%�_�K���Y0��8����W_ȸ}��
���.lۘ��g^ȿK+�Ύ�@6AbJ�w�4��M�������[<���P��FVn �|N��F�H)�Ă�<�|2U*�A�o�NY�ɳ�jؕ���%@�c�T���H(��yc��m	�!�T�躊�Q�r��`�_w5��C�ٻ$�3:��+��X�72n��H�u-�,V'ʓ���s��u�[ԘϽ=��XR�A��n���v�vU{z��6�T>� f{k����!����'��0_3<�`�T�����DK�X��+�'?kP�o)�u'�a2;����X�]n�.O�O�`1�-��Mkع��;���;7�	���h�P�܅�N�҂Ȯ^?x��<��_-σ�&�^ƀ^�xK3�|��7 R���J�˪eg�"�0����>Jk���.y]�E,�l1Z �=�F�i�-���TC�&y�Z�&��0�,�
��	3�y>�1���'��ƪ��g�?DF�I�C�,��"�Mly�݈ҁ�1��_�Qa�-Y��%�7�/��(���5/��[����f,����%}}���F�W�Xp7�����%3Sݠo�9���D�`���@@�����{�����13'����@�x��[=sBRfk��Q�EGs5�B��xֈfVcAkjc&�{fvO�b������N�������1-��&-yE[�b�cI̢Q}@��P�E=������Y��L��Ih˔y���l|��q����9�If�@�7L0��$��.ԉ��O���OC��ާtP���:��Lı�|����Փ��B�I���Ѱ�w�w��Ű�F";��Oz̄	�O{��tƅ/���R�Lբd�N���B��^~�ӈ�L*��/8b�e7˕��ô����uCQ�Y��*�)��u;=��9seI���F�>'��i���Vw.#�|�����8;����jɈY����95�P&H��ߘԂ昣�"<=�w����԰)X�c�^0��Z�p����a��8YХ��:�<Ы��;��z�4�*f�>��G���v��s�&|���GP��(�kC��/�5���m�a챶����cT\!P���,gD��-΁, ���T"�9q�G�����z��'��@f��D?Vyxڝ�5ɀ�@lRa���A1N�1�����?ZD�L�z��_������1!�ݍQ�V�S�uB ����$<�JoW��kC�6�!-����Լ��.#x�V��A�pbfv�'@����X#�\��G�����>�
b�TK�����U��2.�Z�㒊G�.Dʇb�Ÿ����A2x�xE�ȱ�y52�p�<��]���s���%����W�e���7�̔ݟʘk��$�;���1��52�e}?�KRų�O$O��x����>\M�̚l��l̹��+	Fsp�}ǲ`,��^K��\����{�ձ v��!���JB�Шz�"���p��/�)+�MFK���-찒V@N��Sg��d�eF(}3���߹��,Q���M2G�"vel0�[/K�3!�ˇ�h-+�k�8�8�:I��rz��n�@���.`����H�M�Ԙ��)/<v&bp$Ê�b���%�ݟٹQ�'|`���;ՠZ�ыG�|�3�|1��a݈b�)���?ֶ�uM��X٤������0@�bR�)?����u����|t)�mU�Ѱ컐~�o%��}9e�ِ�B���B7YuH�& �em��	�D.�Վ�MX�F�s��U�Ԃ.zO���v�-,�o�q0��=O��!+ba����зI�Y��y.�K@:��p�����g�WfզHx���i#��佂��x���W��:��s@LB��u�� ;�+���WB1��z���޵�s���W�u���Q�}�i`�LG+�q=9�A����vl�t��~g���g2a���'�h]rt.?K�w�����(����+f���*�__��G\(ACMzu�{���J�5B~>'�Ʊ̓���d�N L�Х�x�.D2�I_�e��c���酒��:� ��П���膥�{�.M�n	R�Bj�2lז�m�ݳ����5?�� ��g�>��D���ӓ~c�鸤����3Y����-��:*�4*�cJ*.�_�"�9�>攁��I�]V�Q%��P�Emy^w���Ė��\B��̑\PW���=�[C;@�*q�AUN������~����Z"�Q		>���T��aO�y?$�A����3�%��C��ΖćX΍9�bzo�Vz����'�)H8�\�N9����;��@h��G$���b�	r��%i�\I2����0�Hq+"�]Z̿����A�r��P�"�QjӒ��O��s'���b�RdGu��J��q����"�jlS|��&�i���ۖ��#�k<ǉf@34�(x�z8�J�U ����A�Rb)���M���7a�d-���v����o�����BB��cG?ȝRq,F}L���.��!?g��.�6g�����e��gLtP�1d�&�H?k�ް�VH(j�	0�ÛP�߮�J�1���j-�"yސ���v�zl�G�*<@�%W1Di�thF0(�U�M��S 8��A�	M�]c8`�Ud.��E�d>|C�h�n��ݎN@���"��c4�ůr����*��_~e����"?����y��<��9��&�S�m��)�
R�1�������zƯ.���� k��It�i��	�۹J��Ek����Ν�F�y]�P��ӏu\�hFiڦ{���{��{^�t_6ER){��,�r�9�Ŷ�꽑��M�Vrs<@��L�p1o��ƻ�'���Ȼ��#��ODAA�X�LE��b$L[�r+o%霪��Fa�
���H-=o�H�1��ު�5�Y3 �$����߷rE�VJ����O��!J���ׅ�g^����A���:���Ocf
y�����ʇ�1���;���%��w�,,^D�����.����� �[Z��pb�$�g9��m`c���9\�]�g��`���u��|���I�ϕR��>[.�*����������Be�	o40��}ɰ�̼��F��߷1x��ui��:gK�+�+b'*���خ��}��Qx���ؙ㊴Ec����R�}��)�d�vynFN�ތ?�YQl����Di��}u�%�d�"fn�8Y|o����}w,��T���}pB���-��D1!�-���c̬ĎA,ɣ���჻1�e�^Q�]Y_�<���}����2�^��3���c��-F����pxl���Qnh�n �8>��Mf����/<*n7PJ���@���I|��y��WQ� ��A웲j�=�t5���8,��֑�뜁b��	���j	���am ��7+�x�dq��i,9|X��3�k���h]�D&��ܻ
�Ø�~[z��SD���t��i�e�Qi9X�>����״)�u����5��^��ya��;'u2b 	��:�雤p\��!��ޏA��P�ّ��$dP��d�*:ω���Z������F���b��9�JG�P��'q!h���EU��/愳�=���ГS�;�g��Z�M�$B2��R�P��tXs?9xI�5�7~�슫���Q����&q��h'w�k�0��>�|{�L@�/��Z|"�xO�yE+��e�sz��_�f-k��}`W�m�����|�ev��E�"m4Y�(iÈ@f譎;�����Sc��q�g,�	��f�'���?�sWEYCW޼$G�3X}���kP3�3��9�H�����Ԝp��Ԡ�ѭ��8I.�O�*����%s��xDgr�kj5ƨBq��Pz��4��&G�)�y���PhmP�W�8ӭ(��!�n�ޘ�r6��w�o�����+�O�n�T^�T����s�͠�	Is,�5��7�
`����$�y�	��[C*zM�|�`r&�%ivp���"�R�Ȱ.` z�x�[�e>���{*�!Z�JѦ6'�9p{k4����f_�y�_�֙k�C�5���9��~��N��[�pԅ�:�o��EyWT|�Wڻh�������7�T8�G�V�S�?qv�r�=R��u2"b1�Ej�OiaDSN7���p��0����: 
G�Y.q��kX���Z��ƀ��&�&Z!�g����w��i0lҞu���/�э�� k%�T� 8['�<�}��m�=�L�»�4�D/��`L��̐O��]/�����;� ����_���NW���b3)���ރʫ�!���`���w���zW��]��d�����r�ޥ��)珡��s���Ш�l4:�L)�&��b��g�UP���<D��1��N ���.�!�@;�{֯[Ѻލ��2)�a�(�R�K�2�3(CT<���n纖�@�9��9�ojP��0������t'�HiUy�"E%����	v������Z���;��@�onߩ@���dOQ&�;�i�y1AGkoZ!Te��SO�:!
�{��{&�C@�C+&���rs���XƔ2NyM�Pa*���^���&�pBŧ=��'k����!�f�.�_�����v�+V�_�%����mW��U��8��T�L�W)3 �/��5�����!�����#��0 M|y���Pڅ��i����	�ӝpryf����O����T���=�O�V��y��7�U�L=Q�lz�[y�dK��o} 6�XY����.}�����I������E?���C
@��}�`"!F?y�c\�ߣ��#�a��<�@?�ѽHZ�@��Z*�O� �@�0��@�/{"��y�T(3�������Tغy̅o��j� Q�b�%��;�6��ׄg�/��s]e2���NMU���#�x%!t�/��bJY
�O��8���J�=N[�����պ`��?h`�ĲoN����`*�S����b�a��|�����Nr�)d�?���;y�>f�:�B��ο�X�-DlNSÇ����� ("��8�k���i�{r���i��n?W�s�CeSa�M���rW��7e>��!�3��)�f��^��U��̂�/Ôjxh��!`؞���H�
w"Atʏ���'���:Bm`�.��͉0&@�O�Mt�k�'���~�O5������� ��
<�*��¨�؀��cjg|�1i�pp������P��
��V��wK�^�$4���X�G-���T1`̟�i]4a�D�N�Ŗu]���]u�p��6�n	>�N�m�buʻ��A�_�k3V�M�Tk���08VE��o,�����P�����g����È�IH�Tr-8���Ƭ;~�;�qu7e��&x�5O�� #��)�ܔ�
/������򭲫WC����Tq5���X������ Юx?7��ګ���A�/׮3���>@&�Yeia�2k��/ɂ�*"�{bD2lvh�)��.!#w��~7e�"s�� ߯�YC�X��;C*�$���h����F̡W[�������(8��r:��/�͕pE5������_�GS���?%������| ���O�����c-?�w،����V�uʬl�\A�	��:�(�`��([!I	HdVc�U˂���'a!��v��G�r�9BYr�E)�d�_����hK.��P1h��] B��ﲋ4\G��?'��:2��2ς�-w�l[Gt�J(Yk��׵�f�]Y���w��mW$[r�C�앖��A[]v���� �6�L9%���>5��I�b���lBx��� �c%LZ1_Y����5O��cL�q}R�:aE51�����yVU��Gg���\���U	�0�9��۸�����Ǵ�MZ���ԅN�������-�Qj9oi�Us+Gr�dX�l��������3��Z<j�]���G����<lE!g�W��Zy/�х�v��&��} /=�-��Y7{1�K�7ʶ�{��x��LP F��d�Em���/�b��1+�4`�X��� /���_7k �/o�3��/��"01�d���ϻ+���\��SWU��dy���(̨9VH��Py���lo����n�Nֆ��fRMqW���{��Q��ы�����j"�YT���`r�p�b�o��/d�Z�������2n�����XnD�N�������xC܌��uﱹ��G@	�dsy��v�+�+ *E'��:���Fl-�N=I��R�0���+Z;q�)�Ϝ_�� ��1r־�Y�=?-��M6CN�Ϋ�}`c�Z�����g5?%g��;?�g p����z�@m_���f���TYV�]�g�-Ó]��ZFGU3I� ���%:�_��N/�3�<<�e�*$)�(�˺F������0�H$��K�ZX�1b��l6����Wl����{�|4�%l���>�h�sd-��3	�K��E��N�#lZy-Ǡ�vJ�J������}v����B��,���#'��8���s��;n��;6�S(Y�?S�ZYɥ���9����,����(���^��p�(a�l��'k��PԱ�$����u0���G��`-�O����]���'�&r����N +x��Rl���`���9K���Yx��T_��gO|u��؀��@�������l������m5UF���l��VR��X��M���AȃO� �������i2e��Ep�lg�o������4�7���	�!Rgs�jT�\6<��$�n�@��f����o��~-��h���D	q��W��fͨ�K���`����~{#�@<��t�����/2�+x�_�V�)��ܭv�v����BF��qs@z�3����,O9j����e$����l�i����o�ZyOd��J�d�*�F�V�QnϽU�L��*Z<���;��Pr�N���D2}2���RG�  �um�&��ac�Y�1s܁����b�j^�h���^��?�}*~K2�
4�]X"O��
<�-)��	YX��E�ȩ�d΋�^��yAC]f9#'��v���}��U|�͒]d�2'��9���wN��.�z<\�z @�ȿ�I Ʋi���v��ݗ$ �
?a���?f�h�jYkTwD���Uw��{���\~��0����`������J����(�*��)��a�zgTG�Ͼ�O�nҭ�0�f	yYY��e�@0���1\.�{��vm��}U��S\��bh��|i�>��7	ŝd� ������ P:�i�0�R���j�οc�^�We���:eT�{A�C�, �w�`G�^��gV�)L~�ڀ���c�MFБ��Gt���e�g��cu�����UP�	3`���R<�5���u�;XPp��z�\���y�����@V7��I�u���ռ�m�4�Ve���[z���a`�'���L=ΰ'��(g�w@��n/A�n��J.�<��0�*�c�s��֦���-q���ￓ���;ͻٷ�����{�|����,�����)�ހ���	j6�h/W�[�v���it�v�`B/�deo�@��g@}zR�j�y�ظBPR%���ZE"_���*����8<r�%�����9cX��"b>�\E�ūh�ʵ	�[��Sj�b��	I��8�O?��q��,����]��0O���v�:C�M�`�&�<A��\��,WN@�S_��UMD�6���^�2/�ͳJN����.B���!�U��&v[6=�Z�N�9�7���6��U����PL;5N��YHxPc�?�ι�Rᨽ*/��P%t���� �G< aѮ�K_2�Η7�̫uŃ�lf���kUm9����u�d��7�m]V�J 4�*	�Y���m��!E�2n'�b�c��D/���΢�'�Q�=3��o�ޑ@�F!��t�ӏUPA����o��'e�vH�Ⱦ*�������> ���VV*�'�����L�v\J@ �[iY7e}�P����3�3C��w:R��,�F�d�SDV23z���j���]�:9�x��O�H��+�?�t$�L���8�W������[����Slz[�ُ��~���,��j�,$s����E3-���H��~">���i�����ˍIAS�:)�����0�G,L*���D'v����o�gZ�{t������Kǭ�=�]���2G�!��b��d3�$5h�ػ���R�$Z���v�B�?Z�\`U����-�j�@�w_�φr.;c 09�I���A��m�l�����Z����{�d n��>�3~�d!fwگ��_}�� �[ʂ�}�>����3��x�+����zSD�-[�}�p.�R��5��./�9X���/�v����x�����C��U�mX��ʽ� ���� :
���l����n�7[^ñuzW%^�b�E�;�6}쵢�����xV�����h�#���[��)7�bU� �J$m�u�����L���n#D���� �,�&�c|s�}�T=��u�����2��{�AЅ������!��\��G.|6G�{���C�_J,V��	��1�{�n�ѹ�=����4����{�&��t�{��vf���:Ϳ�5�����`Xx$�7������6�jvnz�uŚ��ꐇ�\�\�DM;��3�����q��d\2@�e�x�{LI��=��$����K��Rf�'���=1�]f?���!v���w~z+':���y���(�Cl�q��w!��L�뜿^��//�VcW�fZ�;=AL�i2f�Z���X4�[���J�p��F��f)�[�a����n��W;.�&4�I��s��ڶG�-�kmh��ńN�xrh��&�aj'����B�Y ã,�6��r�=��|}�R���d�j���o��M���M�/\�0�9U�pC4�MJ�L�.:P���9��6f/�|C�C��0�+]��	"�k��S��C��lifW5�i	.��T�X�"L�>~zY{v�ź�I��w�Ȁ� �Ro�M~"�m�4��&��&x����~���Π�̑�d��v�ѿk�.!�!�S�by�H������:ߋ�1��O/��Qa�c}lgPT���ט��a�gU�8��=�(��x0ak���{����_�V�U:v¿����kQUeo���6wS1�t�*LI�ҡ)&?�Uҏ��ʐ�x�!n�{��;9[1��LBYcH�x�5D�8��y�"��_�nY"��Qq���GSEБ�o����bTLkAc�:V͘� �?�Oi�*�=|�pYF���c<�'/����R�������^�5p̯
���,ԁdɣ%B������ad% ����� ��o�Z��Fo��Ii�?����h&q�����cD���.RZg����cO���^�)�b	M�ak'C��ͳ�䈳��H�WCC�>~w-`��n:9�b�e�ӊ��f�S���tre(�!�B>��_�yp 8nϏ��.vX��~��t0�z,�@�,+�l�7�iQ�7Ә䨽�7[pdǈ���fW��s�O[��9C�p+<�����r����ۊ�sV}��V6�;<���Չ�k?��/���;�Y��*6u�{p�����y���a��R58��d@������gՔ�������͠�����Ԇ�[�L�����@k�)�=�IF��l��e|��/0�Q������߼B�?�ů�̚�q��yC�J�4���4ʡB�PmC������j&*?5�t�?��PޘDwJlΦ<�W�.�t���.I`�E�R����ɵn$w��Yh8O9����� ��;FN"e�(e�
a���X�����-�t�n��k�i��~�FsV�Nk�.3���7�E���!�ݳ8���P�X�Y���ᄷzy��T�3��׺�1�c?�d�׷��0� ��U�R '��>b"�Ӈ�y?܏"��{~Q��>p!����`ґ;t^{Ց:���޾�m���=eT���F���m��$2Tj�4�p�;A�A7�l�L�5_I�NGZ���WP-���M P�%iZ=b�բ����0��b�F���G>'��Wh��JY,U��;%���0��z�˧������Ϻ> @:Nu�œ	�ո+C���E�Z���h7�a��c*a��G�yhaۃ.߶l��ȓ��������Cړ���� �}���j��As^a��?)hN���~�=K̯���4��W��b��7>K��'T���|2��j��	�S�����2hp ���z�o�����Q|?�ߨ���׹��w�'"��v��I��ę�w��q��,�p�j�8=��u0��kx�-�w]�]V�
A4�X��9��{�uh��P�������rB}�t�0����>r3��^�p���j��f�xB)�VAB�1�.��Z4٪�ջ�r�c^�\S�7n������<�<E��}���@ǳgˏ�#Z���'�����F�T���)c��R<ʙ��S��Ȯ�'��j�o��
�Dä�^�k�F5Q�����@`��\Iu��z�Q�BtNQ;GT���B/<4E�	}�_�`W��^��A��d}��o�9�7�Ru�_�	Gc�юb���Gp1���Cm�⒛�#��nY2G_�c/ݨ������Lp~��D�&)�̋³���C���;�q;	��A��vR��7��}l��u�li��=!L��[�W�Z�`I�T2�B�[f�{��r����M\�����|���0���O�{V9�"����\�4+ �d6W�J�@Ոx��|����DN2�o�!�,�^��Lk�T<�I!z��T�Z���i�X#�Q-�E/��k�ܥ��g��4�k�p���J�ߞ���1W,7�_1i��n��^Apq�[lxe:�\�V��KU&>vu�[�"�V��n\��	��k���a��ʨ!���6! hJ��xʿ��l��l<"��g�!:��Ҵ`��:>����j	"��t��BSTT	' ���'��h�Fa�Td�(s�G-7#S��%sm�[��2���iY���l���?X���z+l�@R+��e-�H$5����P�S��e���g#�
s��M1�1���#B��rlZ ���oդں��Z�G�#*0b��%u̣?v�z���U���~@d��̆b����	��w!�U�8"y��͸�$Q�ѓ�!r�v�0�軮Ω��<���[8w��ȋ����z�֍�x��m&dB�#�|�T"s�>�AL�q��~��L�bw�KCy��y7�uH�n�ba��l z?��>CB`�A�e�hi��lV��tQ��Z��μ^��e!<[`F?�E�x{*�%�"��pU�\"�Li��.��l(���� B�Q�z'�44����#Ӳ�u�a*H���B�H�X��ճ�+]
�I���BR�Ah�~��]lA8�X��1����CW(&�w1�&�-X���eo2�gQwP�H�١����_"G��=� nh�<h'{��09ҽ��X��j��>xv`9��{�x���w��(����z˞Y%ȥ�"��Ue��U���j'��.�ذ��V�0���檘y~�Z����#y�<vQ� O,��*e�Ø�y;�6J8�;��j`�gs1�$�Ё��)�tlj}?2��Ӓ���)(�Bj�CK��Q���@���"iU�J�����|����Mul_�i���{���x2��H��|x�@n��Kr{*����Z۰��bN�1)�V�,�H�B�s���G��͕�G��5�{�Y�+l��:+W?��:o���e�f1F�*S���ggB\�B�E��.�\ٴ����F�S\P�����URQ�"��B�}⓼!��'#1�l&d*��|{��~#T�����r��|�������L������k�.';`�"ȓ2�a��gAN2&-��!\�ɒ}�����@�탅�[�E)�����/��g�m��\�M��#iP'�����|A��Ѥ<���4����	������f�l�/����j�b]�I>(�ӐXZ����:�;�������¾7��'��/�����}�	�.�Y��yN��J�ʊ�I_j�$-=����E���H���-�Ln7۔`�K�irR'9��)`�;����w���^�j���U�J�~"YZ`�v]$͎$�mZr��<�f�#��.=iPҤDY� ��jU�X(�	`��ґ�p�dn8����_#�(2,,s/(C��V�ab}&�#`�#���3:�:��h_��}'�� �9�U�:���1T�mƪ�lrM�I�hF�c��0u'(�<�)U>�|��;��E�ɛN�V��y�vܰ��ŧ�ZB��5��/��c�}��A��Q��� H��=�|���o�O�Ae�Pv$4���ڐϨT�V�L��	<;$�?����t^ �mʶn�N���A�n��~�"A�s���l���8� �	�/����n��|����m1��c"/@�V�i)8(���qe��S��*�LM�j҃YK�h�
erm��?�]·��k"���Ks�:��g�����Er;�Q���Pꗋ�{��L�
�АR��7ĥM��z��r�ZvG1z�l��)��Ҳr��l��z�2�N&`�Ǒ��<�Hx8�D��h���aM�U�n7V,��`c�AԽ�[!�l�R%Ch)�4�)�@��DD<�J?t�N�X��>5���P���mЯ��㒡����r�A�������h�M�if$��Zm9�)�|�XئY ��J� k��lqZ��W�1v�rl�gی���1b��+E^��~x�}l*�;�Gb��_SF�V�B����O&����^J���n~�*'�h(����O�Xc?�B����TF��2�C�|�?�k�T���0*�uʅ������^zD���=�k[9b� q�Ry76^#(o�Õ��X@�xHQ�0n�.�m�g�R�߼<���s��	�yp���$�'f���	 (�4+�en�:�.�l�*�L&�L��t+p��$Cq챗?�ɇg��
^U����XM���A�(���_͆P���Eg��0�hgp����a��ކU��X ��CA[�ci$+�ݶϺ	 :Ǎ�o��ږ�
z���V��Z�E��~��A���t;nwl[���-)Td�"�iF&�_yϔ��/��ҋ8!j	��o�wL�Y��m/��Ex=S���ۺ�?pF��ʇ/di���Y���-ᡗD�9 �9z���яW�"����T�F�lFW�J͋�+��*Ȉ��bG7��4�А�*D5��]i�_1 ���Q"3����z�*����_��f�-W����o�j����Ly��� �Ņ�Ǵ��k��*����@�z~#�vC�[������]�F'hB�6��'a"�s�]����Tg��Y=+��/9�r������$�|�EtX��z����Y!7��$����
S���"���x�::�z��ʊ�O@��������5��_+=��[�keu�2��dW5�A�a��]�W��&���+�
?ݲ�����~w��c�Q��&|I��،��.&����VР�� -�@H|۲�� �a`��+΢����:>IQ��( �]v-�%ݨ�ͬ7g��>��v�B��2���4�"rN?�� ��MdR�F�Jh��&��p7Bz_����l�8LM�Hx���H�* R�۲;�����=B�	�q2ܻ�g��<���z"�N��B�c+PWD=2�GE�����#1�/ܔy��w`S5�!�Ѓ͌?��8�QmMJ�߄i�����uMZ�
��Q4���{��a�\�c� �iLa\n�����C�,k#��ޡ�H�i�Zq"���E���������ծ�|�$��AZ���k��`F-��?Oi3ʘ�\�x�M��v3�'T�&��a�P�g̀��Z����Ԧ;6�>~y�Y�Ǩԝ��~d0�?fE��O���d�8�U.�����}�����i�H�#�h�gN����o�$N0��?���j��'������d
{H�������aC����SK'�S[OJ-M��N41���9�X޽j03$�p���������!�h>�d�fqP�$m�N����A-@��DKŖ��awsJ|D���!�ٲ�����9��va!�_/!=k�i�1U|åae��7љ'�������va$$��w	��Eך	�%�;,����U�@,A��b�w�����k ;�(B��zu4����/إD��C'~{dlm��G[_������Z��K�bx���;{)�V��|���-���J6g�PI��<N��M/�O��R��|���$��%�$B��&�ǁ�e�6~׵ݕl<1V2'�*��zMf�!��<�N8HNs��0���ޖ-GeI�<RhR'�7L{m���W��Y���V��9�g!�����dÛʟ|�_�H��j5lU����@�?�A�#N�t�9D'��O�e�p �7�z_�<l#	gڻ\�Y��7��q�;��a��BK�RH�ivQ�F�NQ9��tG1Ȧzwv8q�Y�
-�䩇��)d���ݭ8��Q5͊'���[Owjb`�g�I"k�6X�F|\K@!iF�=x=f�NzB��Ü����8��|�]�#ϓ��LY~4���OA���n߂e���!���KD��S�f	\0��2�
�2�],A�c9�,&�6B�E�|K~�Z3�hG`�<�� p��gRi���\hZf ���g���A
5���*@K�h����	�nV�� vb� �8�5���#��I�9H.V8�0��R�����F�(�ΘFw�B)��{��!ϰ�J��Ȟ��V��<�`o&��i��:��@:*:��z�+II��X;����.�g�ѯ12�͡4,���&�䤩�����0��̞l����m�GF9pd(����������\��������fp�����IO�����1�G<rYȗ�ޢ�3At��z�V��u�iR.ǆ����bnq]>����,\���3��R�D��p��pw�MQ��3U�*�FF���� \�4|��d��"�9QS���c��X�w���&���"�[Z�!6 �B���[R�Y�4��|�ͪ�l#��)��{��X2�e�g��ܥK��R�<6�����=W���������A��Nrq7~/������N�gvVCɄq�J� Tێ��]���٥<�H8�;h�?w�a �Yї;<�g\��Ӵ��wo��nd��9]�:�a��)�`1�ŗ!��-���C�k�{6� ��q�����u����ߐ����7o�k
.� kwmr���}����K��I�Al�e�!�=�9~�0A!��z��
��.`�s�E��䨸���0]�r�;l�~�b#DM��f�R��X��R����oN<,�d������f�	���s�f���b2u���Th�UVR��g�PT}:�J�Y�tЖ�CRNY;�5����X��,�8�8�q�H�K��8:ۄ1S�A�/u��sL
R�C����\�s������W�w��
VV��`�k��p�4�0�V��γ���
Q���� �}
&�[�j�
( :B�w!�PjE��U�#8B!/��,e���)�����9���0�+bb��43�D-V�e����8%�iE���$������&�^!�����x�j2���{�k,4�Լ�N���E�"Ш�X��Tk:*���h�L]y������o*��g:(k`z�^�e�\�A*�#Eta�n�n����=��t���4�t��VT���� ������t���+Z��z= ^����_%l�)��l6����h3L醨k�P�b^[k�U��o��!���*�ï�b��DJw�k^�Ҁ}�ф�9R��S?�����Q^��7V��v�>��4t��O�	6"�b����V��Ԙ�{���NETT�t�T�$����kW2��W)���3�/:���������V���m�� `���{�5��	'�yh��%��;$�G�+�$����5��U����A�Nm�6�z)��Y\�]��'���"�jr;R6�E���}F�㺖pk�.�=��?ϙƖW�jHU(�\O �Z�]J�{w���N��1mĵ��I��ȏ��l�i S	�@ǆ6��m��M�������6�����R�b�DRA���oe���+"Z��S��aΉ_/?�������
�ö�'L��3=�g�w�E<61&�k�n�����W0�5�T/]����`0�t����>� �a�M8EV��|A �ٕSq�-��{_�@�=�T����ch�0�_0M�"���ٌM�<���k�Ӧvn�[�e����2>����W�S�g��sx`����@W�a�Zf:�0�9��n��(d��������j�W��~#	� �w���u`�X���Ȥ)��D���W��bL �g<��py�ܪ?�����{, 8v�.�	]�(�i��a�`��Y���J��I�n���?��"�U��X7��F%���?�+a��ъ�qI��Ԛ]H��Y�W��\˩/�u*`��݄�bXv��pc�"��r[{�叓a�"+���F�K@	x�"@�5�i�rGv�v�rG�ָ� @�9����*����������&���j�a��+�*��_'1h_h��q�����]8u@@3B�7u��l{m�O.
B�������:E��g}d9^�/nlzV`��jT6y��喂
���=r#݆����81?��4h;Gr4�:\�A��k�{���<�J?LaJ�\t75c���m�vӣQR<ǭ ��S��F)O ��o
ȹ���^�m_A��Rh�\�[B������0��C���jeQ��Q :7�A���'���J=��1��щ��-D0z���k�TL�~�_H�Q�p������5t3�i?*�m���!3ğ�k��8����\��ä�G��{���P�"��,�s!�t/�
�=Z4!��4+̴^�U���
ꥦ��Z2~5Rf{�Dg^/��`pǘ���o+5�����S���Jkl���gC3�B��t��,_�������\YE����P�CսcZ�:g`U��}�E�F$�y�=@_�b:䚞y~.�^��z���Y�L�8�<��}KW2�jO,�^�����Ț߳�-�������/1�%����jU|y�����pk<+��!�e\9p!��EC~�v�n^N
�]ik�zs�T#BcP&fRW��W$�]���,�46W��X���W��_�"�T=��1��+�c�+e2��>lM�!�e��ʩ`�A�'��sGz�yo�U!�#��x�;�(�1d�D�0���s�Ѳ0@-�����π�zǎ�=5��Iˀ������K=8�3ڙ_|���(���6A�I&po0�)i�{�Nt�V#���/�I�u�o�O���9�a���FF� +��W_w�ֵ�ͥ��J�i�Pg���8���5W�L[�h���g�܆"4���t�7|����&����� ���٧0R���s~I��[;!�I0$�J('E�:t�[ٟ�M��ۥM��O�A2bfm�2��U�X�Gxm%����Q�)=����
C$L�P�U(0�����jާ��	�+������ؠaӠ����AY�)E��3C�BJю�S_�cF��r^~բ��C�V`���r|�k��23���]�"��ێ�o2=x��j��m���êD���_ �'.��L!-^�C�ُ��L^BY/��m���������""
�Kn��.�1ƜwAYn�O�y"��NC���C�1�i���ˤ�]I����ݎ�:�|`@���g�	H���U��2;�$eϣ󀫽�Y�wR����mȭ΀�M;����E_�; 7tc��]�}w��s���Ԑ���P:���9��0~t��]��!��%{��x��4Y��Q�I ��HMȎ)��Y�ɬEd�l�xG�z���p�\|%�������77
;�5��<^e���tMg"�{�?��5`.����5�c�l�VìNN}�}e/��:�%�Ň�j��Ou"�L�]PO��%#��b]��kռ�j�$����}p�%�eN�9:���	�K�O�14�!�H/ϔ5��&�>g��_�u-WOʱ;Bi$��I��[⥟՜��������i.���\+���)���E���+�u7{�w=�W�uK3�B��:�	/�?�
���������r8qI̺���t}���0��͑��H�#4�v��ڬ��fl41��6/\Ԛ�����(�� ��bӇ�*dGy�|��jȼL�5���y���Ǥ��K����8�4��/B� <:���������H@���Ŝ,U�n�ͳ>��Dy,4Y�Ĺ�4�"�UW��:=���]�/�ɕo�H�teGZ��mp�\D9�P�G��У��ߐ�@d�Gۚ���)���D��qH�k��^�R�]_i{��7Rb�".�D�n�0&��M�xF�so"96������ǧ�ߺ�¶�
�ۿE
T��Bsd���(8�V����be �xX��Α��&^�H��=�C��s+J�o3}��M\ei�S���L�ԟ}��ASo<c��.�X��e�r�a#�EBI�X��k�`8�����Ϙ��sW�8�@�xfu����:��K[ͪ�y�7W�e2����O$�GZ5"w5>��#{�����j�m+jv��TV{Z��hT{���R�.��L�󏘙~�C7s)��ڇwM[����HݤgX0[8������5�T�ag>��<��/U����t6?AOU�u�D�y���l{K>r+���8ݐ�1�k#�L�a��<}%hk{%O�%̣��|�(����
j����}��0v�:]�R!��n��*y
M7�)>��o�]��]�tv��K�$�G��$#����}��'��	��D���zq-d$aCoE����/Ԕ�%u�ebY9bXS� ���MFp�&-O��W4��z��ִ���@�|�Ucz���n�&�-�Ia�:��#i�t�:�MM1Ī��ӹ⭐-�g�M�Dc���J1�왺g0+]��BWI���@B*Ւ��*�Ժj}+�VZ��&͡4Hr�V���D�{j�[���Em}���?e�����)5`�!	�\ ґ�Y��*��b��y�� /�y������Zw�"��8~d���?�:)hF|l���g��/*���:W����e�%�ey�4�Ҡ�$��L6!��]��ЪrB��9+C#3�Α�jN��i�J��h�8i�侱/�,�̹��q�A�5�Y�0�D$�]K�;m��j0we�
.-�F+Xr��H�\RZܢ�-�3i�=�p�yYv8�'���/֮�a��{J��*�T4oH��nk�m"��L83|��z�ʷ�UD�����Y���	�U>/�#Z�&�� @y�+L��Z/tK�&���@̦�f�����*Lb<C>�zn�#���;Sa�CQpv�W³
7b`�c������QQ�D!0��Yr`ߒE̽���/"�K�gec�բ਒�0���b�cI��"�Q�%^^��JH=���g�S�ԃ�t�tS�$�2[��PP1ck����L}9��PG��t�>l�=9����m�NV�/ .��1�3A"%�Q츱���8^��ʺx+��4q2�9�ʹ\��%�c��&�ɔU�!�'r��Й,�p�Ww;^��!�$��:��{f�>|x,RpWMs�dRH*�ߴ�d%�m��F*ۈR�@g��x�姉�>	򃒙u	,���aۣu�6|�|������(�F�.��k��4:=�L��5˞��z����d��L�I�]�1���6��;AL
K��u�P���:�	��_w���$��WW��-������-�p�n��הZ�D�=%jC��Z��QT�`y���_�ȾR�9�G�'4:}(I1eOE�P�r�!96�\���{��^�jC7�۷K;����nx�s�+�x���,/�(�@��q��F�9��%��*�ֽ	�P�v��b��*�`���α�Nʤ[-�8Ge���������&�[izt�!J�p$c֑�l���,��
��M�h�M$졸�I�f&���mT����0�����j��Y�c.\��ބ���u��Owd zl��k�� ���Ru>��R�B̯W����*Zv5}$Ծ$df���xg���onI��({�z�d���Ⓘ��[�$���`��Y=�$�������J̶��5�C5��I��f-iX~3J[��U��J���,w]	�a����;�*1�`�#��u���q���w*�)�$��q�r��}����*&��@�Yw���?�F��tj⸺��f���B���Oػ$uɼ2���,NJ��G�.� m^��� �|pY[�>U[I�=�I6�j5w��Đ����k|lv�[Em[��*�m:̊pO��mP�X��v.��9|���Q��	�eWၻ��nn��C�"$%x��DϹ���]FLv�^f�R��1 �v��<���ֱytW�=�V���r������d�j}Gp�s�)M�|�=�� BB���`��µ�/�v�瀖� {r������/�x��p)9��$�vN� �j�[��O�G�G:f�,sk�p�	5�|��[x�+T-ڶ2�����+큶��<�{�~Ϡ���0�w�qxa`����ۑN�?N�����5��d<����B��/͛��{�(x�is�;����&�����
�S^�F�<%ѽ%C�ι������26.�0�R3��D���/�C��п�Y</��F�+��vS�W{ᲣyV)�0���Ya��3t�,ߑ�G��sy�݈k����D��ԃ��d\�q���?��J0��ϰf>��j��<y�w11��#�+� ��KC�����D�aǺ���D�j7#�wo����}9������?��*DZ��Y!F��p����Ƭp�Pg�yNd�z�����˝O2� �Ql�r�0�;y�#OH�{wb�����^zi�7��8�^�bU��zI�� 1�,K9�J�l!�B�x��*�z^����sK�17я�Df�7r)��0N����S��,V�	RwG�$�7�蕻��-���I�ٗ�I���k�d=q��k���)��c��v"u.���1|��4vqw~�i��2�5�$����\����p����k]��{���\��D����,�W?�y�$�mɰCa��q(>�>�"3�v�.H��[*�E;B�%��Ա�Z�FB������J?j����H줱~��k���pt
�^=J�����?��2�P�h�i:sX9��%��$X����w.��iJq'��%%k�#J�Cw�\߈������W���-gГ�u����d�M˝��V�5Ԙ0pOIu<�-�[��C8��'f��T�$�ur6���d�{<���G �8���b�Z���r<�k�	����v*0V,����L�X4�̝c ��b���z�zd��8�E_'JS�-h�ٚ�є4{���*a���W�r�A�p�l��)O�ɟ����5����j��m�BT�{�z��(�>jaZ���xrJ\�ṉ� r2� �H��UylCPQ���n�J|/FܻҦ��oL������g�I���Wd�"�z�3�����J?`�#���,ْ �dQ����g7 ȿ���PB�� a-h<q��N��)`�p�,�d(�¶U�.&U��լ39R���j3d�3{�Ų�X����� ���w�k��׌�q�E��ѵ�{���+�նW<xշ�:������������?N��u ���I[vQ<XO�l'�5J�uI�{�`��!~�\�?�
ZY�v���������/ͪ}�x5�.�[AD1�Dh��4�zz0�զD ���$�;�2<��p�|�1��,!� ���Ep2��x��v�>U	�K��G����z&(Jz�+��%����B[��Z7*�=C���RZo�;��:�3��wxg�R32��X?!�"���E� x��I��_`�S��r�>g� �\%E��r�V��!�:���񗐵 ��+|o�{�x�M��2��I�If�>�{����锜�J��w�J�2��o��*��h��߼���
;3�R�����n��70A�A�XkY^D�P��q=$w�:ʀ��&�F��Iĺ�JϘ>B�'⏘��n��-�hv�]F|@���l�H�(;]W��y~H�܃�յK�%�A�w¤0�[x� i�s������T/� ���ˁ�t��:�Qº��|Ng���]���u%�Y��vd3����o��qU��.hqT�a�h�KԹߨ���%����n��
9�( 5�8��c&��LS���@6�)+H�͹,&+rCSO�$��đ4P8-;��б�n�4�ݠ6�:q�0�j�W�KS�? ���*!�
�$��W���Y�4�#�@kL�D��F�,^��쁁}xחmy�|��xng������1IЌzo�Z� ��A�g� ��ȵ�'��E�<Ά�0)|5�U��vy��E0J��� ����.�)H7f0�*S<$ݐ�����۱1�R���zЩ�9�$���V�ϻ��!~�:S�iZ����{3pǺ���[�0�{wh��=?r�lϿal�M�:�\��l�X�.tTU76���N�C���L]�/Dc
Q����!��¥����]}���[�~�=��=J5K��L�)QA�����J�8�OE�A#��.[S��u^:6˟�]��w��IJ����Ք���f��|E���P�����pyla�q+��飬�l�	]9Ϣ�t����0�,(sS"o��+�=a' uSY���}7��|[�vüoI�B%L�x4�zHC��8E|��E��)�]FWL�FHW�H���᝝㡰�̢va�Z8��C��mFU����<��_�N���?����2:�$m6�H�I;�~ɦ5����,�8��{\���~V����eU��hpO�3	�W����SC!��a�ĦJ�?/+�Њ,��H�-����	���i:�;�B�� ���9	�Ԑo��R� �gk	h�o`B:UWģ�O�-,�u����f�~�pq��Γ<����t���S��0<�q�|U"��Y��!=����n��e����<�aj�5��0���g�&��d�ւXZ������Q������-��bPě:�|�a�B�۠8�fr����RW���K��