��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�?�"|��lQ��Fv��}��|�T����,A���L{ƕ4 �B�[u���1�Oe�3���ٹC����V�v�AؗN�6�ۆ��IJ:�{�H�i�3�r��%�\� �]!�|N�b�� z�ZD���-���n��'�M��.�I$^�U�&�8��r��wl�����?$ \��EM�ph57�P��@�[�b	�3s3@s���:�̖�lB[%���b�tm$\�#��.AkIv�w�f�V��E�Z2���c}6o5�ؗ� �u����y�l~	��������P�;i�݉���_�>q)G���?R���kxuEh-8�B:F� �ׁ�f{��_�IB��{�84��'z��{߸#`β��N�p���X�J4ב�*U"���}���_��ׂ���T!�u�k���i�����E=LoI�?�c�~ߪ�62�-��ug*A%�X`�Ԁ+�,�'b.j ��'�����]��v�e�kW�g)x��W�_.�t���jL�P�`T`��9]��[���J�1�9�C�F��<��o�̼p��Y�M{�8�gVV?.4�x6��)_w�Ƴ륂����VL����A3e`;��4���Q�����yV���+|��p`�����/מZ���\8�4�����*DW{bӟ"��9t���&�����F�ь�V�5��$.��֍�eo jT��Aq�M*���*��'�ܯ���x�2�F��8hf��{��:�h!��Q��>�0�N̹Y�/��� 	y��XHLGEb�W'�����J7C�V����E�md��6�4�C}��5	��m���.�����ֵm���Ox	�cX�$#w�L|����@Z���Fg�X�,هO�W��ٵs��!}���k)Hރ~얌���Ҍ�w�dO:o���4�1G=ݘ�V ٹ�P�2����>qC#qk��4��mT��tk�Ü����8�=즠k��YB�%gSIc�ϕ3��8�r �����.X�}N9GxE�&HS�=o	i��d�%����R��!$��츯���h�4��K�S������!5?u�Nn���������3v�Ul�=Ϻ��}��N�)e>�[�I��B��W�U�����O"�������g@��m`:	u�Z�DiF,�MOX/ӏ��d;`��_8C?%�>4:Q��w�5
��.0�}熍7��a�Q����[)~��	ADB`��B)*�r�-$«���h\�Mp�z���;�;o��RW���Ύ�'�4=v����"�W�CWi��Q����"1&M����6��0�L��Cg��'��7���3s���+M��`ۉ B�V��$�rhH��{j���R�]�1��l���^`&�MI; ��?fw��ҟT�hH"�7��f�r�R�����-�.��"�WA�I��>���0Ey�J
-<[��d�*W�U�H��E�B'��hd� �(��q�44��<o6�?S���Q�:ү��Y��m�\�p�?H�0��@�>r$y'��c@
��ސI #=���&�mk{�9T��7�Y�9I߰^2>��g��Nϻ����ILR��*��:�+�AYZ/��T���u�+���0a���:�/�ǐ̻�� %V�uT4?K�넷�)9��	Ы(0cХ�!����>�FL�s�(�v=��RŔs�G�6B<E�[P�Gf>��j�ch9�V��m���p%Y�ո�'�����Qt@��)@ڍ?��z%�W��׭>��p��]mk����\~����"�;%��6�o���pkì>��7ZBtľI~�?E�<I�:ض�{=KJ�~#�� �^WqP�K�R���\g��w}�9�ԧ�~qU-�qx � �f]���V�>j�So���Tˡ
��j�����t�*��d2*c��($�U���ӯ��?#���A��3yr�Ȣ����Wn*��,�s��y;̱�[���e�����z��R<��BdZ�d4q��Ęu�v&��̦�R4�t��H�3�Q��݃�v�i��#1[$��k�B��U:� 1&��Yйv���>.�C���ɠa��n����F'�$�%_�hX�7�/>���T�C��N���>��������ww��y( �|��)���D�?p ǤvnN���!F�Xy��C��WJ��V�7�X1=�m�q7���;��!���;��� *��"�B��"4�Kx���I�N���9��@����6��d|R�H>��#�`rtk�B�%X��O �?��^�%�g2�(h�Q���Q�pT���#�<6��m���'��H���B>Z;���Ȓ�{bT&	��ɚ��|E�����sA�I�?s_� `��$��E�!bG�G[�x�@��}F�����v��8�X�ΗX|Ι2����WOD�Fe�ǒ������d�Gk�q��(���,`����r�h�������"�aSzدi��A���p���/�d
�fn��)��1���� Y�7�E�js���1�����8nv"R�ʻ�nRX�o�Q0��lTW^�q�k��g��J�+� 	�3���`+
�􅥵�u"�(���G\����h-�c��_����\��Qi@��lv�	�5&�x&Ⅺ�?�����m�����U�~�LEDȥ��vR���tM?���wX���w���j���~n�En���rB� ���@�:���Ë��h�B[LO�����ŀ�AP�q�27��8�q��V8r���R��a��(�oh++d��<`�~= u-8�C���!X4n�[<J��_��VcQ� pfi�
ۛ��鷷��O�T2��|�T��gk;)	�P4�uC��|����wOUx�*]u:�;���R��q1RlMu��x�
\d7��~��$���\V%C�=f�oc��Y�sB�����P�W)��5K�aˑ�/]��zL�4r::��m����_����`�og&rp� ��� �j C���4�x��n�����2z/0@�F2-��!C$8�@�$y8��������V�U�`���BFXFU�,�/tA��R�O^Ȓ��ɺKƍ���i���҆z�֬17�k�hjH��;L����Nh��o��� 1�\s�����sދ�P�v�)���U������p��6ۜ��|Ԥ�i��յ�=)�RU��`ɼ[��,^�/KkT�E������.���~��9��O��c�������r5�$y��� �4��>_6�i�N���xs��/;Ǘ��z׹��ؙ��\��,�h	b"�v��1��'���Z%��:��m%��jc�<|t��<��K�i�)^�	���zYcz�5��,�Z�o���Q��� b�go�=m3-�����2v��^\ϋ����M�zQ��V���"�u!/��>���Fp�f�[���}༸��t�-]����@{nԀ݃A�涢k�2A��E/�>vz ���6�-�g;ޱgَ���C����s��b��Kb����2�o����)/��K ��)�~��x�U����4�q��2Ţ���2@�������,�ף�e-D���f%#�o������yP���QT�p|�R�D��ǧ����"]�8H`��z'���S�77}LVś�2q�륟����������?%��@1I�JWף�p��yt|"���MУvy���0CHE�I� T"���<�R�]�5��w��ո#�=r�Ǐ�ԙ$O�cE�Z���!��ލ;�|�c�`����xj�x�<% C�,B�3�3��#���{�=��צ���_#��ι�*dVA��E��}4N�y��@.�z�)Z�1��MZ��o�L�iw�Tm��6�(
�/Bf=T��G3P���3Ý-��E���`���߈x�a�cf{�V�"���M��p�>b'���p���Ƕ@׸ bvS&GPƜlAl]=u�?bG�M`���D[�ι�3j�C�O&mzF{�9����!
�q+��CmhIj�RMR�=F0���+�ewiY� �d��>�G����w����E��]]���8��`j~��$ޛ�B������|>Xu~��?Q�hQ��<�+f3���=k�w�q��^�B������$b
d��S�*+'�{^��^��o.�!�A8���r�D�a �^��b�qqw�#m��נH��`x~�فi2��x��d�ܘ�������,1�]_�����c�hK>�>���5�@��^��T��A��9�#�k�E�]�Y�(/���]"w>|u�"��}<��&H�a�%����P^�n�v�|��J��&���`X8Dp7���vy�cuV�lf��H�3���А�E����_�8��N2�_�?zQ��aЄ�
@���[o���e/��p9 ��r�a�f�f�`��,}��\\��=��0N��z!YTˈ�הz]p����]r���GVl��A�e��4��H#T~���M�p��G�,8^��'ˬVK,����'h���7������w�ˡ�� ���:�0Y`Hl$q���v����a�?f��#^�qs3A�m ��3񋱚�k��]g��B��)�<�j�Q�]+�(H�'y�<�c�AnG��c#cLҀ�Z��N���O���Mt2�hB;Gg	���anZ���yI����G�">�1��}�?ON�����@?��p�����P��S��^B�_�����	9�E}�bV���Mn��Ɯ�*�#�T�����P�g��|-F@@i5 *�M	�D	2*h�����D!�ѭ����I��87�Ŵt�[$Lk�B �t*��1'������o:!ީ�,�۬��x*%���(�	;�"ci���Oi�Ч[P��&M��of?f%������:��� ~&���3꣄{�����~^Vw����'�)G�s��5H�����Ἥ��S^��J[a�^Q�����#���Ex�8�̹��BKi�C�i��b��(�0��E�u�^�d�e����_�:�N׸�����9:�*�ث�n=�T��>���ҋ}����^������ŋۿu�	-Y 1���'�sn�Y�j���*��p���X:�$��Sq�����Y�V ^'�������cA�'��%rx�8�t��^�������^Tz�O�����q��k�-�I�cY�f�K�UJM�<^y�b:&���6�b��>�|��v�m�E��i���4.���Ȭ��:7)~�w�BZl|�WwǮ���$n빼�~D��y�:WG�eh����t�Sgbp�}����C>�_��x��LK[u4"A��R���~?T��r�<$�~�l�JƎ|�$�P&�zڣw�E5s�������E������4�+��i���>ޜ{r��WCLł*����:\��
�5���2�/�YL���^֮����T����:�xVi��;�Ta��+��"��="NU�����OS��~9|�Ⱥ|S�i���Єm�+ �X ��iz`I�F\�(֬�!�S�wR0�D 7�����^]->)cAV��D��D�?����~�)Zb[�*^�G$m$���ǂ������M�LN\������$Vl	��adn��uvZ�*q0"���S��3�,��%%�hG��&L��T��?s�̖?����7P3 �����#bUo�3 ��G��˥�2��f��3���vQ���E����hM��U�\<��g`tuU���(�8��#-�!�	+CH�^k��.P�z6�N��oUp�"0����A�M�B�*R�W��H��N)�y���{虶�*
<��{�/(�}�3,v����Μ��V��de��	::<7���3nR���d�/�y�'�N�1L3�d�"����6����`_4U�ԛ8��:����xe��M��x)�ج��]9�A�<�.\��u�����^�:��aΧ�0uI=��v����#E�G>w+���O���`�2V��bȀsN�Z;�0�1�t2��7����J{�&�ҕç�F��-��աOu��)*xu�77z"��C*&��r ������pn���(��'�Ƽ鞨Pd�O���N�("��GL�:;�o2��Ƞr�Z�Υ
A��*�4Z�:caXj���]yp �	������J�|�a2���e�?s�7j=��`��-��-`�Sdm����{�n:�u�B�S�'h,\�<�D0N��Y:R�W˘ФP��Ѫ3��ft�b������>Sr%6�����\h|e�A�	mQ�����b��J&Y&x7:���5+ӗ($����\�'�؛j�C<x���]�տ�7����Sͫ�D�`(C�1Xz �U�&�S�x�����kJ��������;�d�q�}�c��'�]��Ou;���o���b��rS�G�km��#sh��JQ��L��#��7�!M�9�2��"Qx���������hq��PЄyV�P���F٪�0!�tdq>y��+�̢��䠇��E\��Ǆqu4�ǯ������f�+fk,��T)LZSh*��s>gB�ŉO�D�Cq)�A	�d<�EP�\Qj8��^��՝P��K4�0!�H�>�k�fƶ�1ȯS)���~Tw�Ql�0>M�_�F��s�7`iH}$HË:��d�%j�B¹��s\̎��'d�����p��~G@	�>cx5��o��TZ�$+\�@���Ra�"h��1-�`�.�I>_�ꧫ�zw�⇌tj]F{m@�_�Ճ�r��B�iS�|�)�{B�j��As�0����pA�iA�����=��v��y��PID�-9=�q�&�K���8C��2��l�����o֝���O���i�j~A}±�&[��쎛�U]bLGG�
�R�-���%�����\�W�k ����gp��A3酟�𣷷)T�3��W�`b��0�$y�f�72����=\E5-���_�im���?�� �F�S�����JAhR�l�[�d�fk/��p��.�Iv���9��5�
��-��6�3���<H�eK� �����R�( ������V�:
&W���F�Y\��PU����>�6oO�����2��N�$���!0��G���cr���+���G�eP���R��4Š,^&wg)�|i0�����zj}96h)��v�M�U��@�����Q�K9� �T�#3��1��#pqu*}BM�mj��i�����^�&��2b&�x�S��L�ǣE�/aTa�W�$���$T"�v"l�
X(�N��+�I��.��.x����]kU�݁]���g>��LF��5piI���t�^�� 5��H)�a Y�wv�d.�F+w@�Tܟ��ITq�#�z�r�)6�l����=ٝPѰ�xT�=�Wxe��II�aƿ��	���E�(�5���7��a�xm���"b�T��� �T������+�>�_#T��Z�0; :|ۓDO@����s�}�նuw<�>=��_?��a�k�G��(�s�3x7lN�,���%��_︓{n����1:��G�a��-�x��ö���:mK>��@������"���f�\�M��6�F�f.L���W]"�&F�o-�����������`Q���Ll��i��&"�r�> 9ώ� 8��[R�]�1�܂�:��\�B���U9�L{�R"9�#z�t%������$_�/�H+-1p� 9�t(b@o���j��B������8�,6����}���燨��9��k=�TPÓ�w��躽ῑ�_j�\�>2n.��Z�>�O Ǉ�G@�l�)��b��ѱcj�ԴĪ�	0ۦ��*�2���%�@�SJI�Ѿ�-I�g���Ro@��m�6�����������t�gO�:�7�/���F��)tc�>��<x(��A8���7C�����"W+����X���-���O~I�o��X��ѧw�TM�:�ڙ����9��,~ ѧ�BJ�{g��A����U���;䝏���Md�����D5�1��z�1g���m!�.��R���$����>��]��0D���������� �YSy�}6���d�}�*���b)��� �eO��dA��#{��TB��쾘���H���ԑ��"�I��o���)F��?�G:�*5hq����*�����2�Ϧ*Yу��b>kREu��D�ZN/��t�{<���g��/	��,�v^V^��#�Yp��t�N3�{�^ſF�ӏxT�;FU6���.��@W�J�0P��fl^G�gG@
��r�"[�D�p@�;H<���~�	rRJB��L9�O ���n��3�`��T�4�l����[�0�C��b��UX%�p� y3j�.Ʉ�n-ܭ0�~��U�4z��̵�Zitv@_���~B��hnƕoC�%����ں��3��t�*��ywL�bi����U��MC�!��|���not���4���>��?�J�~o����jM���T�F������?̳ :νo@��D8� eVpHR�H���}�K5�\DI�/I����z����?�x|X�񕑳vP*`�(]���*��0Lˊ��H��B>��4y����-(�mTχ�Bl�)�׷�)�N��FZ��s�3N�*�WG)m(�`ml�B�5"C(��X��CwjDU���ɐ=�RI/���#t[E�ƙ�S�fǀF��P�":�9�3ަ���𾋫����gR��U�ۨ��|�N�D�sh��A�l�^۔t����n�!�Y�]��%x��	�ӫ���S�������č���D�%��c�H���:�I�d�/7+�ކ�)2�C۰��͉2g�2�2q.x,R���sA����=� S���n�WD�^9�t,��*H-��o�9��}���������bRWǢ��(y�5ttXhJڧ�U��s���;��-��6���ڙ�lߵ�R!"ܿ�_�c*�����
s^:6:�LL-n7a�x��C,�<P�Z�O�ơ��g�-Q'�2���eQU7ݾ�����(� �3|d8lr�SsX~���k���Mc���q8���	�S�eA瑏������<�.\/1�Fz���U�H"�R��n���]܁�0���@)�Rp�Ԇ������$o�p8�r2�k'��� �`X���	qC����&����ӏ����I�m�>9ޯz��W��6b���>}�_����Ǖ�R9d!�`�xW��3�x�!�h#7A�=��;�����>I��(:r
Hbs��Oko�c���vM��������	�Ą�_����� z��U�_5�7E���mޫ�{�Wʽ�G�6o!#��7�C'0�t�hU�����rА�4)^�d�����yՆ���Jp/5��!7e��k�롇�F�?��F������xn�Uv�ݬz�������m<p^�my�麔�Ӡb�Akr�،ţ+[)�!6�v�oJtr�z�g������{�7ڍR�'ؓ�/j���!Zѱ#|[u�����'�t6
ʝ
]Snc���+�m��H/N,{R;�2?L��*�#�4T� �d���.��1����Dr����
�V����h��Ge�bYp���U`4���[���~P��)E�Ej�e/P]vA�$`:�8���h ��IS��Y�o�a
`or>z�Tw`D�Q	�Y�[.c�"�P���i�	l�2�_�m�4��Ew�jі��V�%���氲L��{�[������U1�Q� � ��y��o�;�+ػ���ժ"jDN�0*0U�p�F8a\#�4<�-���a��08�EXh��݃��n�b;��a���(�Z<u �$:��<��@Q0�i�?�X�w�� fW�d�@GW%�H>V�'����m؜fAk��i���?���VT�"u�:b�ܒ����Ԛ>RSяu-��νB�)E�H��NS�R����������T�����x��YE���"�D�I����&l#�`W����)h �P�ο�A,�:c��� ��\>ܩ���ۛĪ�۔n�T�
0�C���T$�zO����m���}�m,C���A��i��D�ߓ� )��P��pbDY�eKpKcx�qXΠ�$LfJnp �?(i���/M��VW��8&ȔJ!l�j�ݏ��3��K��ԈƟ�"揓�����:Ym������%<�$�!s0.����"��4B��<&F����Vؽ~w~/$��s�ߦ��Z'����Z�J���]��!�y26���0�u�7C�M��xDE��	�<	HKY�-LB�桄�4y3��>�F��"ZY�M��G��;�xpH�)��ݺo�Zi6��&lI�
��Ǫ,��8V1��<*š��LgB�w�>��RdJ=[�ڕ�XX�����u²�R���^W��,�PE�[����:%̠ܷqΝ�j�a�l'S��ڐ����t��B���
�(�|W��o�_�J��ܠ�؞}���>�4s��� ��Ϻ �#��H�t����'rv������������$�r�G�"���zD_�*s��^*f+��������7�� x�4�R�9$"9JFUD�#kk>���=���r�F�y�To��m�Sƪ�*���E�s=���v��8�R��
.ԦZ%��h�yj��پml4GÛI�C��+" �;��u�up��i�Y"���NXn�`��z��%���h�W�tp�Q�[�@�V8�˜�~��Q\wx��X{u������X'8|F��!���rt��گ��o���G����}q�.�ٕ��� ����Lē�M��*k�VlǡU���Jk
4�=d�piq�qlйk��U(�bY�8TZ�g�nl^����(�9M_sR:���(Č�b�����Ϫ����L�h����j���*,�j��N&��Ԋ��M�R�H�]�r�W�j������c'�������|���[pB�7�Kަ��=�Q:.=�"��}��O�ɒ�=�q39�YP�b��4���z8�Q�p��q������22���M��;����+!�>��8�t�j�\`�&B)�<���W�L�#������)�K��';��榫��W�gSn8��,`�q���8�3���1�ۊ��M��������c�P�����3'hBU�w�1%<Uu�K��v�%��k�9�e��ȑo!qz�n1�?�J��[K��/�(l1曫K�t}6��T᣼t�Ξ�O���)Z+[6Ltb���[�����H��}w2߄p�ـ�1vb٭��_�lȦu��P&�����e�9���7�&i�e����U�d��c���φRj�/X���e�~�C|�dZ�����'���qm�p����Bw�8Z���������Y�`Jt��A�v	�_�i?售��X�8�9O��ث|�*+Ӌ�:�Gmkc͂]@�V����ƛ5�.���&Em�~��C\.ӊ�1�BF�S�0�F7\c���M��V�hg�YMâ�9u\Φ��+g�@�7�vN�b�J�!d�4YUTr��,��������6@��U0썲�
�:Æ�3���g���ki��٢x���EN	�����ɾ� � �	R'�3+B�.�!�Y�_�O�Yk�)>�F��3$	���_ߦL��~�8i Rw�W��lj7�C��0܋?|
_[��*��v�Fsh<A��n)F�t�J<�������0����.� ���n2S�>�$��J����XrE�U?�f�ك��������<n��L�4��䐀h\7��	��0y�Z�i�خ\U;_P�NN,���ʄ���IjT>�BQ@��k॓<�����+- �5V�D���, �R�`*�����2X�:��:���0�y�is�Oj�O���p�Ee�B+C���	�b��v����N�`��]�ڜ7�F1V9jz�q ���D�_f�\_� �6Ѭ*DHj� ?����?(�z�e�1L���2��9��I+U'��ח��$S��\�Z˾�hs�1����n؜�� y�M�R�s�<��ɘC��]�_���5�rYΟ^4���P���(X�������'�R��-\�?��Y��y{��З�@|�'ᬱQ��1<�fz6�|=��lZ�؄X	2�1�����eC�%��9	��k��*�c�皼hU��@���PQ0�	Fǘrc���k���
�p���M�ߟ�ni�U�RO���"N�6�/�tU�D�?�QN$��ND����.���4���4	�
i��{.�l��֎ @��7�m8>�peuI���V��KX?ժ��^u?Mcޯ��c(�D ����qdD7��(q.���f(<��"#c5J%9���ux���W+�r�LǼ2L}���(qJ�:�ץ���]�qD��^�qܹU��Yň=(�)5���&�<BiU$*tR{H���KК�"�YU ��}(���>hP�N�����Ekwx�P�qD��zhXBD���w���:� }4�8V�h&F����(d�G���f����B�9�����tz��fC�&�<����0V��� ���"���2Q�4}���.�:�|��@�hUa8D�[���;4��w(�c�Tc�J|ռ4�����?%�J���g郘 �L����vO���#�p�T�2G7��W�T.a�B�(���Æ/�|-��ď���Yw�%ݖq�U��� ��6�^�h4Z�W�m����Π�8b��	~��7�{fI��r1�$e?�X�|��)L�Ƈ���@�ֺdH�xRu�ӎ��r��T��.I�X����@Ȃ�@���OH��D2��1��Ї���2Sl��f���%����-�n�ic���+��u�j���_��JR�^�����Y��C���y�����~`j�Y?4@���!`�ı�Ձ�0[M!��Z-�0���̓4��A�� �I�?+��;8���w�'��n�iw]j�nb^_,3-c{���r������c؞ͳ0\���f�*-�@-��9�H�Ru�� �����|�FoQ~)��x�k��7Ng�5r�x�8P3���Rw(,�@uG[������\��p/?�������:Q��6j,b��6߇q�^���A!pm��N��P�p4Ǿ�E�V*>�~�!�|}7��6Ɲy�-�=R�����R�2��ne���[rP@�T�<5l�Y����E+�����L���͇�����;�Rl+�Hf����vqɀ�_�_mZ(�K�"�z�qPX�e/P�D��]V��:�߸}�g�6��W�1��o��K&�l���G��XY����c3ƚ'�BK��Ďz������:{��S���_