��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX������`=��u�#�{�m �;�:־���(���.�t�3�ya�V��s8-�2x��z���������+ڦ�!/Ӂ+6�C@�#����P����B�8��L���ͮ�tMs�v�U�8��DG'��k�t�7ZV��j6����OQU4�?�9��V�y�?�W��M{{wi�}��:��ml�]�	mX�R����S
T������zh���G)_������23�k���/��	Cȯ�+�������3�� �h�%�X�4���T@��cx��8��|BSU�2v��KK�U,��+H��yua�ǖx���W�SH�Z�H�9�7/�`�Bt��>��@ꘗ3�q�M�@m�� ���0
�0�[�G ����&���"���,c��t��޻���,yyj���vQ�D%{�ä��v��_���%�Vg��h"��X"5���G���flc�g�����2��,�Ќ�?]�pD�%�xR^�}ն�:I,����1� ���?��F�ӱ���/l��0��zv(�<��� �_�q7��(L�W�siu( |�î�ZU/�@�����G�~:+�7*���钝&?�fJ��Wu�In�j㛬�D���W0[Y�P�{8>+%�DL�����O�v"�d����6��O�1���?��O;3,GQ������U�̆n��_��n�	cx���Tʀ�}����[�
�A2�Uf��\�8� t6�������C� \K]n�*{÷�?�"J��:Q7F��щ�a�>�w1f$�[�r;��պ���>381;8A�/�կ��PgHGvW��|��]y�8hȊj"�LC�'"O<�8*<1�����_�j~B�
k�i��M"�&&���3L|����K�٠O,.�4�Sw&�jP�R��������~9�Rn�c����GH�� �,��aaZ�'˟)��y@p�=��7`�4r^��<G�uJR����mʦA�Ǘ#��?�3�p���ъ֟�u,Ly5���������b��:�$>����g��V7w�<
��%���G�<����6B�|��m̀y��OB��l�)� �M�a�pd�ɊO �5;��$]�*������cpD�W͓�%�:h�� w�ǋ�ٯn�ڈ��<�RJ�X�¡Q){R�y��n:�n[9G�֏��^o�����4<R��M������D��ﾆJ��a�LWn�t�v�f��طya��$�f�)!�\59{�Q��U�m��M���#m���W��GP}Ƿ^���cP�t�}��bte1��M-HƬ�j�3~N��eGȇ�����?f�R�g�sm��!Z�2��(�'brN���{f��Y�އ(�8ȓD�P+���]5({��@�Uf�n�k>����?�ly��L�_3i�F�`�	?�B �ϳV�U%��^ �ܸ_7<u���گK�?:Ih��O�C��q��̢do ��K�חl�����o�1�[8�g��5w������h��bwP��G`���?��o�"�[�Y9E����ԃ�T�o��]�*�_��x�h��H����\�Ā�haOӋ.z_��!˲����v��r���<��:p���&���d}��ˤc�Mt#�M
���7mڃ��������|�W^N X�s�$��J:J~e{�_mAB��� YJ���b:��ܺ˕���H6]g/�(qAp��Yzߠ��}OL����s�D;�;#���<X1>op�21+�Y���B�/oK�
�6vQ�-��+��!�S��Y��� �)�蹛t�E�4j��Qߥ��<2�4���/+�P�v�Kr��l`�~��_�hce�tfC�Ȁ��(�qBb�Mm�|�*:�&P[W��~���d���$�P���26��1]r��,�&*��k̋���6H�j�ϕ󠍵��?w��j
?�-���Ճ�yJaz,ot	����a�-?Ti�K��-�!�)��&����.�4�8�?��`K���)�D�N�}���(M�
������*GZ�98_�`�ʁ��0�zE�}����WM$=�>�1!=䯨5��U�9Gk��˼���BmS�e�'2�ç>?������1/O�2����3���H�Mij!mb�����U>��h��M��{p��i�p*��b�����
N�B�G���t����ޕ9q����\e9�[�ߜ�9)No��Gޖ]��Ҝe�ӥ����U�1~(�70:NF�ώ]I
���k��7JO,q�?m�V����Bz���[�h���|	�$�W��L�,>�J�UTW�D���':\� �}_���*�t����+)�W��
#5�"'�;F�
�H�C����G;�"Q+�H�	����D:���w���G(�Ґ�1�]V;���\�� �H>F
s�Ʋ�͆Z��d[˘�l��9��V�m���%�b2���u.8� Ɵ&;����3Q�ߨ7sfS���ȒFUy��-T{���PY�`�� ��S�����+�2��9 x�{_c���H�����nmu��bx����9s���r�ִe���d�C����ʆ���/��4U�r��_ߚ�&��g^�����a�B��&|*�]����i �GwMv�̌S`3g��:�S/�N��[Q�j��Q���$;R��8�쪷m��f�F��H����{�D����)V�w���^_�{ό�:6B�l��$�C����k���M@�Z�
{Z,�=9/�ߴLW�'�i�:^�g��9�i�}'9�^,�ț��,�Ǽ�;�Hޠ˻߶��6(>�O~A�����.)�lr[Y)px�?����zr��oIi��?�bQQ�������ι�����F���@0� M�\�N��Y�.i�z>Z%;ԫ�O�unq��{t�.s ��ja錛&��H$�9Gn6�_´������C����4�I��W_��)�/��~�|`Co�W4w��&�7� � ���h?�["��+���3��QZ?�2\i��Ք����,����	o:|)jr��Zx[p*Y��CM�T��Ym�Ғ�2����S?��ˣ�>�
H�1��3F���h$ծ�L����s�@�GA7��,����:�J��ِq)�.�m�{�h�NN��K!� �6|��Ѝ�H�����P���F�(������"�4Q��Iy���6�is��aRL�1��0�9�Ӯ�}�i4�	k���pc#h�/!&��ѭ�ؽt�C��l��a+k"n*Dy9oi�P"5:�e���~�,����=���f-G{	1r���L��ak��h4�b�gz|lH�z�!O1�(�U�ק�.�	.։�B�����Bd��4�y�u��I�dK�v؉-κ�S�<���o��-��T��Oď��#e��/��8a�:�Im:��sxT;O�ַܜ��ߒ�8�w�ޑ�Oq��R�����wƞ���x�L�@@1���|�ZM�Q��&��utH���3R�B���,Ӽ�/|�z��%��������i�+ ipN �r�D�=�u�7�"�f{��9"g���c��ZJ$���{1��F*u
D]d�G�(��S�j�D��)���kʬ����sL����>�F�Eŏ����A�0���C�h�3R�/�k3���bu��:y#�� ����\ʮ�ɣL��̦���K{^A��XP���!-,�~~�������.�+�/�*����-4�}��VFG��&���s�� )���a̽�Ҹ��3��6;����������:��Z{�%���Is��_�"s0�A���@�>�sqwS%z���Uڕi��T�R�f�i ؙv;��t�($�[�7�P7��N4�֬�@W�g�V�W[^Λ=��a�^ք��c��QЧp�t��s��fdOѕ�@��X/
*���Z��DD���0拞�W8ea���*�}��ѥ@Q�XX�U���;�=U�[�jh��]�  �}<�����J¹}p��$ȶ�rn&�\L)�ӝ�*鎓�� �X�¼����H���O�*�K�$܈�6!��E%_�	X&�R�	��o��YG0�)Vr��K%������៘F-��ޔD�	(��g�P�9Z:z�i7�iܻa��Es�`0� �S{K�dbCr0L��l
��>��`�����G�*S$�y����[��<ed�@�B�@��{��Q9��� ���K���,	�V���-|��ԉ��޿��*���f~	U��Tߵ(��O��a��[�||�!�&�����C�y�?�
�jS�/3-��b���>���uvΪ�[��(��)����8UeL ����D��y#����aI�H]i߆d�y�#��ЁH��uɯ�K�\���>�N���H+���.[.p��ޗ�*�[`	�4S��qh�3E�H!�O��+�z.e8o���+�ݿ�W�hxR�fF�R^6i�V+_=v�Y�_=�|�@�i�^k��*�K;$'�o0��{�����jl�-���܎Ҥ�Bh8���<�E�8�6-�_H!�Wi��E�89h�y$�� %��^�J��y	���k�J�O��0OA�ݦ'��l'�#�1{�����V�b�v�Z�p��,�Jfw���ū��	����.JVZV"2 7�8�#����E��������|�W�Ad�qU-6Q��8;v�EY^�{�����{s��,�xOKz��G�A'_��y�2��_�F�EM,5�Eo�bb���&B�0��)ܨ`O~X�����7�}�i�N~e�d�O�Z�Gס6�;�Kn[p�)׉�@��4b�7fm��/�0/�F+�M�6���^��DLVn�<=,�ބ'	*�����-ji��|^n��s�?_��@
	�ЏY�*uAr�N5�_��D��?����Z?:M�R��S-�=N�?)r9��u���.�#�?�hq1>X�s�6ώ'�g������O��eװ��>-#C~��������K�!~W�]O�7W��s�gIkh�@x'�7f������#>��z�Z�@X�P���:����Q�2�?�\�s�*�z�6�a���kK?v��	��5�G�	��q�EaQ$��\&ԽRY0�K�p"ﳇf�2�`�����V!9�咈*%'}Y��'xY�,\���{^�������ѡz�x�w?X}��E�W1��ٟ�2ߨ����Ҋdd8�X Đ���	L�<��%	'�S�#�����ѷ5%����2N��W4���`x��&^���2�ةa���w,�7vJ�3����U>)�(�����Ƌ���M^�x��:��B��2�+d�����K��"�\S �.�S��F�2}6�z�Kےi5*p��w�����I�?��X�����Dxk��)Ȋ+u?���"�'��3��~�e�щHZ3a�:gh�p(K������=�W	O%ۃq��,'
���E?$u4V���������yJ%7�yX���Zt��A a�/e��I|��!�c�
�l�{X�}��B=ީ���اP�1�%�Z=<�Y���
c�Zn��A��_��\.;٤z~r'��b���	�Է{�_5ԕ�מ��� o�üVІ�� 3�7;R-�u��ɏ^��'h���\�DW��*2d���}+�W�����@���s}#�~�F��Z��g;h1�������),K�[.�����D�͂�B_�|2���1�{��v!
00��fG��Ř"G�{c��~�9�KB�0�]�y�N�����Ֆ/�sI�@B����VI�1��O#�)��Z�)[�������BngF��a���y.[:�%��/e�9�yz�7�ygt�oXsǁ	���6sҏ�OU�#g(�e$j?�$1�_�~�ѳ��Q\�$T�3�d�B��' �%ļ��C <ٝ�7y��9�!^��@�Cj`״F�ݪ���_`hm������k��/6T� ��|��5��C�f����(�5�Dfph6<8Z/����I��+^��V��hnk���۩�h+e�p�Ȧ���ff]�^G�;�+>����X+��+X��23~���ԸH�f҄E&:3j�8O��R6@����%��?|�'�6�J4Ż��Q�?0�4)L�U��S�z`���]�W���,2��Ko*��$�8^J�F���]������=�;�j�c<�Ƚ��_3
�9���X�����@L�j���\RT�4�@�	-]����WSq�y�%2_L~N3[�m��e��}N_<b�����q�{D�(�e�#�"�~Q�]�
�n��s�24�?��v�Y|=�o��J�]ؼ�wV��-���SU�<AW[�~n�x��c��8X"�P�<G��2b���GN�~���!�<�m�%r�X����eh��B��z��#RŹf� ��-iQ XqM�$F���s[�JvNd��Po[P�S0�W�����[	o� �j��6�����O��:{�g�Ŏ���Mr���?�[jv��iT���( ?/�X�c��4��R�֠��I����
�]���W7�6��ki���q|�:#���uuU�v�����L������e��c���aΤ���<1�A�IjA�F�_��N�4��ߙ�^�U%����aL�y!g���a�����fs.�	� �ˣ�y�J�:@�%��ey�֯g�1]Y�͵O�U]���߶��]=��K�1�k?,Y���	2�P�v��g�΂p�k�5�c�>�0�n���N���c��b8��¸�f��ź���+{K��c��o}L�B�Ëp�ɶ�/���'+�|u��=�R�Ϝ����o��A��No%����9?;�8�O�Hp˵-��ʵ��]l��Ki�$�t�@jk	t�˘�
�����{M�/���_�]8�c��1 b�qY%v��q�T(Nk���Գ���4k��3g[�l�$��.��e0hv�Q"���Vk˾��U��WO�ע<q{s���\xz� �
�K�N_{��8F�F�K9��"	V��%��a-����E2T2O{���8��g��`5�:Dd��B�،"i�a"����˻�@��us?0�)��&<�W!���^\9��6����߁�r����[��^�H?�B$�%#�B�p$C�d���0ڲ��K�/}*��N�W�X�e��=���*-H���mh�"�,b[% p�o�ԑ�Pa ͕iR�YZ;ś�X��H�Bnr�q�u�X�Q(R$���~~�㒼�^JoDA�9�c+侇z��/�2뚵! �!�׀��p(�]���eBs'�Ϩ��#}�X-�m��Rqh3��
�2�A�;�*Ő���􉇸�����0�ʲ�>� >���@�� �G͘�q D�w[�@�����Ȫ�j�����(��8���[8b�g|N~�O�:�2�^Q�7"J�W.������U�&4�dz( Q��5�gãҠ��<{a�ϟcR��M6up^��8B��'v Q3=�5��ڊT-m���MT]���X���^�g*X�YVѷZ9�������[o��1��sS����͏�"��j�4�k�Wf&U�L�4���x��(ֳ�=�����XĀPN�.��U3�v>v4��wI�f��U�c��!��]6;t���:�=�m�B�鞦��x#b��L�J�bb'Ө�� ��W�+�[���q(�|N4;$��p��w<�AƷ@�3�(TB.ȱ׫��ȇ�d<�Dt�	���"a���|f�^��'��S.�zT]%U/$��4���0j�r+��6kؠ
g;���8t���=��Qj�;#��<��mC��>M�ք$B1�C!1�a'�)��ƌ����dy~߭/.��PL�g=�S�7kç]��kg���:w�<.�����B��\n�.x��	ʞ�f�p��)ɫl���,�����\��M�Xd���i���{�����z?�1��֏���N	��
�1�m�l����>�UbɈ�������:��"�R
1n�� ?a"�iq��w�l���~ �UX����X"���}6�J?�#�=��6+�y�$���=�SQ����/�ȽS�M�Z�PNz�u�F������S�S����u��]�A[����Q�#�tY^{���s�*�zBB���5���`�<_����uk�G�Ql�1�5IJ������ny���"*�(��8!�{����n��Ƴ>�C���sxș��V���������2!}��o�ݨV&�S��9�Dá��f�s�'{�Θ2�k�IکI^�CE��
�v��w�u�hW*dRP �EP��(��Z��XpAf�x�Q�A�����n�J���u��u+����'A,���h�;�9���{b+�ݿ!j��n5/[�3|���9x=�'���2��O�7Z�K)(#��z9��)��ϝ��bϘ����?{PMw����Il�&���.V7����޾l˰&�Fݼ�3lj�V�wl��5�C�e�2a�1�Ƶ��t�6p�VH�Tq_��uq5�;�xE�Z\���~�)�~���&�|�W/p��@V������ˁ� 6[i5iT� ;TG���3l+��0O6���9�Z�Pu1�K���*c���[�5I����Ӯ�ف��,7�M�&$J�&#��	��󾌣�©��\����4�ʋ��VP��̅�ƼKZl��B�X�e����E@o����r��ʁ@m��G�/�#̀3��6�R�Rd�%�*�L� ��5�������	��R�]P|�u}�G���<,�}�����)��>���	�Ӱ���7���Ɗ/	�����GsҚA=ڄ�5��������i��&}�gU��	D���]Xr���.���:�P;*X@��8\]<Ea���y���w�3�RXO��D��ԤH��´[���[WC?p�qO/��3���[ն��D�N��m�r�xאC)��Ú��0k�8��U�C�>��n1��Ka'1�U���V	�H�����['�y�C�̚�a}WbȒƉ.�b-4��C�����߭­pD��*�Ï���8��>��g�K��@�0-��2�����Tff�b��m�an~���ެ�q��1�p�!	���`�i�X� �yŔ���@WV;�����#<v�d���T)5�*F�����oW�#Y�&����TF���Z|+��.�1n�4��fW�LS*?[f�b�X�2N�k�B�]V��qR�\Q��1
�� C����b����\^���p���4� �o1m�!2|6m�H�ʪ��KA͂����P3	n�뮇AM�eo�R��û����_��{��C��-��17���*�,NJr�>��k���0�����˚ob���G���P�k����ǟ�mv",[J_����8a�Rƙ?l,��&�m�����5�#��JĠ%�����Y���M�Hܖ�1�d{��G�[��WLIH^p~Y��d()�R9���qT��1GP*�����$��J��"�m���b����ċ���䗲-��}���:/h�~�"���x����U���΂NP!�{��ۙ�v�����bH.�unԬ{��Cy�Z��W��@8M0�����W���8h)����gy�>�;�9@Ƭ����?E�~9��Β��k[��+�H`��W��L�(����\ˈ�F\ɨ�0�;���_��< l�
�F��XQ1�Y��p�p��~�	��Rۦ�T��h�0/�� _*4j�݁�0��{�]Eh,�kR��}��*���y?d�Y�Y��l~�95�.hG�bG�eTt���s	FJ9����O�u�OaR��l��)�op	�G�kdt�%$�i��_d���cm���7��.s�Lb� A}����̓t��T(�Y[������%��Z�(b���#�I,�2�j�x|[O�Ή�&�U�"X����tWA�na
��9��ڡ]vor��Xw���d��C�eVUk�� �|�g�JQ'a��[�?E��ݓk�=��7�<*�Ba�M�|���$}�o/ic4TB���*�*�I~JV��rm���"3���m&q�>�_���0��SV�%�;_�ڣ��ٮ�oI�2c��k� ����*��8�d�e-B� u�]�SSp@7ő���r�÷�T���tR��
=!�ԇ�Un^/*���U����%��6���P�B�VJ�l�Q�� ވ���b7X�ulf ��R>f�4W���:�r��;��(]gz�����_�H�8�*GȨ�� .�z�%m��/\���k�;`^@F+M���5��:Uu�A�p|A_���^])\�#���< �8{��Q�$��w\^v���i�q�̵?R:ñ�A�_I��U;��0���B��Y������s��k�	S`��$��oDĮӨmpDYjd��X�Z_��-qB�h=|�GOx�9�+1�s�0��{׆:Ǔ��G*
e%���D�T*EwO摩XM_ݒ�3�.w_r8�A}��.S��I��{$4�_zڄ��b/��pg	н��"�_7���g}��D~qj�>�e���ܢ��C�T�c).���Ta�.��B�)�����%h5�r���'�Y��Qɓ��Ir���

e�[>�ԫڟ�Vx6O9U�a��ǣ�A9��=�O!x�u��N|M3��7+�8d��?�ىG4S~��4^����Zs��;�;�CĹŻ�lP��]qw�x>ʱ:PV�a�U<)��d	y$V�`L�KBk"��9^	"&,�̓��o�F�!֌~b�u�O����;y�u�I����0�H�`L&��鼭4@�%F�֫/,T�}�(�&U�M-Yy|9,\��$ {1��9G��m�'�3�^��ߌ��l�: �@�Ծ@��a�Zh�h���N��	\�Z�ҜT<�	���xp�r���A	\����om�2�C���G|J/0i�L0����t4�B�Y�6˙���ᬕ,�o���U����H���V��B�#QLOL����R�-������.��P��E�؆�	�f�E�}��K�!��%z��"z�'��vϳOnM�Ͱ�2c�Afg3�/�����́dL��b\�~rE)������գ�zt��������s�HE+��ǭ-e�RYɀ���1��>�3RD�Q���]���0uⲞ*� ��Ƙ��t����	�7��R��|��W@&�����3�Ýj��t`+*D��g#������8^�;�{���K��uw����Q�S����tD��4Wm
�f��k�'R�����\�	li��tX_#�^Ms�ݤ|���^�wa��d��*��~R���[Nǌ����7*i�y4���� ���U.c�1�����[1�E���|I�q�L��'zm��g��s
5J�81dU��cP�X6���#���u�n�Mn2>��࢙@$�ʨ�����&����IT���9riqf$�`'�+��+�IQT��I�8~5��������N�䭍�9��/���K�AI�n�t���t>/u, L�;���4�9��F���ص�wd8�e �)r�tX6�LH�$��oE=�ƙ=@ȶ'X]8T���@��G!����M�1�����Xr@�X���6�Ⱦf���n��i��mĺ�wOl���e�S |iT�A�UM���}��)@6։m
�|ܱ�
j����ŭ#�����I��u�#rmQQ�Y`�;��B#�\�֥��9"YH�������[�Hb�'����ٔ�������Eޕ��aG"�O+�θ�59%�І�FP��{i^?����$� �M������D�X�m�HL���>P�?����_���}>mi5�ˆC�+��*W�$���q���� �y��s!p�_�+��g!�����˰�$���e��F����f��m���|���w?{|�w或�q��>�
��`1��I�>��=h�|�o�^�U���Mi�8����82�y�����J�4�N#h�����KdT�\y���d�`Yw%~te�(f�B!�DH��GI+L��_ωj\�p
���H��O�%LΩ��5��O�.e���23��m64�<�E�:���Ϯ����8a����z`,�3U^7ܩP�6�G��O�3R�.�O�*�-ީ$Z`ܷ�k�����Ki�����!ĭ� ��;C��?8��%'��qn�u9Mq���$�(�o@����҂s���C�k.;ZVL�h���e �17�y�6	G��J��Q���������-祼nG95+3Q��/݌o/Sa�T:J��3��k�����._0���*Rv�[ `�yC8KPr8<���j�p��ef0��m�����/�l��7VWR�R��WP��2w�W����]�~�QX���3���h�"�����[)c�G
�{y�f8�$_��0�U�	4׬8W��_��\DX��ߠ��x�c²�Ca����--_�Zq$<�����G��p���#8I�f��}�\,Gb�M�g&@��GG݂DnXy����|HeUI-���|'d�	�e ���_k���!�+��'���$/���h5$qT�O7;�_�o��eY�<��.u.�cwAfΉ��庪.:�8�R<#O�#�B�T�ZJ�|�eR��d_;������p;���sXi�����K1.x�m�Oԕ�ӀǨ=۾rx"���by5�X�����9������h��)��X��+��>��/|�FLQ
-Х�!/<�����
���_��Q6�;/�+�,B���S��<���G�_�6������"� B�U/��ͦ {[9�ިwf��)��ę`�B9R���:�����,l��b������/r+��T_w�T���^��l'jp73S�k��u�5r��V5W��8�E���,���]��9�g�Y)Q��6N�Jg��%.�Ǖ;gG:�O]w��$�]j1WAiH�n)��ՠ矎+�V&F
�膜	8v��J:p&�Ǐ�EU��R s�7��%�5m��l���z��ݝUB�jx��Je4/6h���	J�i�o=I�=]����5믎���}.��T���(HBv�S�������=�#_�:$�Hʧf��w��-O30Ed����ڝ�c�Ұg��#*a�p�-}��zx��`�D������~c�b�0�
��Л�L �u6(0����
�
�P]��*bF�}��Uyx�d� `���ky���_1 xOC����Ⳉʪ�3u Mvn���؎���dT&�ZAa�ܵ�jl;�9�I�^�@�gy#�g��JH���3=��J-��u/�I���Ȃ��~��@jq�IM��u/e����Q.���O/���q} ��!
^�
0rT]�U�I�J�J�ð��t�r��P�ѵ�Ȭ�ʲ�-R��d����U�]xR" ��kckOH
2����B��Y������S�ݲG+�~_��{"p������S\Q�	��y�17�Ϝ��9HQ��.B
�v��I��{���Ս$:]�,�D7K�����7wp����[i@mo?o�۽�Q��0��N8n=w�7�/RLL/���'�Pk�JFz�t�2�^Cg\f�W~[������@K�4;`i�d�KDy��K�"C�zy�oNts�_1p��p�R_H8fjݿ��ګ��n��@W�;H?�4 
�v��	��W�?�p_?V���lO���XX�3F-�Zo$^{\H��5<*A�]�괼?�z� k{��䙌Q%*�=�\�|D�o��/W@e�j���_y��H�fѿ�G��V}�g^�h��p4��zZ.Ԫ|��PFaM[Ac�����xkS_��n�1=�[��K��7�y��t�!�9ei�л���d�hї�
�˖il+e��~�Y����(�g�3��Фv���>�ٜ��m:��U���L6Y�	K�#3�4ŧN:;��4j��ʾ[z3~���J�T*�2�/?���؛������ߖ�`̨J�ej?ID�
�N)�_�:��)2���=�L;U��u�<x��TA j��y����g	�#�������O�=yj��&��e����}�jZ���#��u��e��(�V��P�Z���V�U�L�2�#%�]�f~�>ux:P��."'ː^->�N/��Z]�Q c��l���x�����Z��!�5w~H�rs}�#s�?s��m��
�#�uӝ	�|�T�G_��o�ٲ-\.�y�����8�6!�:�����J��83�D��ǯ^��}�%�Ba��i_����uS���MH"��bs�E���1�РN圝�%���>�f� cS/t��^-� U�KWp�N:.�#�;��m%�J����&L!*��~�c �AA�d����i��@<n}&�u�]��|�u��<y0��6��A��3�B�7_6����<�ޛ"��5��~�@Hz��y0�XXHHr�_������`�͇�� �[H�dpV�6I���}�O�?U�6�&�?^VcU&�Y����b�	e�xi9Y��M:wOT�$��1/�[)'��vNn�հĪ�3�M�u�ҽ ���9��k�����Z^�~=}��h���7�hsh�A�;�Y^�o�ͫ����ޠ�����!OA;��r8_�$�+N�Hp^��$
��B+$�7��!�Z��ӟߌ��O�9$T�����vW�U�#�[`yP*v�r���5�@�¶�!M���f�U'-���~}��ZRH�a�i���I� �w��S����6�ѧa�@��+�?��Po6tK�m��)p?Ŏ����ތ��x�|ݛ�[�����\ƥ���S�"<�v�,s�4qV�߮#��������((�_�x�n/�����'IZ�@��2uّZ��w9�=��fqb�w2�x����)n�#P�6&�J�}�N!G�D�X�+��C��;0�P��}�xR��۶y}�E�+���}��3J��0����~�s�qPĂ�*6��X��Z?�dI�k:sB�8�-4���v��6���m}ϕ�>k���(F�Iو�SI)�G.R�2�nv�c�S@%��-��]�N�X�<������>�5�aA�1G焷�ד
s���ӻ���;����'h
�c�5�fR.�̆�6�h5;�G;��V4&[���oH?��sg�S0���-i����FXKR���;)���m*V������
6+
;�H��㳶@F�7��#8�s	׋?)���>�qg��4!~�P?H��o�
oJ�z)��Q}RQ�"�R:5��/�Ѕ�8j;���rY5H^����-PZ��g�-�	eMÌ��,�;�5���[�E{p:��$�K<�e��^X��L���a~}hs>J��ѥ�I��T"���K��ҵZ�NY���[B������h�d�?H/��p�� k�kb����R���[[��(.�Jc��ˣ0N�����H$wFr�|J*�>ۨ ��p�P(��l�œ���}�
�Dț��e��LJ�۹�5��َl�����VH
���&D�o��ɐ�R�!]#�Nf�ΉRpJ�)�tw��մ!̴x�5v�GS��$c�ptV��d�,f����G��Hq�|lc�-�<�_�F4M4؎�I�Ko%��6������� ��Iԑa�Ma�,�6�������rɶ����5-�P��>��!J#PQ�)�'�1.a����TLM+�^ %@���
��uth�j{]Y#~�8�Ī���9��a���E�B���R5�O;�Ge�a�Y���
�V��ƧLl�ʇV�hL7R�F�u|�t��ȶ���]��0�ҥ��ި��M.���\�ë~�-cK�w�^8��r�k�����HYD�p��~6��+�ܳ�G%��Z��{�\��pX�H�4�K6O��Wp�_/}��y9�U}Jq/Sy��X�I���R��c�>j�����r����j�f~-��]w�w��x\"%�����f�Q��9[�2��J�C<��X�:��}r�"&;$kq֯�	ݶ�)3��C�KN�R�-ޜ�j�� �犎��Y��%�܉C���[]g�Vy�r��6 aX��Dc���̪Z�ܞ�%�uߞ�������=e"9Ԍ+��3d�fVkT� �U_���es�>��AsmZN�m<�epw`M�	�:�������?��t�2��L6�$�*���r���e��u��A߰=K�7��,_&D�<�ZK�D�
H�����2��B�x}��Ϫ�2����,�%�j����:ÞP|X&W\���J*�h��}l~��)�s&<��
1<�i����V�Ū�R���@���r����I�
�:C��w�a�$��f�L�a��+�������ܿ�VĿֶ_l&�Xzϒs��w��р�y^cLrj6O� \W\�����\�(8�hM��y��y-N�����8 w8������˟����6�H�NčSjV �$?�;�ED�^���.���}%(�� z1�E�����Yq����m,�J��˕��1mHe5�5v4w	�G6!F��{Ė���4�S�͟
8<�(�������{��NiL9ig���jݰ�,wQ~��P���VUr������ ���D�a�ڣ�1�]��+�ɵ{'�C��/`���d�U*8���x>�����}/"���A�Т��Ԩ�{ILd�����2�~n���ׁ
�5����h�k8mp���k����� �HT�dK:�������_�̗�)16����	���T�:��}l��j�	x*
k9����&5IÅ+\�*on]Ms7dI�8v��t���s"�*�'4S�M�BY'�+�?������/S 3�"�[y�)�e���a�Zy��Kd{�n��:�,���B🋕5���b�0C�����Mj�Sce}]Y�$�oS��Y�x�4/T��Z�B��ʘ�5��S�5Tx�.Q�
�p�ґcB33�#�e�����ZDc�dpπ�RԺǁ�^��q���6ΫjŅ�s<�+���fTa٫�]���؈eVQѐ���"���R����W�1,��t׆�d�8ؗ�&s�3Z��{c�ۮ8$��֥�b�3y0�6��W�j ia~����d4�:�^���p���>'������NSl�*z�W��7�br5y
�H��^i�0E� 3	Ϗ�����h�
���z������	X��z��	}QZyӪ��|�������o���X��B�Xg��R%��-�.�I,�'�N�K?��%eU��Z).�K��+��/t��/�}w�1,0�0g���H�Ċi�9���������@)�7F�b0$��`��el�i#8��	q()4&rh�Q�w�Ird[W9A�@�j��&/���M��Ց3��.\ӈo=�@����(ذ+V^�^�M?�:�0�<�T9�X�B��{�.^����!�cP���^�o�m��P���~Br!����b&)�%|E��H�G�7���,�#�]D����� ��{2�ܢF�KN�~��{f�J[Z�'�W�|�X2PL���"�.	3��q�r�)VRQ�Q!���M<�u��ݣ9�U^�����!���Se;����\oI�Z�3��gl�MΣ�����5�:��U2t�^`׺�N$y|rH���$�]=�~]7r�*n2���������=�:*���l rH�֡��2�έ��RSX�F^|�q��+v�ҥọ����3f�~�@U�&9Kq�:��k���������K�4ȸg7|R�:Y4��w��T�L��LN����FJ�=X���t��~�OJ���*���H堻2#y�W�ֵ��b]�Sӎ��Jbh��,�ܝ�X�Wb��������H���<H���*p�n��3�9���F�2L����i��O�6���w�{���E8B�!5w�/��/�(`��l���ߺ𺠘�p��UA�sľ�v��v�S�䌼� �[�$�ܳr�r�9�)a7,��>�>=j��F� 6�x��.^S�.����i��G +�J�!#���Т���ҳ�qގ��yC�o5,��.L�P�T��`�qJ��6���0��PI����Y�1��?si��<g�ak|?E1̈́�vV�Vy!�ܘŢ�,��� ���9�gE�^�=�͂��E]�؎Q���".�	!���,6�V0�Q}�P(�J��	�@e���`t�3)D�I�~��r@���������B�:�����UČ��Z����WG�n?�_W�?��r=$�2�/�"�cs.?�-
��X1�q�Mt�}9ٮ6��&�d�]8l���;�<�`q�	D�� 32*F���E#mj9d�z�c�~F�!����l�}�Q�*��`��^���'oS>h'�	�����#Rc*�&�x�>��ɱ��t�B7�L��@��W�� �:�����/-r����PPIUZ(靻�^oQBn�mB����B&e��+� $�-HbL.���n�S�Rl8��gx� >�8��r��Sx$
��F��b���D�/��p�}#S�&�p�b?!l=�%��!�B�7gHA:jG�����/� ��a��v�� �4����4� �@7�Y�������٠�� ��;�w��j�37���iE�@�Hvr��`�a7ݪ(�Ul�,����S�$������T�*\B��r�t��e���z�Q�d�l���޲�C���1�� �w�O
�a�TeH�t��C$[��hj$�-)ܮ,M�/��B�0�I0�����td<1`���z��_#vo��NK]X@�z�wD����F�C�#���u���җ�;�����.q��Ic��b�*�K���]p��9��!^O5L�\�ݠ���}��j2o�����Ă$>��:��~��`��E�V^H�O�҈/)�=N�;�T,�!���_^<�,>W����!e�p��x����r��&��āte������$���V�����D���'�@�o�8�����{�z9�C3F�Q̛�h{A{A΢�JÎ�m �S���$�5>����'3�E�$YR�b�hE�_�&�#Z�y&>孋�$�/00Gi):���a<��'�2�`f��8dL鄞\}Y,!�Oi���%��Ϧwd�����;q�Z��F����V5]�w͊����Dc����eS�}ξ-�*�fy�_揞������S-菊�n7fbګ��!g�UR����z��Ma�w��"�F�>gd��+=w����{��b[ɴ2�� q������n⒵����U�L�Xi��RD�sB5�GJ�arʨ�wjr�ss*��MVJ%��3a��ݢ&�MJ%X���7�$H��C�KPcPM����2�K�}u�1+�@ �G~�j%3�+�(*®��/�퉨1��%̻|�!���p3ʂ_�bad�eeD� V���i�@�P�D�
>;S��TO��j<�\t�-ue+EC�w��ӧ]���A�bG��*U̍PlF��@'�o��.��b��YQ��Ec��Y�!P���a�\�T!���h���j�cO`�����Kh����u*���� �$��(�.�B��3�g��jU�嬐�%�OT����E�ӄW�Q�^��G�b��G�ZL e�m�e��ǃڽ�r�E��	�Z��1�U��G-��)��/Lm��uj�)�_Y��D�3t#�L'7d��*b�������8;�>�@+�/��l0�"������J�x$����/��瀎�E�%ڢ����R�uGӻ6be����sSA�u�����P�gSj�������$�������8A+�L�Y/��Jk��<&X�	N q,v%�8�X�J���*�M�]X1�%�F�y��X���:H��b&�:�F�����ҹp���6�j�Cc�	�"jF�jÞ����C��՛+��||��^��I���F2�-{�(�r�_ɹ�B�N5=%�!�T5�+̗���u	ң ���O,J-RBB
�o�;�l�|w� 
3;�7*�j1�F�O`�Ph-�
܅���oH���d.���ya��k�S�����F�J@5��u�,M��{�g��u�_B0��h*�gc��]+�Hv@1�"�e��ݻ�7�����W �wEr���E��~�����;[���������D檦�bGE� �lW��',��)4���UJqK�V1}����-�3V���ۭ����i=zY�M�1Ge���s_��i	��
�0��j��e���>а�tm��.9�$���p'�@���w�'��(��1�X���Y��iiL/��9��ϔ&����-�Vx17-b)$�輻O�~��� 	 ��I%�o�M�`��V���[��ݎ��
��a���S�Cxdw՝h�sa[���SΩ�_cF,D�L-����S�*�ܑ�SH�y���j��è�.�P�]b(m�09���K�+#��QO��� ����Q���uu�tzMR�l�����ƃY��� x3ET�0��4�"��3���@�C�n��{�K�8�et�j1����~��-��	�E@ >���S��1����FN{Qj��E\�j��o�$�Ѝf��h����֗
F�؞�����-�{&R�K���r��%�%����
G+1���r��<��>���u���ӹ��0N�iK�$o듣�V/*.�QՖ�Ӛ?�1 �u�.�yP�8i���c!�����{w	_6�h����~�$�T����\&"���u��2{8%�E�F�X���1h���c�Љ�JG���L��#��@���9z���3#���:�Z�F=o�:�b��#tkq(���|���b�����l�ב\+
G��V6e�R*{՞��!�yw�E���m`ƛ8m��� }��dJ[-�Ipm6�-�����>G��2]ǨOXO-��b.��T��ued�,	��_5��f����j��9�4�萘�i�µׂjq
MK�����&��4���;ұ�yp����2E
k������%!c�!KG�آ!'\?->~=�S�᝷���C�Ǻ��/&��N(�ͩc9��a���+�]�+������l�Fl?��*�(!�{�l��{��[B�����>�"Xo峒<�%KVtlv�`a!֑)<jt��PiL|K��3�(4y�V�}
dp����z�m��h�_46X�^u�UY(n d��%nK�.��2�ria'y�4 ���V8���)�ߵ
�#K�H�I�Q�M)���G<7̿��؝��{��k�D_��ҋt�&i4��s��� T�6XU�����ȹTB��\ �7�_���ҭN`l�m	�sӕRT1��D�5¶�Y6�n�pA]�e�K�<X'-3&���r`���C�3��Ժ��� �r�N�;.|�Rk�8�v��l!T�Ɓ֐Ԛ�����X��I~~R\��7�l���m�X��	K�ԛ+v*ۓ��һE���*�Zf�^��2���o&�._�d�Ӟ=��w̯xޘ�R#41XQev����Η��efa�Q�ӤA�f�^���x���y<�"�'������4�Y�F��I'�]�!�B�o|d;�Ǘ�H�����ӊ�!��6I*�(M�Z�E=���F�i����X�ʖUa<����2RD_�z�0X�v�.mW�:��rٗ�e���R�
��?���_���6��6^���|Ltb�qc*,��m-�$�ݡ9p?�l��2��vK]�	؊��UJW�(�n\�3тӂ�cri^p���)�>����j�kV���1�O����^T`?p�f~�2�I3��Q�f)w�y=����N��!/�8�7�w�V�2����M�z9�]��Ǵ�w�C�I.�$�7 �N����@�+�A+��� ��iL�h2`��Wڢn�������[�^`t��PP��r�^꤬I);�]�*����g��g�Q8�|N�1X�陰�پݳ��k�B�]��mη.Pȡ�$�|�7H4I���1��͈F^�K�ប�Z��_�-�<v.��z���V���6�!@nȈ%3�Oә����\�e�A�t&vT*��VX�H�`�Jo
4/t����|�.l	�D�;6�B'�5I{ݙ��An��v�+~����?p�ZP�W`Ar!�ݡ���܀��ާ�<���cLM�(�GgP�m�<�O!��Jٶ����tN���`�ԝ�'��t��Ϣ�A7(`3�=�S��ڞ���S���]68��z��WuUf��B�pF��*�Y�j�!F~���� �9m)X�.eQ@��3�/``���1Ȯ���	���oP��E�5�U������E޽�����΂y�����0��4wT�i7���`с��<EG�lɎm��y��&|�M��QA8��k�w��j��C����Qa3_aa���*�\�s!&utaf۞r�p/G�}�`
��T���G�ƻ%�
��ԣ�Q��!��*��AH�����|���۩Cf�Je�J�>r�A�o�N�"�u}��Y����m9u
�c�Wh�&~I��͸�hxs�7*��{~��o��ҥ��#k�z�y8��덺�Ca��(�j��S'�o!���N?e�������/�x��K���k�Z�S��#1k�s�DdS1� }˙���; �y!}�tH���斛��uT�H#P�2a���Ƌ��do�e����1D�7��$��.Ǥ�h�����ٲ��2K��y�1�8g05A[��M�q�k#X�8����8��V�%�����?�=�1�&���e�a�	�|Ԝ���{������ X/|o`�}H=z�$_b��d� ,$��0���z^�V���O+<��R��֘g��+G1���6�*�J���1yjɭiE�C�x�R.u���.�߯�~y`�r*�I�a�S*:���W���g,�A��l�����c�����'�	�����~8��b�,i]!A糆Β�Xд��]P��s��!D5����!g���e)Dt%�;'1�>��4��)�HzF�������ml����j%�X!���{#���_�m�jSM���`^��bʇ�%�B�p����o��U�Feƈ��2��*���ʌr�V��p��l2���K$3Z��B�ɾ�bz�7k�����Sρ�5ۨ9s4Һ䋌��h.<z�{���=�qe��Ǘ8�֧ȓ�Dd��8�X-�ه�M~���C�M��q�� $��*%�����A��H��-�"�Ge�'z��ȝ�i�T1�k����fǕ���M�E٪�O�
	26;@�jש��_�7�\�`coͽ�Nxg����1Y����V�t4��p�LR�3��bj�1��sg�� ����V��X���l9�8!Lb�v�hr�*�8%_IT-ҁ�J�mn_����o؆)����_�Md��w�Yo���P	�W�����Vږ�y3�zW��5;\x��9TO)R;v)��7��3�\���qo�����Y.6ј���F�V?P*/L��������}g�A�H/Yӻ*2z�Y�G��|a'���h�+���F�n���������i�
t�3E8I*oR�^0�z��+1��s]*q�=��s� �����K!�Qާb�1��0�13�B'��\?AO���u�VO��IC?���z�am��&G��bD�Q�}�I���Բ`,�I��Oͻ�0-|�%$i�W���3�����S60�^�e�;�%�S�LN�I�k�Pw[^p�C�?	�Z����	�Є��~z�}_��x><�Y��'���𶓩j,	s��Q�%�����x�G��]�g���oZ4���rn'Fh6ũX�j��e⿄�C�~���;�u&_p�l�u��/����Ħ`�|�����/��j,�Bц��˶��n�����N��9?]�ϻ �3K/�V����6�9p�����g��]���O,7�R�P��h�4}��C!���?�D���ze�Φ�G�i#�FR�z/�|�ޛ��1sFs���R�n�ee����:χ�4��T9\���Gɸ��{ =�{�!&�0���'"y�/P�u�h��Ӫ��>���W��^��z��q�ȇPY	4ۋ�*��BAWz1߁sAp� �ġA����e�K\�o�����F�%)�#İƏ%ӵ�!}�44�ovYH���@�ym��qUX�`�Ū�rID�я��K������ĒY�v�ֳ��[��.P�e�|:��SlY�e@�V�H����vk��,b�'Ucvt{{�۽^��tbv�z��3����K�
����8�y#�Q�u�[�_g|��j26Aa"��������;!*A�=�X�8q�|!t=pе�\`��Ֆ|<^�ܜ�V��6�Q�ڸ_��+ �� i5�$�k�߉�N`f��Ht;�Ő���j�|�3�ჷ�����ɡ�LOV�g�o�&�]Şk�<dh��;.������<U�EH���ŔY {
ar�;���{�2<%��'밫
��`m�zF�.ǖ���-70R��MX���t�n5���0���U�h�9�n��Y�ݢ�O�z-����}��ܑ�1�T�.���+Q���T2<��N�j7�a���SL���sy�	��(6d>�ź8�e�OT��ב�rC�>�r�!�L�{G$S��I�d
t
�p.IVŬ>X+���&�hŔLK���=�I^�b������ȴ��w;�T47T���A�ۆP�� f��Q ���-���R,�Ws5�rZ�ׅO�k�e�����xU�2�
��$[mrďA���i`;D[ɐ�,k<=��\amS�
�㣣�pۺ�3ex\<4y@���e~�D��Sa�Ry|1W�^`�$@�~&�ɨ��3h�#���N��Nj�}�%Nl��"<S&w��i>�s��,�m��R��#�ҋ�g�u	��R:p��n�f�^x�hC��X=�#WG�Y�����\���fu��
e��:��y��yo�Q��.ֳ@���˷�]��6(1�w���x$s��J)Y�;ݾTl{ϋ�Ъ��k��3��6���j���+0��t��BVBe��d�߬�M�>��kR=.Z����wh��^��������6C�,��׾w�"�I?"�4��^�f�(4�W�A�6!8j��p ��Q_Cd!&�#�4! <��5��$.~��%�6�4�DЅ��a�7C?������L<|���+�,?rG����`�\��z��3+��1�Eƪ��G�<h��S��L�c��[�8�����β`�E��%��k�����ǻ�v��tcg4W�
���O�"�g�נ�R�ok�M)��~��9j�ZT�$�uj���;(I`��O�;JVs�{���{��ڠR��8�*��7��-x��czfU����+�`�����I��v��K�ĵ�-`{{��}l)��6�C�6�֧ѿ$w����S ��w����0�m�2���-޿G�+��֚�e��W�����'(�'q��<�9{C����WM�LO������A=�5R��Qt�B{�3��]� ����E#fgk��Y�zUL��-b��M��A�䊔�B5#hd+�%H�f�%X[zr��n���E�'v����\�p�5k �b�ej�0�TJ�%<�5�1^�؛N��U��['r�Bj ��}Oq���p;�G���	�X�ۡ>]��=_x��`_^�,>�#�B��O]�Y|�����ls��C?��?�ڑ���g6z���9���s��MpH��c��L���G��D�����0�ɉ���Nͅ��_�8|nx �FI�al���J�1}>�Z���}V�] �6ܚ�ƌ�����'`�M"���2+�i��l$�h@����q6l�2D����3{2+`�[�o��=*��Q�D� =Я���`b;P���pb�=�v4KJ�l}1p��I���lQ>�x�h��F3�W���깓g)@ω���uש3��qH'v;�T=�Bu������T}��h�aϐ��^��R�@��E���.��9�sR0��JF	A��s�$�q�R�lK�@_���B�a�7[ޖT���I}S��&���ER�&IL����pJ�.k��)j���>C6X�G�H��9�L�W�%5M�UDPn��!�FU��ɺe�fc�2׾D�an����S��4��q����F�ꁡ�IL��>��s�(�Eb)�n�p��y='�K����6K��(�m��Z��"����UZ߆L	ZMƿHz��de�ν��|&-�=�@��T��ّm\ ����p��4���I��K��v��M>��e���Ȃzl�~� �Ě���k({"~�Sf;
w���2��Ľ�mǂ13����Z��;qgɗi���-W3�6y4��G�p��(.��8�t�b��{+xm��Wvtb�w�AI�L)GD[N��.ݠ3>$�$��=�n�p�-�Y}u��;0J� Jmt�|1�U!�E~��U���'>�a֊H�-Z?�J��(]���=��G���$�$jb!����k��������=���N�{��pIp��:��<���m�s��M��5!C����@�L��ɩM��{����Gǔ�������΋϶0��eo�q����h���jm�t5q��<���K3�:�an �O!Q�x�K^��0�)����q��ܮ~����]
ja\���޶����> ��+�OY&���J���,��D����̗�ʮ��e�M���s�����/�����a�[�+唏.�<h'����4��{�������3�@)��t2A쩤b�TiA/������n,dM\=w��Ck~ ,b��ų>�M�]R��n�,{R�����#����!��)͍U� ��V�6~��/��"�_�ӽ�y|����w48����Ǫ��j���^LYT�7J��P6��NMf��zuL�@���m)�u�-�Wb*�e�4+�N�?��Mde��n=�0�<�%��DY�s%��v����:�6CB!���hI�K�W�4��{�ߖ庒n��J�:_a�Ș_��R;��j�ӳM��;J���A�[5ykW�)��i�B���>����X����&Yձ=���)vi�y�'�F�I��K���HQ�Ch�tJDm�O������f�\L���6�L������8�E���@A�l�8u���z=(�u<��ǡ��)���5�j/G,BO��B�g��)��XE]�~9���W�Jyw�q�i�	M�h��������VJ�C�zWr��_�]y��1��x�pD`��i5��k&̛�7��f���y� ���3��x3����>b��.�R�z	h�rp�^�Y��P���\]�+Gx&�]�K�:H�����.bB��1P��S�{j�F�LP�RZ��{Z6C�J���C�Ո�Z�M%�.����/?F	[�h>��D�O}�X���1CB������MB5�M�y�f���%���d�x�4�YF�m���8 �����L�W������.dR��%����JgQ/Ibx0�Q/p2���Q�	Q�+~�5DŹ�!�j�P�Ȥf�hdd�(�m��|����#������2�`��0����$�2����n�7&�XZ NûC�
d9�FJro��RU�~��\��)���_�R�,�{�P����>�o`� ��$(c�R){������9�./�j��π�}��#������/�I���2K	 hh�d�dX�)�\��%T�N)�T�������uN�b΂�&i��X�H��w]@�t�rW�D��8;�f�X"��H�R-��).eȢ})�#����r�#c"M��. �����sm��Y,��t{[���P����2?�^��GK�ЗY�Vo�Ɩ� �#���rm*��sdX����A�	������������.V��!�/!#��/���a���"/���y֔�~���̸To��'�*i�.ɰ���fu���v]�ۭb��33T���	Ū�
�ɖ���K��qU�njfIX�۾ ���y;�	��gwHWZVCJu�D���_0b�c6�]\M5��u��ԯiz~���қn��`jS���}����@)9"&+z1����<�.�S�0�rt�{�_�ޔ�?�пK��j�f�]�O��c	x!��W�O2r�2�&U�7Q����*l�0�_$�� f�������W��m��{j	Zk4c8s�i��yL+��l�,�v��tt���/a���4�. Ū�·���RE�<dħ�T�����;A
�A���X�YiX�$��i��n����o�l1���']H��,�Pيjz�و��w�,j�Mx�X=m���=F���*�@DF�V'����-���26�W�e��x����� ��i�ށqď�E�N1o<7��v����V;���bgв������O?�q�	W9�k~(z�*L7!����}�Sn�S���� ���I�
���z��#�����^h�:�q��i�6Mϩ\�����v���0���������a��G���bO�)��,���Ix�	�3����$�n�-�:��P���1ې��̦5Ӵ�dx�G]M,j�m!��C�3<̜���c��}�	E���e�p@���d�afo�G1�����{���`���wg`N9�ſo���וN5rwE�_\��ZQj����2Ģ9`�,�r�d�.��D'�ƥR�%��hA����)�v�Ş���-?���6���A����K��]����v����n�Y��s�ꥠ�Zj؇{�ybJ�����ߔ���TV��=4����J+c��RT�K?���G�Q1%,L�FE��h�ڧ�F6D����Q����>���=�65�GݏE���m9x�� �r��N��u
E�I��p�S[E�&tn543b�D��#8���v}�Lk�(3M�O��@��
-��6��G�g�.`uF��4�=�i<�����5v�[
�rw�DA�I���CB����4J���ד�'%��Jf�7M~�~&�/y�o���, �����0z��?lbXG ��0�0����h����_h>�5F�\�i�"��D[�6�
ĜEWU�]�E�Ri�(a�@����u�X2��:���oB�0�Y.ko�ێ�K��\��N�� h����c_�9������Yu'¤㶿{�w<7#FHT�,�dy� ��'�o���6�6IKꑇ8hBsS5|A: f�|}���f��bT{\�0�r����X���7L96Ǯ�ċ@��o�K��ɴͼq�a���Wpkև�-�j�'�h�b���hT�=v	|�����|g��ȹO�<���x�3KӘ7Ω�z�Df��;Ԙ�M���2�͐?�YR"-싯�x.V^}��]��M
��
��!�"n}��о;P1�Y�hw�_G�<�{C�s�^	�����V�U3���b���f��Q=<�K���4o*3Zd��������?�ͬW>�"�����V�߭��g�Y]����k?�i���&:��w�{���yܽ���b;{J��b�6_X�Ima�Z�!���\kH1�'�Y�7�V�$hK\�;m�Y=r�
�Lb'�4/��[���<(] h7��D��9��K-r�+�6���e��\܅�Zcw>��w��1[�+K����r��K�x�=33�Vz3W��w�h�"P-�7˽W��U����]���e�g�ʶ��,u�Z�E���M?�x� X
oB �v-Av���ñ�VK}u�!�Ä䖜�=��� ]��[���s�3��m���a�>'���<��#��PBHe5�R��+����e�7�}�H��kO�NW�qq�U~B��B���c4�����x {���?&�3�:���[����"S5/�Q����ddf[��}�nB�'D��	�l�-ve��6�:�a�#��,b=#�'�us7������?E�_���P�D]���1.)t�h��y
�ǒ0[�y//V��pU�T!l�`��'��X������u"j�|%j����$�[��|�	��!�`��p�C'N�C��ƴ��ς��|eGKE_�ZX1�E:�
� Ժ�r���N�L4�5&��X2 B�b��%j�%Y�<��bi4��I�"(B�J�〸:��hG(;� �����[0�a5ua>�Nr	��TzՈ���^�mrGo�^z-o?A���D9�� ���ϡ*�D�d�æBi�M�4��o\D��	��$xt/��Z��	2��yvM~��[�ʣ%e�+�����9�����`�3�a�*���qk��ϨD��p��)� ��3T^Ȅ�@2��z��Z��R�4j[��d?�\0�����zk����{���_��F�����P-n�[�ϋ�BIm��C��� f_�2�b�� I ?����G�|�l����1�����X����*Nf���S��!'��������K<Rh�X��=v_���x�g���FUҔ�/�Bī���mg�ۧB)K���^��GQ��Z�����,d�z#��)[2����645U��Ź.�8�hǓ��)�M��zR��vZ�_ݵ!���bsm)}��1�����A6��f_�W�R�xM��������O��p'T��͹����Ł��}�.�J;���ͣE��'�َT��*�HvI�� �(�2<w�V��v����SK ��`���/��};�b^L��������}�V�]��6d�j�y�p��Ɨ��� ��D��]�T.Z�j�������ՠ��禾e<�)��qS�f��9�!sړr�U�~��|Ҭ3w�у�RY�"�v���NB��W��p�#%���й!���/M�A��g[HF��m������@��<Et�Zt8ip��Y.(J���F�@9�V������Rh�e��U2�ݠ�U#g҅s��_o�Mm?_iG����!�k�eq�%�m��߳!̛�4X,�0ǟ1��PL$E�	ڒ��Va���)Brw�繭^��p��R�]�pZb�7S���"��Ju<z6
�S:���b!��v�/����8�}7�0��(P�����~SS[*�MUH���-@�<�("�^�(�_�C��I�Vw�Ԃ�@��A��v�Ε^c�B�ͣ�C�S}��d��
�.�x���֯���6�J���[�n�!J ��Q�)�@b!q�(H�o�q����6g��S.Ğǅ��ph����Y������@³>�Z�uq�Y;�O�D��O@�*3R��Mnռ���=�Q�4��7h��[(�uw�,*~''�m��	͞�;B2�B�-`oAK�֟�S��Ci�rJO��/���a��: j��:��,�;�d��vEK���Tb�񃃆�t���(Y8����R�|�j���x-#n�9X��x��T"��$�ͪQ������z�����?�]�z0V�K�t���a�r�Kb�.�7�rm�Qͬ�A`�0��#�؏,�a��|<���H��H�f؝8H�Ǌ������-b���@���e`6�l�9*F_��	(��'��RĐ��Xl�$$��Ly;�5c���^8f��I{��gkf���nk�؎�~�*/g|�Ѽ4��	VU}���Ɍ~���H��?O065��*='�i���<1(Ko����i\��zicC�3�fe���b|���L�}ZPR��?���S0-��w�*aϙ~�F���[m�	���1���B����/����>`�Q/ؔ6>��z�ßZneǲ��������Q�a.,ֵ�Ki�:�[�qh���WQ߼3fxC�b�@m̔s��o(U����6*0��*�t�=4y@������C&���<x05�ؖ$����~�K��o:��0��\��T��OQy����A�T��=��!(seK������RPFh\棭�Cv:��5�f�s�r-�_�@r���2g�c���oD��	�m�2R�u��P[��^��S��q�=>!L��#��uJ���(���O
�f<�උ.��b�)p�ԯq�1u�h���ꛑ�Wo��e]:zܚ��KC�N8{�q}�,S��ˎ��V�L�9�%��*�򋛭�Dn�7j��(�ǒ��$ڗ��.�qfےе|���XE�ˬ׍I�;_����zV֏�.4�iu�-��w;kl�V���Fm��&������tXt\���~Q�_�я�8�]�ጋR��?Z���[,��G�w�\����q�����+C)��H����@���^�׌J7���;T�X+��x�6̘K��*'�8V?	�zbu|ZX�2���elBÀ9b��ޗ����I��Wc�Qt.��N(���tL-��w7�+9�
{!�+���AeO�6����gn�����Q�eqO(�$�G�ih�_5{�*K��X�c}u��ƭūT����6C�1��44UJ��;�QS#s�b%��S����6��^�:�x*�{�s���bT%�A׽�et{P�_��lKQ$�m?ɇD�G�ɷ)�"|$��2$.�p0�W�!�JR��B��o��;b��)8&���ҩ68w'�5�Uj�v.���p���J�@�/@�1�^	�7�l	��O�\_�Y�r��/:J6�����*F���|L���^��0��0����6Ǉ*OR�2z<��7��<K�c���p� ?Űn�ك3i��� |4�w"�D,ک��Ə0�5 O\���.��;S8�g`b����x|���\&�&9��r�'n�P%��*��=�8�m�|�8r<gX�CMw_:g43�+�ɺ��"��9WMQ2�L��n/d���O����\<��Y��j@��}�.��Hê���OA�Y�J;�W�s���e���i�ύS��F7L��H���lRh���G�X�Z{�� ʍ�	y�#����xp�{�t�ǵ�M�U����"9��S6C�7�媢�^��E����f���7�f�X^�̻3	?��S(�m�i���Q�{�1?��'|nu��t9Ő�<�ʓJ�ϫ�����Rj�fg�'/��J:���Y����3.W ��K쇗)� ��fsPI9Z��)|,�7��L86\���$a�,<a�de���z`©Z�_(�V�]�jϹg� �L���q_v��4�Xcz��Y▗�H����`�Z"���n����ow���#s*�_�W��.ŃAq_oVA���>uqkPI4�3�_��,+��=ۣ�C�
;,��\���8�s����-�T�3��ǖ�q>�illۯ���hOOB����9k�����+1�ː��� U%'�l�a��+}�����ݽ��285�����⣅��#��]� �m֕uX�~5�?`'UF0�
S��F1��3مHsbVY��א�tS���k�)Kk�#�}j��2�����3�kߖ*�8�o���8��A"���1�҂xy��%��c�L߮��63@�J�8�߀������ꀵ/�8����_.����@É9JUw��D�9]xɠ�3��GSc��K��] �NU���'�`^���C�8wo_-�L�Ξ�U'�)��2���I���:�?�	*'|��Wj��XD�L��z��,/��N����!;Fż���hj�ro�3����ϗ�w���T�h\�ɗ}�s��ҫ���2��9�pd�gì���e!��Í�q�<E����d�2 Ckf�m����{�ϕ�� �aMk��K�i;&(!G|���q�|lE�x	���;��H$%���h��1v����̹��I��.�[���_;�
�0�z��D�e�3���0�"*��y`�p����t��������EcQ�+y�j��(iplUz�踇���ZF�,��YsJ&�7�Q)����9�.�%=��
�r��խ�m�	�B��μ��W���
c��ey�o����^�0�?A`�����H�n����YYd��m�3���?����X��������l�A�2���-�#�������og�^u�>q���u8��u�PD�	dz�%�s�]�]d���$�ζ��7c�J����Z1��^T�g�`?z,���;�%oZ����z�9!�4��U�����(
���#�r�GsA�$��� �D�l�ߤ~��5Jh3{��ӟ��"�5���PU	��&d�e�u ��u�L4�\��kZ��"'J��ig"jAJU�k���X*��I��57��iwj)�V��m@�F��H�~�cW�if�ps-�U�;2$џ��p[`p1c� ��E4T��X�ih[���g!0_o��?�Ϋ	e�`��?�Ϣ�)H�&�VsOs�i�9ŝ��)9��ى�[�k��w�)\�b��3e�黴s� ��Gd�G\�� ���3?����ez���>+����E�a7|�.!w����[�,?"��fR�\�n��|�/��R��J�\;�����C�+9���q6���W=.�>܌D��:[�F����L�n�Z_����	� v�sy���	l@3",��UPSj'�A��Щ�f����f+R�>>)�Pt�E����_c��y���N�m���*��B2��I��E�?��1(6���F-��s��](���)�"<U�,�E%\���ؙ%��gF��A~�6� f����Z�R*��	u�&����Gr��ӑS��I�:��E�;���Lf�f%M��e���<9}�1��!�/O<��fe������%�O:n�8ȓH��Fq^ܜ��ɕVÏ,���TT�P�D:��n�F�L��b!�X��{ �'C����ީ����pK�ZQ
����!�$�����ѭ�r����tI��±�⸢��]��Դ��o}﮿/��-�]]�G���s���s�����*;u,>5���d6��9@ᛮ}xڐ��q��&��լ~���%xهs�x��88�Ÿ��;.D��#m��t/}��
�5�|U��6��sI<?-PX���M�0qa8�)�|Td�-Z�?b�\
nD����-�U����ko���]�9i;ЯQ����cTQ;���Ϗ�Ѭ�I�Mf����H����A\�j����qU�%���>S��#"��;�}�*��̨LX�\*�M�&�� _�BI�M�ʴ�eU�<��^D//K��j�Z��A��3Y���Ф�����s8|K$'D�~ސ����T��:TI����F�L�gU)��zH�0aӐ��g�飑b��1U�W6R��&��@�n��Ѽ����[m���K�K�ng�����*�2eU������+iX=��r��y��0�h\X�D���A��3%���g?���x���7���'����N�If�񑰻 ��g�7�'����ކ�h� ��@�8������uO�!�#��V��Sj4(S$H$��SM$q����'�Д�WS_	>z��T!&팟�~��Q��@��н�9z�㨕�?^ا����*�5A�GwW�K��V(�&�g�`��􋨡g��%$���Im�	�$n��%v�5Il��n�#A0p�����,��e����w��T2��J���B���f�͒���)~��>�&`�r6�
�EsK�G��خ�L�}�Տ��f#'�{���xW]_��6|�|I�����0U�g{� V���ܐAɡqWP{dp�7��"�f�)u�'+��6����c���S�\���)H�ᙷ��4�;=���&�x&!t~�MXL�����O��9�:S7.-�yB`�<��>�����V�l���|>.J ��yhoR,	>�縒3�[��/�cO���,%no���B tl[[#�#ٟ�z�����d7(B���R��ƽ�YO�]�8$�?z�KQ$�F�˶K���Eg_2Z3͙��s^�����RC�JI��8��$�5��ٟ1��GkH���*st���Y?����Bq6���wK�7a��`��?�VSt*KIyp�u���nG��uNx^a$�:[v-�>O)�$'�ؐ%�N�����	�!�wm�F���+���׳���J4n �R����,���j^�6�(�#��1;,�G�p$"�Η&�G�N���9��Șɷ��f���#@Rj9Dm�ќ��;�sI�9�F�w�
@K��0�V�O�CB�䂙�8{��	�����t��ɞe�k�Yp��A�?U|&�h����3����Z��Ɨ���fS�GOe��wj1�҂�J�ǫ'�VH�/���5ƒ���X׿cn\��w����<�u �a���+-�cEk�����YQ���P��#Ϧ���;P#F���*1
����t8�o׾�0�z�`W3~���X�~�
[�~�L��s~5�Cԓ�����.��������?�ƙJ���hDC��R��ӕ����E�[4�s��f�Ge����.�$%1�WW1��P�D�:�����л(�ؒ���&N=�����d�S�*gB0�W~(~��Nb��2�o]�40Ѥ��ҿq&D͡F���&L�f����܎�&*������{�V&��_��b��贇\�ƴ猄��r�9�a��(;N[�������~dS9J�ݟ�؆]v�->�����B91/D��h?^ԟ�y��L�ȕ�FwU%�������ײm\}}$l�u6X�}b��0�k��cqrsg\��z�w��3��ˋ�J�l��C�ܿCj�E��)21ؕع��lK��J�B#�����	a�g�J� �ѻ�^��ö����Ջ�0�J������' F�7x�0�C ^�]���J���3�פ�w�vBH|/���|���'�c?�[;�(���?�A @��w����}��́m��>���?�U16�7=��%��u��,�>�X܆��n
��by9��w�qH==f���~��c��x
X��v��T����C��,�%z���'|r�7�����$�j��X�d�s�l��5�����L�[�OT�>3�͢��-��q��`�˲�*
�y먭�ΐ�i XCY�p	?��?.�n\���7v��Vɫ'Ϣ�]�,� �;�^;�0�	!��Fs�	��~��U��l��W���릦.P��_B�gȗ�	^RH��W�4��j7�H<���8}�����X���$�+�S{T[� �A���2gu�;ث��&��Ai��~�ĺ녮�Z�[U�շ"�8ޛ�n���y����g�Y�;�f{�2a���B�ȿ�C^p�����x��R(W{���V�f�q\dn�5�4�0��"�/Q�@qw��P�C����������0E��{�?��|0�Ox�R{��/$�5�k���#�YQEjk�62�Ч&��A�xxu~�Q�ԳK�����m��r����q&Dc�PT���\~�} �����v4���+1�em+-�NL�b$mԋ���c@0jΟJɥ�rvo��[�g\x��D��I��p�[�LOnOI�F���Ao��S�͊�<e��o��V�+��é�C<e��h����F�TZsΗ��6����OC�Gq������6_R��q�^
o�C������ut&Fg'F�������D�AL�.��=N�6��4���P^�/7`*��\�]�j��F���G�ŝ�s�
�V�,�D��T��]�_l���Uת���I���m���EX�_l''u-��׼2Eb�*��^�ȏ`@1�{��܌ƃ�.I�� :��)֎g[JFr}M�U4��V]�2,��5?�*��H`l�+r���}�$x��%�w�x'�_R��b���|ܼ�ߞ�i��u���A#lƆ0�^�{�H��[$.����n�P�?ޛ1���=�q�8�x<Wl�Nt��h�4;{4���}e���X�_��|D=aV��%2�����&R2����q�M�Z����^{@�Qk@�!�ulɪ��wp�+_������U8��,b�w�v.T4̜�w/8c�|����
�Z�n��[�t������٘���V���|hƭ˛����8ͭ7kg���S�j5�Mf���lR�;��[
��\ŇI�ܡ�m����î/fh���Ў0=N0�,bd��.��}l"K4�J�54,P��p��"�)���$�9n��T�g6҈D+���AS^���
�~�)=`���d�v�=^CCI�/�;U���%-�AwM��㸪�����.B|�OMZ�v'�� ��j{?\1w�{��@RQ9�э�����0Z���@���$��,�jM�qeY�(��c]l�ww�@��m�Ȟ��ʯp_�L!&�{�;	Ґb̢(���߁��->�^�e�B�ʑP�f�:�O�הM�T��A�iQӟ��\�q���N=d�y�i3?T����e�!05�t����*S_�/�c(�nK� �������d�4D��#h���|b"�qX�z-�/���)}�ب���3I�$"�Q�z�xɌ���*-��2|<��$���aEm\"^$�y4�t�a�ȭhw�$'�=�t��Pkc�]'��3oT�@���,�2D����1��'�&i�]vT"�jH�L���W�<���w4
ףּ�?���Ueo��<	\N6�%*i��=��]�r	+&�Ϧ?v�:���rNԭ\�0o�S5�@f��j�̤P}d'�%U��Sʩ*�kP���^�R�v����5�����
��4�7����)���R����C:�m�Ζ�F��
�_�h� eXC�H�D��8���S2;�8;����V�:���i�n��\�e?1��hJ7e�m7��R��+��H��ˊOE��b��8���$�5���!*���f�.;ʃ�[�)�đ#_��Pg|#�2]x)�|c����K�p�qQ��>��G4��ӵ ������<cq�q�!{P����m/*9��nVd!+ȋ���e��AyV�t>�phl�p�h$7ph�4@ȞEZ�2��N�ʋM�N�0@��'*����'��BH}$�#����e�IK��`�d}�qŶ,X�[V���w��9zu&�y��>%!7I��}�œ
4E+�xNu3�5�Zf.S�h�SR�¤X�D.W0�BR��v�\F*V�T��ϥ����5�E�+�źR�����Q�U"��<R,���쨓�T�Ie����yz�A�����`8!�D��@w`aX�X�f+����R:Ŋ��ĬZ4hY���/��Q��K�����Dh�捴��V[/�jb\CR�X�e"��7sԶC�7�+�����?��XFA�qϾ�>��`z��|)&����*ȿ� ����W�����/!ң9��ВIV�i��Y�s|�R-��+bfr� ���@rb�$Fv(z�����a�oa��:t��աCdR .��[�FCQG��/��g	m���iJ��Y��sl�⇞+�
�w���5c���R��+�MOj���P�Z����d�mDW� �����=�y�V�M�g7S�w:ц/=�R��D�V�v��
�\����@��ذz����(������?x�{d �� JrX�B=1h���8��m�+I�O\w�wޤ�Ѯ�mZO4���À���{���J^��a�#���,bf�Y7�,`�7ML���j���8@j 	��je\�#W�� ��AH���[�%��}[}m3�B�6^/:�Q�)�Ԛ�
/t$-���B�����B��^�g +@�[IeTc��|G��M��.a��!�?k����#y���@�͏��b��4���mfD�KZS:�m�4�B��K�v�h��_>��C2�f�T�)U5ru�M�B)޽�Jq�}C�6����ZeF5M���N������k%wG S5���P�����cA����䃫������]���|즔�U�w���N[��B&ʨ	/L�R3Pk|fh�~�Fy"����9�eV��h���Cn:;�!j����s,%'N��{��W�2
���|��N�:�U.�_�|���i)*E?0 ��T�g�C�i�>ƅ ��'랇2�䒧a"-u;��lh�|֘z�7fJ�R�����g��]9FRvx6�e�� '�,2tQ�
��Q����#ݮ�O_�&@���_wށ�9�#~aѕj��-��J��h�r��w��F���sl�~$���.v�&��f~Q,��V��Alju'=�������sf��qE�F��-����[���H��P��q���Sn�I�miL{uފv~y����Fy�,mkzJ,��:46��#�bZ�j�F�c�Ke��>�a%-���Wd�����
�)$���?����F�ƥ#�w{/x%�=�C\�x�-{ئ��ћXj7�e*�j��ܿ`ڇ��"x'�q �Q�a�Jxe�S���O(�5A~rm� �0���(�����c�?�Yˡ�-����6Z����3�$�x�?�M`���� �1��o̓RL�p}��ɐ�(;�]��60�3dǧ(:�zF�Q����U�,c|UOw|E�� ���m�G=�aݒ�q�%񺅱9@�v
4�<{�[?�ǧ}ޱ��f���K6��í	9�[YW���Q4&��?��T/��@>�?*87nw)+9(O]?w�b*p���h���o8Sör�tA88ަg�(v%�ת��#=�=��J"
qگ������㦅xN/=EHajv�Bʞ�қ��2�E
�} ��b����G)�Z�S>S{��ݗ��q'97�׵��3r�Y��T����<���-�h}���W#R��!g�3hw�eu�T"sJMP�����������m�9�ױ�G����׹��)�g־�;��d�sykd�#��D���&U}c9��H�:w	�-����u��-������E\��W�<�l��sj;��a�?���-!����!0MO	ڂv2�8F�߷���Ҡ��zĢ��R�:�)�~K��,�\ a+�K�I1� ΋��K�Y����R�-l�%�֓-I[f���}�r�q��8 ����^k��[�N>��h�7Y�´���]����˸�~1���W�]?Y�r��F>p�� P�4 ��Fq��fn��_�F������(ؤ:�fz2"*�����3c-�X���h��<�䥋3�Cw� [��b�F(0P��Z�V!&&_��=E+��;|wjK/��p8��#=SbE7(�ۋ��Z�0?�Md�rg���s���y;��5�E����f!��5���JbK�Y ��,@p%�k��N�����v�2#Q��R�覿n���wV&xøuδ7���ڛ��^��K�[MJB�)嗩��9�<HE���$	B�,���B�R�K(����+�w���rV@��~�1�ĉ=V9�\�4Pw��:��I[�lK �2��f3�q;�ѿ�(������}����G)ϔ*8��(O*�g��1iM�S��N�����!�k>b���N�`|�+\E�-E�>��W��;��"j�Ѧ�#Ϳ[�n���Q	�͵�� ݸ�3N�(^�%���Յ�s������L���{�;艹�!8[���m}0���^�z���
�>��{�#����)�!�Z%������Nk�T�V�mi��ɦ�+�I��d#�(Z�̥���oj��a�1�N ��{͓���C������ay�n��l��4[��G�=7��yf�gi��C�,��I����(�oP����dV����ڃQ�����\0+Cs+C��Y��O�*��;�s��?]�rr�O(�,,�Z��Ƹ�>PC8��%zc)��&�4����tb�Z2�z�["T,f>��'Ӹ��-~�%5��y{M�|�6��=iң��o��2��sy�X�c�%Q��M�~�i见���@�9G,�G8R�g�G�z�V��Q	۵�	=�U�_.h�ؒv둕u��>�O��~{��9
g�F���H?��,�
Q`�!��<�PS"�Wk:�����̵�
��#��ֆh�P��:ܚ����̩JĶ��t��)"�3�\��hR9<)�,�58h�]��R����I����8L��I�3��U�C��B���{ �vV�r�sט��l�}���8;"l����\@�p����GƥB(k9�6��܋�^3^�tW��c64~�}MŽm�Mng�]v��]����9;?-b	�����]����(��g��9$ݑl�&��g��F,2� 8�{�η�<W��������ι�^ ��Da�TuM6k����n;��&��N��0��ӳꮤMm�>k��8B ��8lF<.S���K�B��dZ?��r���n<�V�cղ�;�Q���X����,@ ��<��X�*�=�A�C\3���׳HN���9��4&C�F~:��T�5ω��x��*+Y��g�ׄ�����e���V��"b�`�:O��"� �v��0��BX޲G�EF��<n�k��+O�8��
>�
�[v|_=A��z8�k����?B���u7��;x�(�?��D*���JR��F��YۃX�F/>k�$6N4���y7��+�
���\�]h���J�=֣k)�����Z�i�7�㽲dC���N�p	ꆄv ԣ��a���$���~?�I���r⫝���4^�}8X���(�z�=�L��􆜷YgT���-^����� ��R,)�
�{�"���bN�Sy�h���N�+����%>�����{�{����R֭F��3�D�?�ƞ�t_Y�����c�\�y|t�?�[5-��]H�+��(��,�o�ܨ����9���� ��f6@U�2C&݅̒+����Kf��c����C?N��vicsa�<O�V�X����9/�|5��~�Θh~$�"�s}]�e�X����	#��,���ua翧˻}�A��?/1����5#e�fk_���?ӝp�R�\�֧���{�:�˲t�y����Y&R�����f���`����P?�����clyk"kYh��+�⬢�
��^r#���ӷG��.�d	���ޭ(��OGC~p�Z���a�9�@�����6
�O�6=�E�~as�pC�+�-4�	�ȵdRX�rL�0�(BM��]*�֤����_j�j�:\] ���&����N�@���4m�=D�4���Zz�s\/M�4Is5�1Y3��-y^���J�[�O�sgcu��g�q:��x�[C��=,��qî=�
�B�}�X���kf�E�����;@xH�b��tf��B�egK���;Y.��S�����o�X�|Yb�U�~j;�l���J7z%:]�U;7e��cR��Mx��d��"�x��e�p�t;-� �p��&��+�	��#��r����eE�Sɶ�����ɣ�?"@K�"����t��� �nF 4U����4YV[NZ��Fo�%ƢGp�
����ڽ�;�
� K"�V���
��X��:��4�*����@�W6��(7������)q��z���5�n��A6d'#�Q�0�_��
0d�f��fR+�qd���p��ٳ�u�@TL
�3H�F�x��SE��� �\���f��Zi�a&�or�����Ƭ���.0K�[��WG�I���n����+�\9G��Zȥ�۽�}�����2����Bo�7���yjw9o;�\��f�� ��n~���`�xX�F��v�p�P1,�e�&~�d�Fn��S4�����ѧD���EE(�_B^k��}Z!�ŧ����`���ZH�v"qY[�R���h�����F����=]Z���(� g�,E 6�'��P��P���<숱��@�v�	t�M��O�r驇��hu�`�\9x��Uo?2�ן���Ӿq<�ğ���W(ɠ�mU�D��a{�p�g޺f���?�T#�Q�iL��vi���9������[�:)0Ƴs�G��(|<�H���U���z#�7�)�Ԃ5�,�`�
N�v#0׹���EE�Bnn�uXG��`�w|aV�����֚��]}+�Yk\o9����(d�����o���� ��^��a4�q�Ʀ�͔���2��i���&���?y1�+�+Ĉ�
I��^xϙ��C:A�G�^�]�Yew�d	�(
(�3����Hsd�U��賁�f<+5㐄xg<��1�2VKwgE4/�2��X1��g՞$�A%QC�&�T�>ɤ�>O@Y�v7B"D`%Ek9{b�Ǖ���"�dO�g�؆8�/��sL����y�$SI����R�ϓ��M8���i���FJ�"��j��ῦ�����ֶgb��Z+�CiޫyX�AS%����f�7�$���a���p�Z/�����AR��ˆ�+4��Z���~Q;�=� 1d��Jd����%�W+Up���#���K�e�42#B\d	��z7�H��F:��<ˊ}5��l�=k��gVk�rҪ����-wd}*��H�1�����T����!�c���5�E�Λ����@�PÁ�m�jR<�RӞ0!��$����]�Z��X�3"����
��7���m���g�-�`px��V���?�V��F�F��%��V��cR�J��i$��D�t�{��z�,2�ĳ���G~�����	��R�����ayWKZc��K-.��P�^F�xA�4(r�(}-�ݶ4�5�Wj沴��}�U�$��iƘ��ׅ_���&��� �x.8F7i�cŰnc�U�m{�m�c����y+�=���g�M�c�h��ǈ-�T��e�Bdɇ�c��'�q�v�_ _�rO'ˈ�3������\��)I=�'�J"�����&עai���(])�鹎=�8jXJ�J_�ǲ+�͸u��\̭*���f-N��r��U��
�/���.Kb���p�����a;����1����.�S;�),y7����Rz����j��A�mH���Q�M�xozu��Xƻ��Lg4�"�w�>ɘ��zD0�����瑰�[e��	�6�	�=�&�Ls�Ԑ���S�{*�?6.d�~u�T#n���Z�({�,��Ft=]��Dq����K�t�e��W{~�
K^mA �@7!شka�?*T$�$����J�Ҥ�/��9�*#��<�
�mOq�!��>#����T����yg �֯�BCYs�"	����נ�	�I���ؤ����L�"������U	KV|�6>�v��ng+<����M/�b�f��ʾ���YE���!;ͫ�$�Cչ�^1L+XB�r���L��R�	Y��ّ`\����h��f��)Z�l�_���TH)
�dOO-��sɟ�-Y�S0���"�z?�xt�q����Ŏ]����|��$�{��o]��9�+e$C��!�]&����|&��|f�p�5�T^����\�tx�k��wp�����J�San>C-M�ݢ滒�a��Z�DEx�ܙ� �+PYI�����\��;�����J~�!���]?�v�av�;T�vw5��Z3�D�W5��#6߶�\�����/}ݓ��¯(�^��mg�ʁ&���6���d.������7�\;.�������B.�_�&C�aq��A����J�#�Qו(z��n�+���,
b��E�P٘�o,:a7���
���κ.y��/"�v!x
swXxg�\���>6C,
I����\;f����x����I'��ڕ~,�тBzo|:W�:�{�(��E&�0�����3KN>|�0*�'T�*ՀZ��UP��k��b�ox�;����X�f�=���=�k������b\?�p)7�7n�A��������>,���f�H�z�������&�hޓ�~~+)*<sΗˋE���n�H��^%q���g�R��WnJ��"�Y�քGbtj�3ĝ��7;5�4�T
P@���a�\����g�&�A�������6s��[�+�V�zj����Fy����#�t���Ѕ)���	�p"!�ϪY+@otSKS0N���hŭ�8�ìJ��9�^��Ƅ�E%�X��E��.��i=�h�`���˚���|�Fb��6�$����C�����F��E<\�2h�T(	�>�#��e׵�Jm��yXt_�������s2^p�@�-�0���Y�*�/�huߟ��խ�H�����XE�q�N��$�*(����i�I+--��bCً�@3aq���,�'i�1���C�y�ş��5R]��z�+���k�����f�4I�Y
�6��]	8���\D�����m�G��\z�$�8vĤ�0�/�7\ʅ�Lc�p��I9�K�]>�{l�7���z�� ٸ=�BoT�`��-l`�2y`=ζ�W�
���Gj[3f���ok��5�3N��20HqF�r�7��O�y�f�J��\�����$�%T��ֻޯ��R�" E��=Y�w,��_)]��ڢ���S��i򸳖M*]�.abݓ�;��{�;f$p���\5p�ta��:��̴e��,-�i�إ��j�8�j���$�Z��g������4~��Xa,���FC�]�b�0R��O߿�G3��!Tnk�e4֫��ʨ��jiP���n<���;ޯ�z�[)�#���*���%�^���Dx��nqhO5L�yD��7��~j���Ҕ�z��l��y��̻��6��dS(1�s!�w��}W�[�S�Ԃ�%^�%,؃)'��Ӏ񾤍�}ү^�|/{?�0��m�5l��¦�E>Fn/S|�1>.��ŝm:�����;r�*)�$�Y��q�/�x`��n\[����`���n묈�w���J��@4����Ǿ���t'��|�7�� �y�Ї^�����T�}Kpo<�i�oG�����4!�=��'�.���5Q��t��k����b[U���v���9O׆}�,' ��B<�I�����TC�X"��!"(����]O+�(�Z1C���XbG��U�%��*3��~�n C���GtBY`]��<rN��1�:��qt|�����;�~�5x��e	+��da��ͤ�ѹ{I�gtxu/ˇ���y ܳ.8��3�*�mx�y���]2ٛ�k��&M���j�NW��yc��
^�"j΍��	�ӕ��ªY� ��i���x���n�s�@�h[01���������C\JU.pt%��AL��E����&x�(��� � ��¡�M�+L��,���r`��kq��$쥋��𠖶0�9dJ���/��� !��=�}x�x�^�.N���Ֆ��%�㡣~0	�����N�HpAg�PS,�Ka��z]͛U�8��/�z:�N����KYn�.�a��	�79
-�^n$(4���E~Z�P3#�����8A��gԻ��4��M��W�-���q1�����D��2�6B�@�P�%,Ě���g�����ya��i1����!"\��@�f�Fe@���%��Σ+���ȼ�j�Q�nx�8(Ǌ!.�,=��{V72 ��φ'��j�mS�a�ޔl��~����3� ܇�|9Ngu��WAُ���/�<���e�[1�Z��|�������ӆ��ZwJ�<W�?��V�d�^u,�A"^
8����_�#�jc"�k�뺄s�����^���t��7�Y�s��	�a�᷉��
�Rj�����k.�"��W�W��^r�q��"m<AwB�̈|�pc(FJm��6ll�����`Q5&\��{DE��_��`�+r�ff�4���������na�"렑f�C�ÿ@Y�D.>�/b.P20���F�=j�%e�p~�nnRҀ��g�Ml�y}�#"�Kv��}��s�	���s�A��j�V�-6d�D�m�4+<��55�_��iҸ�"�yj�p/�GtC�M�Xo/��o0��.0+ϏDH���U�JL��Ѽ���#l�,������}��3�1��t��j�mʨÒ������e%�!��г�FT�Yg��&�?�3�MZ:?�y�{��*�Ϭ���^įm��3�{W�p��%�zI@�M&$ot��W��8Ϭ�[� ��y7�߼\G�dr�`�^�����~��`��C��yH}������<v�j��!HR��}��0�t�<1�;��*\-F��Z'G�|z35���<c�=�8:��_*7�;A\!:�2�������{/���w��]x�M�ǁҝ��@��xH��wTX�� �`�[��C��wr!�YZS�:��Ƴ�J�wL�E�3����n��x�&}Zʉ5c����zK%� B�Uhq*s�z�8ꊫď-�^�x��2C[�m��[G�V��Bv�r�7��t�w�OS=��Gq%��"�i��*E}V������/ܐ��FA��3g3[��x��n�(���4J���K��o�{O���� �3|?:K�&1�;s&R ,���\!��ɠ�N-�A3�1��Q�N�%��¬'P�M���S��1S!W����`�Ý`l�y�4%��f���c9���O� �)�>%}= �la>.��h������^t\/ i����j�g���8�Q�Í_��$�"���sU��H֟�ex�6w�-W=���)���{ggeE��IP����G�
bni�p�Z����_�����5���6i��>�/�,��3~[���^J�':i�N��jz3Kh��ɾ�@����7�2�&��JXea}��)OG��o�&-p��Y����Y�M�5�ɾM�ki�j�����M�{X�nP͠'0��/�b�� K�T�v"�S�U6G��yCh�#Qh���M_L�0�`��;�
��>���c��@K�!%6Qd�����4	]mf���>Z����im�������;�[�Max�� v��p�n���2u�if�7�-Յ�u��u��<ٌ,wꜘ¼����z�ʷ���&�Av����B]T��Q�a��%SW���T���;�_R������`�:�7[t�	�gF�����WP�OC�IK�(6�)��>�~����a:ND�%������Ұ ^F,�$���%^���/�c�.D�<�V�c�j���UA�v��Q`���Y<q(���i��?�6Ӵ��tI}{I@�T����I6��@Z�������e\��Xb� �Z�m��hDk�ߠd���sU��*����.��@�"�0���\r������چ �3�%ǰ��O<�AF"܍")��&����Y�ć�}ֶW�#%qJ5B@dv
j�gB?.u�0�����׸� +�[:�;��m�����2��y7��kw8܊�NM�@8�6'��|�|�Z��}7�&����3�`~Eݟ�cC?�-�l+]�t:��n+8d��+R[@��ы�L0�9Y�t�O���S��z
�%Vo���dP颛���Ș��<!;�G��o�Ձ&�w�H8�89�n�MӚ�ۺ���P%K��Q�뎮���^� �do$�l�0d�,��ڛR����u�ʜ.�.�'�G[)g������R�8j)�Q�<���w�#�G)��*L��nh����GN�ޝ�w,,j���z>�]�7K�<�3a��򭟀�uQ"���@zD�z�e��<j�SrM\0�/��i������neC*v52�M�1������O���r��9�TTj!`Hz �.��	|�����@� �؍�r�U}M����6��H�Ƶ�T�v�ìE���et����A�_��4$'�F A���`�L���۬+��|�rw���}��oN��B��?v�vX�%$�i��,/mu�ў�]�2�@��9dↆ��֑�va�P�N���δ_�7�j��vX�eWi������2t��y$���E�����7��.�7��cm�鼅*�!�ϝk��C,k���ՎYGXȪ�_=;���A��t��}��f�Ӎ���Z���2������Hmw Hx��WT�9�	(s��59oX���S�j"�xOP�;�(HU��1w|^m%Q,6��2%�P�֣�fY�{W��S�5Ay��ާ^^����[# ��I�-"Ԣ辈�������`Kt����+q+�wug3x�J#��o���2�@�k;g:?���㟙��@��c�ȵL2�����٦���"�a��_�39�\�R3���á�$�^��y=5 f�[_���b�=@��mȥc�-���9���q��d_Q�Ï�B8���ƌ��]4��@gu&�Ƃ�|�|H�I�S���8p����l.'���]PF�gQ�WFq�1�>^;1;�� �/�@���ب�dJ4@�ӽ�	l�Ƙޖԫp&{���3u��wt�ַe5kJq50_��n�L!AkF���è�G�[�!?7.��u%�� ��7�p��3۷��U��ʂ�`1&@)����SQ�ߋ�8��$	y0G�%�?�A���]+O�&戞6K����Bm�ڶ	�&f�m�_⛹�b<.dw��k�z7�ځ��~�rn�?�����V:-VU���2xigT�{D{����䬗���Ɇf�� �M��}O^D�E��K$t_A��||�& �Z�d>t��+e㜠��"���]8�%`'����E��u�<@�É���ݮQXO\ֶu�C�%�ܢ�1��ϩ�5`"�a���/���y8�&�����ʼa�a�
T�:{�
p�Y��c�Ck�h(��T`A2�9�j�<�o�G�������K�?���;��w$0k��ȱU� �F�X�wLݹ2��dZ��m��C�&�޿� ��=\w�h���B"�v3ު#C�6�
ھ-ud�(�ڄE���0�����:����0o�v�
'��R]��p�QlZɊS����B�]I��1^�I�>J��?���D���P�5�V��m%5�r���޴T������^"�]J�,�|�;�80��T������0�lP��#�$���Ҽ�������GwD�JߴM="��D+0��&9Z��������fCDCJ>���?��"ʫ�5�t���<?I�~>ݠF��&����`W��L��Z���ֳ�Tb�c;�<��;>}�JFkj�ۦ�]�t��l�)6����򴺈��,��YstTbA��	)���.�9��!0�R��zq?�~��Z�{��Ff$��'+d��$�Y�!N���>-t&�(F�vn8�)aTz��ݾ2����>� �kT�r�r�/�C�Kӛ���V���%�ӕ�o��ܞ��k�>1�����]"�C��ѐ��.;
��Z��MD�O{�uj�Ba�����rw��)BH�a�d����'�pۆ��N��߯bF�V��J~H+��d�3a��w�|�����
��sٰf�A�r�B!�:����u��;|{�iSo��{
��y`��N0��|9zuf-�bz��>��^/�d@r�.l��;�<��v�6�\X�l��7Aӟw�]�꺺<�p�As7Oh��a��!F �/[B��n'��{�mg�b�/��z�u�뉖���N�Qt���H�i5�#1F��<������"��b^��o���a&d(�H������-JG���d4ѻ(I�H��5ƹ���6��Rx���h,�������׸k4�0��T�C Y��M��F.� `��z�^���6�_p��Z]�q��;2hζɞu+�G�^�Y����[ȸC�_���>���'l/�p��WQ���5�w��O�,kvwi<�J�$@�Ůpcٗ�A9cC�������1j����pMA��e���AZ�8�Vr���ҵ��fQ"�?� A��6����޿�`�u��E�d`>�2B4l�,�}�e�gu���\o��3�L�u��`9�E�+3����$`��;�>��� :���>���BbE&�!XN��!Q�����3Z7"+�X��H��
�r�����034�`�qۇ~bC��Qϟ/d��� $�<�iT�^>! ����z�⻟���e]-~�&�d�q�k���ۼ,d��� �;�I�`b"�K �.	{�{��	o�/�R;��O}w�i�J��q��*Ō�������s��J���/녾�ع��Fp���@.�I]�f�!q�*d��'�y��� ݹ�mIQ+�JI�c.B��;2�~'2gbl$8�0��AÍ(�6.�Հ�3��v��l/���H��؁eE+\O��y��k>�������	��6�P#�:�x�D����	F(���6�g?�0a�����{��b���*�<����o���Ԕ���I�6p.�M��>��A��Ņ�A��?|a�1_�j�MX���=1�8�ܮ�"�!]kjX{*��ʈ¡c����\��v*�l�Z������`ځd몰�@��v�H��h�׿`W�><$}2�b)@M-Ev���X���Nb��Ś��9�^&���;�;eM3���BCG�1e�qg���9N�m*�
տN_2'ZT�&#w�Xy��%�)h%�F!u��48GSW����K}w k��:O��P��.U���sP&��lR����(���?�J��ّS�\c�VK����V��U�,����t�H�)�����죲й�{AZXO����mZ�J��"�}�Փ8��zk-~�Q�N��	Ͼ�#�a!f�>��W���6��ɟ��T6@���f��Br��}�| -�%*�?�����@>wz^��N�EX���|�H7� B �V�A]||EI/��t-����D]i2���\!%7������/��� ��\*�����υ32LKH�Ǘ�\�Υ�u�x�����B^�dVKL�*�L0r��n$"#�"6ڥ=�C��6H�X�t�q ���A�R�Ϝ�M탞�>�i�����l��^�5��e���§��.�U�r�{�9U������)����7>��P��!r*��������>���c�=�,%��m�;?�6�g	���[ʻ�ˏt�y#=�) @6�2Z�Ϣ��ӽ���l��,T��.��Z��=�v�}�SF��j-���~��o���6�%�E�w�cHε���e��6M�P�]���*J��o������&�3p9���Q�D�6�%���7cP��-<Z��*��WvSp~��݌�y��~����?�o�\�օ���J�]:z�B����w˳l��{�O|�r!e�n�g:���_�߿U_
�1~�d�I����QH�8@C���DoiQi�XOC��5r���_��i;��(����N}���&fH*]׵>g�[)%�퉏9�L�\:)�wO���>�8�<��_u��b�.��(�<΋t�~�,7kW��݌��W��`�����Ɔ4Qibsɋ3����@���	濅#eTǫe}yQ�i�˾���o�Y�ܭ�89'^���i����ޯ�,�H��E���ih�F�|a;U�BiTG��ԵO��f�
����k6y�W��,�uc�8��SiC����R�2KJ���� ��ڨOoklg)����{�	��7����f�A�o��q��� RéTt��8-#���O�L@�R�>�^]|�|��7�C"F�XH�'�	�}T}�x&�3j�Cb��,ykDkiv��ň����$�_���]�7��m�腣J��4ȠE~��l���h�OXM��u���D�f�P���B2�O�����[Rp��[)�h���s�ƈ�zd��Bm�uX��0�hc�>���$��Օ�,zs�G���(Z4��t�9�bOR���#�B��ES��)�39�70 �(��Q�)���Θ���x�	���]�l}Bm���~��4 �w#���L�|�����I�I�]����b�'(;��������j��Uu|b�K�wGZ/�]��� #�B�/���&XO& �"�y5 ���a�w�\�&��6�o<������)�]���/�Fc�v&�ta<B?��8��y+ce����se��O}x'Ja{���L�_���+3r]�,3B89�T��n&��Co�̈�&ݯm8��3�:�D܊�����g���D}{%3�T���{ŏ[�K,��\��y������Ӟp��ÚЅ�&J���,'w#�A��pI�4�L;`�n����Z@��O��d��!GU�n�M*P��������y���tj�xz��v\z�1�|v^�lN�Ob@}�bd��:d�I�Z�/a0>�}��O����,�,DPF�[�1��?5]l�ք�*��zM�B�L��2��Ӧ�O�fD�h���f?AM�Bs�QŋbiS�q��\K������bh�i�����?�HP�[F����}�qY����S�Q!�!���a}?i�n2Lޱ��O����U�l�K��O|�c��A1���?A)*�@ 7R�T�CM�u.�M�5��#dN�8*����ZD:��p�~!Q"���i�>����>$a~��'۹�F�_�N.oI��j	��v~5|�ǨnFrM�ޗ��h�.D�sw�Y�*X��n�ۙ)a,���V듮���m_�%��H�ͬ4$Fkk����#:|�VB�(�����^���W��͔]1O�Fҍql1�m�,��t7�aT�*��6��A7�RSF4*d�cA9��I�:*k����ҥY_��|ɖA�MB>Ńy���e9�B�M����G���Y�B1j��T��Y�z��^�d)P@I�ą=����r�9��◀l0�#��y
����gSD�i]@ht��{<��ߕ�e��6=s��eѐ8�`�$|Ƽ�s�
��#���q����*�&�L�9�ж��9����S����`����VY�M�%P�v2)}N��a�rծՍK6vߣ��c�f�����՞�PēO�]��W@� ƶ�=w^.b��E�0�N+gD��I�n���h��\�M�:V���8[,X�V���[�&��r�Qn\�?�N�ƿY=A3����ǖ�I6�_᫙�U��[
�N�@K��3Z/a\ފ4d�A.c[�:��+��n�V����O�v~�un���ubKÕPٚ�k�c'1�V�e�Nj�b�-i.�h��um�u�Hs�@��?W����\�
����Dn����Рp��vG�W��M���֮���8�-�pK��I	N�w˖P;bȱ�� ��#��Ƞ���Qɏ\L~8�W9��/#7�D=�e��RƏ�MA6*[:����g�生�<��z\ՈBg�.�(U_Ȭ�<��V$s�����>��H�p��@��ӹ�K�/�q]���6�le� d��v�L�z��(�U3�ҿ@���Iޗ���߹�>+(@�	�RI���0�%��>ٜ��K!>���|�/�*���Y�ػ2��ӯi#����e���f���R��r��u�����I_��ߑ�o���|�2G�� ﶔ.�F��-K�yG�<BҏcgY�^�.��F�\�ߝ�CL�^1�W�Vf���4	0z?9F���<�DX���j_��A!ȄYAELY�c�ҠE��^�A����܂��4BZ�&.��h,�P`�Ƴm0@
rG=8��Ú�����#����pl����IF����̜۶����q]W�	�]�������[P���?���U1FH���bB�$]Jk"��L<~��a�5/-ko�xM��0�'&�T�i=���s�Y�t0f�����S�ƕc �I�m\���!
l�2~Xb�03��Cb�O9^�:o���ܛ��QB���*0�'�C�Fg�m�:td��J2�v�KIu����й2 8��@�S�6�+F|���I*Aj���������H�ϐdDn���4�s��}��k� �j��Q�="�R�H����n�����bJ6ק��Jp�Z�Ok4IfN���9]�Š�T��:l�4���6�ϿX�7��Q,� =w�������.b�]�# ��Y�	hI���э�r��hȏ�\���j��qf˦zC���`�nm�?��eueaxD�P)�p9#V�{ll"[�P%��-͖���`��/�%K��:���X~?�*^�MV��	'�8R�#��_�?���@�>��x�^ϴ!q5B9L�P���u3�`/��F8ԝ6�*���N�'4irX8:�C�=�@���+ r&�7�_h|aB�_�@�xLߌL`�h3,�m�I{5�.#R��'@��-�X&[+��]q#i�A_���B!�y%�s��1����]u�*'�T�Q����S��w]�����}�J��M%Z�����S�mA?�QE�y �܂�5�����B'��F�U��?͏3 ��E�3(#=2�c�v���#y [oe�1Mnx��Ǝ����kN;���֌k����������Q�X@�X�\�ڔԪŜ�;|}68F��o�Wo.X�|�W����"4V1�$k�'1�i���B��d>�̂e@4�s\+BEǴ��P!gm:Wi-���c8�'k���$>O��`:A�ɕI���M�g�����)�,����α6�uCu6T�/O�����38��=�uE�]���ތ#��#Pn3��?���wS
�N�&?�'��+�h�p�լm��"NX��r�͕�6U���n3��RDR�Y%���Rr�MA�l�t�h����W��C7\�Y�3����I%�P�Y��
eʬ�M(���S3�bw%y�Vs�kYV������ϓ�v
�/��]si�B��HI�y<GҌ{�t��vPU�z��O�h` /~��t���F�Z�#A=�����w�yϧh�$�gYJ�P�M�����!U���L����_�r	p=8�?�x �:A���W�{-��G"z�~��S�)��{��G�����7\f�N<
���J�7G�v�&>EL���T-,dP�MD�V޷)\�g�L���#.+T�G۳kr-�z�"��/�/�N"���`���	� ���I�u������r���"�D׸S
u�%�L����`nk�M�(t���	L-Y�������F35u�	X'.�//�gzm�%�Kڒ��+��&�T/�����^������X_K�Q��X}�+S��Q�&�kW<��q��G��c�q5���1: �ز��;tAi��s�Ɛ��AF�F{Ǧ�A�C�|�������#�q��t\��u�b�u\� �E�CoQv����>�zgL[������d2�W/�Z�%������`s��fcUu�M}K��;�|Y�8�˥���~ˋ�I�db篩���j���N�K�����]a�O����s$�!�7�*N_��Xߵ�D�h�����U��ո�t�Fn-�3��Rmh;�ޅ��5�C˽�U��>��VC�j��r!?��'��V��Ϡ_ҋ�P��6g��"l6D!��8���CTq�$���-��P6V�[�������r�A�2�m@�{�r�$��v�Yw�'�b�؍��\`��p[�-�i(#Qo�6;���̝U�G�6v8~��M���`�����tq���Z~�^�h�糤�{� ���%(�	�3��/�|��[e���_�Y�FP��=�ٖ
еp����?�Lކ�87�+=?N�/��Ó*o�\�{~���)[߱+sGI{i�e����͝��*����X(�6�p2��	曟n���(0�y�U�*I�xt�����6�\?LD3_y���U#/�4���\.ۇF�*��5OMB0���7劷1��O����مI=��ցa�qA����=(�ycE�bO��=����
z���x��o�<��F{\@�{~�1Ǿz�
���z��{6����&,$E	e������d��x���Sp���2�#r�/��)/\ǝz�)T�CR���`�Q<��ȅ*JJ�Xag��`0�k$1Ё g�gl�
8}�@-��'ze�v�1ҊP�x�a<�%/b5a��ĬG���&{Fxu�7�'�vY��O�*�0��vx��`�r���
z�/�w �����V��9�gO�i�������!�����-Sˌ��gT�6G'�Ƕ�1 �O�&�f� ��~��EkHS~|���m����򺲚��;ڽ?���UE�H�vz�t�.��s�ʱ��y�����l��li��Dƚ˵�����X8z�r�!C���_��^b0�}��^3�*�	�ճB�%i�"_���Eq��;cZ��e������t9mlb�[>����Ӛ��8���W��NJw$��Gʽ���'~�e%��P�D��=�aF,������8O�y�!�Ƚi��*��IX=έÁ�,S��#�����8L^t`K)!7���ܥ$���������բ���ׅ�����]��P�Le��z���&�d0 ���K�����{�����Y�Ψ�d/X������Ye�8�i�� �{=����L�ԧJ��v7#ԨRz��ĥ����5`H�G���K޻�w�ClE
2vq���q�v�i�i��w]���J���*>��塢Ytk��1M0>��-4���K�⪠�;����>�,����>���q��-���W�umF�]Y����Td��x"�z�I2Z���&A�G|�Zy��_j�a]_��y*S�&?]![ \�D���H^��i�a�L�_���R�Г.\�I���lE�;)�;z��$u�LA#�P��u,0��V�z�O��:1��J/�|[�A�6Lռ'��6�_Ș'��: �?�̗���������Y�ޞ!�2JɲH�u�D�+��w�
������߿�Z�v^�Ը���`zyy�E��?��]
�'�>	����*��%���I�?�"�6SF�e��~I�sT,�V�N/E�\��;?ġ,��pռ�lms�kZb1L��_�y�o�*^Ki��@X��.bN�p�Udŀ���vW0k��e�*h����8��?�)`n��3/������?�l�NbqH� E���F>2�-�#러���0\��޻�n,ag�*;�������2�ׄ�Ї�l���f
�����/�}J���1V��4-����Ơ�M/H�&S�d�����z�z�k�Z�w�G2�M�(�Jrph1��>T/Q�Ŏ�@�K�֢aa|�ҹ��)��D��~q>��?Q�	�[7X:�Ec���g�N#�ęoNkdl!"���1}��6�W]I�?!���K�7qo��O�u�2�(����`�ڱ%4��	
�%u���e�4���_nߵ�xnG�0��c���_OnO܄*y��xy�FE �K�x���%�Ԥ�:A�C��"#I�)yWr���F��i��ۂ��x�E5yc퐠�{\u�o�V/Uy����h`�6E��mD9d&���69~��#�Gu�E���V���6�%m��X]K���;'V���v�����y����ȥ�|�m0��!��Ȥ��)V�E�aK��}�
���5;	Z���r�?�[�l�٢$ĺ�G�!*OV�dn�$(��$`"��E�g�D.��� ��X�=�Z<�fm ?-�xe( }�i�2?��HJ*�B� �wT��q$��>O��Ըc�e��܎��X6X�˖���D;��������k��$�_$
4����[�`�>��F�~�pl���|J W��&�T�_o1�̝l߃��/�5Gy_Bo�g��c��WLw ���8eB�R��P'h�(M�.�)��k
��63��^�EYI��l��_#�lA>��M�2w�u��:�:��'q�_����s��xK_̝ѩܻ#2Ԋ�yWy �t�ZY�!;JV�e�T<�T����#$^�dW:Fӹ=г0QtL�Esthɍ�����2�V~�8H(�6�r�!��c���WE;�
�]J��$��:V��*�l�U�|8/ն6ƟI���u�G��Y�>���c��Ova�T;����[�d��ٖ�<K����/��RB�\�~���+�9�.�ǔ������tz�Q�<��:ߒ��[�?�����o��AVa��FQ�/��0���qS�[GD�Ww��^ ��O8p�&��1��NX]���꒓ ���)8z4��p�J�����?G`3�!��HE�jZ�C�(�;�%�S��(���I��ӆ��w2sq��poR��T�(��3�vjsݎA|�uQeGeFt�'j�!�%��@����r\���5J/�d}J�u&@�V(��U$����1�% �
"Ҍ�Mo�O��*���#Y~�����|�߸xj}�J���M��P��xS|����6��C+a7$�#]x�N�nO~�ٙb'u
U��i�|uQ9i&�߂;���yˆΑ���}�"���S�d*<��1�w��F3{�,1���60��C��\#����?�j��:k����.��l�Ǿ��r�°��$�h���_��d��x��_k�H�G�����ث;u[��G�+�^E{@��Sl)�v����9}�O�d�6y]8��ˊ�M���G5�H,��c����ʁ˄�g��RW��l e�jļ�'h2�]5$U�����P�4Q�����>������yP
��	�ݱ�d�<X�*���k��_~9|��ɞ�5�+On;���?&9�7���ͻ',h���Fʩ1��,���lגuaK=ajA�T9�ˮ��?������5W�;r1��J���
C{����e�"b1��&�D�~�n��%�t�@�����K�k1L�dGnD����N���!>_*_~�
�޻1��1��"Ŕ�qe��£5����,Q��K��o�yh����[����s��^���"OF&�=�%���_�%.~r�h �WH�?p1G�����<�m������ٔ�s���z6���8)�J��n����vŧPI�,pV��g��X�2���>��Ɋ&T?\l�b��*���=����bc�"M��m��X̛d�J~�B��t3h	pV~�T�����,Vn�N?�x{B^�I��5�G΁�)�d�p�D>5���_��0��
��Z@q�S8t�T����6��:�?��JlޔDł�={��̠�T����B��Z�����-�2�C��v��ֱ*3R��x�����pQ|6J����7�� XSk�]��x������ �Н�0��Й&�׸���]dfb �X� �3����d��k+	J��ɿ'���u��:1fP����/L����H���I�k�S³���kWCS�h�|_-���ބ�LzI2�Ne&s%䇬i��3��M�dqhQ5Xu<�xk�ߛ�dz0��i�_�B6-?���Gh�g�$�t��a�ڄs�t��$��C$��-�{�%����Tx���Q�l�(�!W�EU�㩒�J�JԼ���T:�߫���x%��f��N%Gb.
�`k��(Kr�r-���P �]��D↫N�8����0���J�!lǢz�<6�<<O��������+l?���Ǉx��>	���8�Mܪ�	,�e�Զ��Q73gNO���� ?�V]|�sާ� ' �.FO�x����[5h�=>L�O�]��/�����ի�']��u#��])�C<������-[=�!�[��� ^n��p`
&H����(ҟ'��Mω��M��V��tX�hn44�; �n-kK�Z1�nwǄ@��b���64�C�3��ot�8
v���T �×���%��{�^��G^���rZ�Y��PJL`��neb��F�1к[�ο^an7����L�]���Y��镼����{�Gb�6Q�W���6�'D�T�1{xY�~��r����&�K��4�T�F�T�Yn�!��y�;�Cj�7�;��a��D($6�!�.uK9 "=��S�ç�<Š�2�3�́U%��� U��[L�tLO1�ţ��ۺ�^����%�����+�8l$a�:��Y/���l��m��H?+l�ZΌ�$�n3y6k	p3B�IZ�h۵>�+�0��@\9�@m��zk�fʞ�!�M0�ZA10B��H�X�$@�U�hc�>���\�0o��D"���(��װ�O����?� ��@��J��?�i�m|��.�%�x���e@�:J�ٰ.|�T���k��~Ah��ߛ���TܩtW/����1%�v8�WK��6�b/���D�B5��2B�ϙ-���ƌɘW�zښ��L�����o�Y�d}_U�>�N��>F�J�ǩl{s8'�U(YTv����٬B4cB��(�%�=��<��c���g�� �q�yv8���l]?"�p����齦T�Gq����{]_����������t�FXBQ0�.S�AB�:ozL�	}�E�l��`$�cW��U�űy�0c�j�p�}���/g����=7�	��f�\��΄�]��Kw�/�s�(2�#�]0+�d�A�4s�ܢH�dƩ�D�%�O>e�����pgg�-o�Y�)�D(�f���]m�zBG<y�
�xvm�jd�oZ신�<2��;-�{C�dǧ ��@p��SS��D�d`)ϰ՝� j�q��=,���rD3'�AV�89��;����X�8X4����Z�ֿ��WD�)�_��Ԫ��z�Os�@�7ڏ�����x��6��6!ϰ�hE�5��M5��gk"�MV}1�M�9c���M���s���J�	���I�@�6y���!���Z��BI+#\\D�,���<Tf�_���ܰ��U{��A�P~�z&Ah(�P�<�jF�c]�w浻�.4�M�`�}c�=�ʁ�#:eY�~�Oy����F�+��Ɉ^���}�X�8��
M���?��X�������pR����c�uW�aFN4�1����嗦��|�=�'����-|�S�;$�E��(sI/��O��;o�����X�Ix�@��BcF���C�%�1�AseiP�A�~Pђ�2Bɠٴ�����s�x��E0��ӥT
��}�_��L�+�}��4�Xi łF����1_��*S��OrsEݖ�$`K���I~,A�������ᆮZ�E,$��@G=`�pD��4X"�i�����bb���-�ζ��5�~k e�I&��[�z�J�m�����Շ�%ɆE�Mu�u�6��O�2�R[�G���⪟�t�8֫DN�lJЧ&���	�J2Q�ko�Z�({���pG�aH@����i�T�<����M�py�##�:r|r,E$�]%V���)+�s��iCb�"���=vs�%�0�U@�-d�(@X�� 9�Ѯކz]��o��Fq�r0ߣ	��1��7oa>/6@�jcϔF��,; rdp`�U	�)������n���J�x�d�$�Vht{̨��}�j<t���� ���E1ctDE�n�,D$�B+'�	V��%�+�;G�uG������2)CO���L�A��$}�T{t�)?�����hE��v�?����! g�9f�K/�ݬ��??�#g f����?�5�����l����o��¶Er�*�X	�퀂~k��`b@�?�<�c��q�,\�5h`�B 1^_�����oԱ	 ���z�gQtŶ�Q�&�ڮu�nޏ���#�'�;�7]*�X���0�U�=\Na�����P��J��Rn]{�������SN��ҲTZ���;c�D*���6b1{d����u�'M�5|x,���*�3��P����Z`������&�]H�U�S�*�#$�'ji[�Δ�0^.��d�����������%��W=s/6�/��_�|��>B͡#�[#�/���/�qncK%?��x��q���m�M��mGT�ag�X5yyZ�"4�w��nU]���Hn�ǐ��w����4S��T�UL�;�N���e6�@lQ��#i?�o��{%�<G��/���j]
i����PC7����fr�,��<K�d4g�dc���pZ[J�1Xk�z���m��=[ȳ>�y����Fa��:���q*�$��}�b��5�d*�ކGc����*;u��d�`b�#�1���P#���uУ�A<�SN���~��_��z�d�����ӂ�r�Fjп�s��F�c��|�P-yw�:�ߋpG��)�E����?��ң����:E�w��U��F�Y��Y�NÙ�)[�s+�7p
Lr�r��e~U�W�n��q�c�r�˙W��K
�I�Z�dM=�I��sŊF �6<Y�j���\�:F*��(��HVt�ǘ��Q�舺�*x:��p�b�Xq�ѳ��,�XY?����]_{"u�z���c����=� ~"����Èa
š^+��&ن�'n0/1*�
���D��۳��_J��>�� ���=�m�;�8/T\P�wӚ��J���UlG��T��fb8N�Bh��oGb�T_����c ��a}�]�������K'��%�}Qɴ��H߄�/$x��Gve�����PTM"N
͠�g4������q0�L0�i��R�C7�r��Ö��Up+�i�B�YNϔ[ňs�u�u��$r���x�d%ў��r���9t����{�V���l�On�I��O�}��s+��}�^Þ;?1�Q^I3/Qs��{� w�,��M^��!h(�.��k��g�Ͻ�	� 5��Tq|�%���w/FŬ�ũ+��j�ms������+M�/��-�65˚���I"˲��S��}�8���>���#~���io�A�Y�,�э[t<��E��5�K)�9)�%�n:�	�Q;��t�F'y��&f�]S���F{�3qD2x�[�
ڒzA�e2��-aL-�w��.�-	��F-ZZD�!���f^���X��Yk��r�V���DY�%
�{��\Z� �6�qdx-��N`O�� Z�W�	8T�^Nv���r�S�W��!�i��*�{��m*a[�7�[ ?����j\�J���!@�N�(C8N���6�Q؆�����.��[pk��(��9���!��:�ʡw��?��P �.�n�u̄2敏b+����fK�`'��� ���L�cO�B���������Z{Y�{�d5)���t��B,� �q҉�b�i�������dZI�L ���`f�[�a�� �T�J�q�}���������Y"F����E�YP~�ӟ<����9W]�/�ƭ@eC�B8l��O��y�f��N�����2��6�x�\.ŷ��z�H\�^U]���cf�޶�#�����k��M�շ
���"�8������r�
��K�]�;��g'�a|�*�oL �MK���Ș�5�:w)F%z�hW���E��_6ȯ��o{ǜ�t�^��J���\F��fBqkm�6�ץ�š(ڗ�_��A_D�#�H��S���pZO�ٴ���j���.�����#~Z�䭜����C��FD�m� ��t;i���5����I���	c7!�4E��箘���FN��ohg�|\H�WA.���N�ZA����W���m����fj�<�/���s���f� ��i��U��-�Q�ᅯ�]	q�_st�����ɐ#pȻm��[��.dQ@�v��\E�@�5(�v^V!�
 wO>;W�0ma��Z��M���r�Zx���R�X�*`zX2j�[,���"�����^����"*&��7��P̈��|D�|�v�kw��>f�ܮ6���^�>��ѻ{���|V:tIg)�'�>���6]�Ծ���#����󭒁;Z!7�}.�mxV��6y��3��9��\���9����!{O��␬��v�7��3:�G�% O�G�X���KI��<EġC�2w�e�����A8|�vG��G��������!�9��p\P#���&hVum���U<n��0�$h�Ⱥ(�}�M4�1T9�`�D�峾$��~y��x`~�ܡ�(�-$��P�0!�����{��T�贻1�>�4E���1���1g�1��(��^.G���U�{PV�����h*�.I�S_ ���|��H�w�¿�*��������v�u�ur�9~�Ń:8�	w1��*8��B� ���j6b��P�^f�2�$�pZ�m'�J�3zH���r]A�5�}n�x����h
a�M��6�	��	��a��!ы��׮Jb(���ﻗԀp[��(��7>�5ݤ�O:O"��۹Y�݋����GU�)�����z	���s�7�*.�$%� �$��&�-F�N�N��..r��+v�*�ox���&����nH�Q��HU�_��b�/�w����P���?�n�ʕ�1M'��5%��&��@j�Qo�tH���d46�6�!q~ ���8��G?���d�3	�W�x���g� �Ӿ�� ��Z�3� ��+�N���\�e֦49�o�$X��l| �5��1'r��}&7?�`w Ps��/IkU�~�5ms��)�3F�H@�����i�1叱K�y $8
����aʪ9��g�q��s̆�����\mw3���|�_6ˆ
��<�1��Te��%J����=�&H���tt�h�"}��+ل�Z
IS؃����CXqpN#C���O�����צ�{�[�ΫDi���c��!��x��'�@w_�j�S\�%΀R] �xӴ9䇒�{S��;� /��� /�Ӂ�<֗Ǝ&�x3󵿛n͒%R�d�f�����ʰd����5R���
A��,Q�F_<�dE���A,�B�z���+RYP@��f��m6���
=��U�!y0���x�aeؒ�=�� ��( �!<��τ���|��zVł��o�Lsk`2���϶q�~�������2�09�m�p���x��<�'����ˡ�ԶOCo0�Z$aG��i��R�>QbC���0�أ�C��5HY�3��{'+�4�e�-!�uշo���ٶ ��p���H��S��0z���ު�{�{ǣp*��c8S��4��64����A��kN��-���&������B=��TW������E�Ї���E���
�8�GC�]��J���-M�w����n�:��_
�`E()/Hf��v�. �S���!��:��t�U�ܝ,WW�tSHM���@�����\.I����	O��j�Nއ�ˉ����y�Y<�ol����-�&�f*3�
���-i�~�iV�ๅ��(��t�z�5�]N��S6���\u�j���*  ���lw]a���a�0k��-Vj��I�P&����͚R��nc�e��r�\dwqe 
�g��E�E�_9'[a<"���^Dt&DT��W�쏳*�Ɓ�d�B�z�B��W��Bu�97�i�����6ԉ+�HЁ�8B>�&�{��ݹB봱���M�[���Ѫ<�>m�$��&��3a�����ٛmk,6]�?1���5�k��~�n� �b0x��vcAR��]'���)��72�]�ma7څ��0�:v�"ū?�E����3]�潱��p�ƱL�у�����THL+b�M��L.� �D�a�dQL%k�=s3 ��T���&�����g]�O�ƭ���Z_g&2&���� d�d�o�]�r��]ki�b��*"W��i���KcE�Vl�+�=ΨYq�|�vߍ�40d@�_
��_6I'"ey�7/ꊛ�1'İ5���be���&8��^�p�X��g%��U�4"�X�����P�q��2�|��B��&��[fQ"��Dq��O���e:V�^:8�K$w�8ڰν�+I�Zj�*IREoWf.K�A�ɢ3�2�^����6���]~��(�N�zE�{����'m���4n.�MH�w�1ֻS'iV`�6
�6��H��c ѧ�^��0:����V��.&�0���E��'^;�6�!S��� 
o[!�7W)wG��\(gU��Ρ�*&�&i��@\���k)�|��Q@���c,�P��.ŏ*[�п�Y�uw(,ʨ˚�CL�)2����4�S��
�b��|�޼gS=��Q���Xn���:1앣����p��L�Uy�=(�� ��i�܍�PO`@���x��!�F�
���3�ۅ��l�$�`�^B�I캒W��?�$pU�j�]��s9��L �3��V�F��t��Z���_��607�ȧf��
�$��0i�=3P�O�X��B�:?۽��L�m|�%Ŕx�1��P�@$�:�9��1\!�J��QG���V�
���.ه�5�����4���C>�va�)�Ȋ���{b��M�h�ۜ�7������F58W4����e#v@�"�Yxy��|�Ҏ^�{>���G˪�s0,�J�I���[m�l"Z�·���0���2�1~+i�t�{RW�r�O�3B��5�K��_�C�W4�/v�Ð���|���48���i�u&��cm"}x����X��8�.���0��4Μ�Z���
�D5���/���I��ɿ��XV��K���d�u��.X[����qki���]/�Eu�?�w|�(^����u%1y ��U5����|>n7Y�xϝ��Ғ���VP_]携fM����č��R}a�H�U/�e���߆c[�΅�n� � 1�GG#nu�����=��,of�:�PeJW���~�� =�	� O�gc����Z�����}jC�·�7{��q:�������_�{�:.m��2\�𒔓7A���p�{sН~�xG�P�η�\�������e���|�#��TB�Xhe�\��Eܲ5�=b�?�G20]���G{f�kP��B+8
-��1��PL�p��_C��ԩ}GJ{��!��2X���:-��(hl�5G��~"��	�;�8���]�w�;
�x��g�=޲U��R��U�`�m%v��)	�A\�I�;�Z*
��CL�M���U�<��ay��Q����F	���_t�܋�e��/���R"ڎi�l�s�ӧ���H�4~��.���U�Kӂ咴���W��H�dJݪ�fū��X�����33����H�ϪM/�fup���Ǚ;�/?8��z��ZP�b4/2��d�x*�_+aJ29����-U��y7%l�m�2F�ݛ8�<���N�sԃ�ke��1�K��}T��G��yIr}i�B�--i�&�5e{�X���'ױv"�~�h�P Y&� =�46���G�C��7���0���+*P�=��+<�"�"��.�+�*@�z�?�KD �}��n~1�%�"��
;��|��}:aT~�s���0DŃdH�����{���n3��C�Q���1v����}�V��e��P�/R� J����h-ف��	EH}C���[��md��+���QD��wX�8�I�5��]���ee3���K�p��Y�4��k����S���	E�7��N�C��\Do��N6:�zS�J`(��u�zun��&�5�
HB��%�h�
�LO#�I4�Ծ�!���&�KN,pm�����.��������X��%Ɋ�ox��L�f�;T}��k�͹Aʳ�LoޝH�7jJ��oP�u�o���I���4��BZ����������]�KU������b�%d`��!�Ь�\'(Q0%�6G�Pˁ'b�PW���I9p�jC�l	�s�9�Cm�s����Ҟ�~'�Z�7R��<k�4�+��=��~��8tqU�� &ɢ�?���wZ%I����e��t"�c��k��J�0��Ǐ.����܃��fXk�Z��fd�S��-���>�$k��l�T`d�f�8~-��G`#�]�<������8%�a�`�˷1�!i%W�X��Aɷ�#?�<$��m^3�V�k�t���;\�Z9��gf��c߮�v\�.�-Ѩ�@@�b0{��1*�9q ���f��<ӧ���Y�����5=��vª�G�/��ߜ�#*h-�+هI�� �vKJ�'� $ŕ�	�Y���j��bq�B�Q"X��]3M���B6���o���a��ӸuR.p������_�O�a��G��J^G�M���)=�ڳ��s����nVN��۹s��S�R9P��|�Uɺ���$��dxI�'i��̲�R�G�?L�NS���s���_P�)�z�mM�b�\���}2�qє�T��銩b:.$�&v�}����'����LA}�](
��_����<^@��m�S��@	�T��Ƴ=�P�����8��%�ŧ�)�3��b�ɬE���e~�m�y�g�deT:����m�����`J�qg����?+J(Cf�� ��{��'a�,E�DH�԰���!B��er�2Tv�L�k����t-�rw����fgDyE�� .��w�O)�IP%�cnFS�\�1���)����Z�O�wD�z�.sSB�Cމ���<ɸ��֒ۯW}��z�ѝ���\�rGW� 9o]����|7�����{JW���Q�U�z��]\����j7����4�:��t-��z:y��r��&���O~Y�^U�y�}�3#1�!q/#��I��̭7{iǒA~���ֺ�t"dz��QHdw�S�4�P���B�J[�f���5 {C�L��wo9F��+�|,LR�j����2V��%���ft�t�̙Ϣ�|�v~�'�D������M��0�DH2�n�*��ߡ�Y��9����c��h�B�G�Sm1� ����1�����5-��	�2pG��w�߈�vV>)n3�0h����1����aJ+��X�S�L��Y^!�R�Q��i
lE� �S̽�)VY����"��~tdU�UMc�����$kL?�j���h�pwq���8�����^ST�a���*W�N���}�� �W�j~h�LL�iת��n~
��5���;�Q�/6����rc���'HB&���f.�}T1/JQ~1��ղ��eB	��`.h[KN���8�IF�F̓��d��Eֳo1�4���%�������0=%6����>���Q	���!�p�t}L�������[M{x�H�ȁ&�G/�:���p�W�h����p�z���#z�����)dz���^��-���ƨ�8Y5}��Up�j\qzgzc�`��_���Y
�x�g���{c���H�a�	F�Z�3{ڦ��-o�bFCP�U��ܐ�.�-���/EdۅԪ� ����,VE���S�曶�L/DZ_E^�Sg!�"���T�Bη\El�!��gt��)ksK�{G��ۤ29.�O���	�:�9�����м('� �/eӷ��� �� F����Yn�<�B ��|����Wi�f���vM���xO�B�����ˁ����qrN�c�eG{��Q{��'����Y�E�ۋ�׷�P=�.H`l9������2��y�9����+U7�!�Wl��i��K���<�����'����)�IE��P�fL�M���K�~h
��j��K1M<�) ���xf�:u'l��C(�P�^CO�@���&b�܇�#:�a�l������Ĝa�����dI�X�v���Y
��Ki\�̓��� �*9�R�n0sK����L�-O��Ұ�����4����M�d�H�=0|#����|�W(���y�ug.%��F/�g�4ZW�?	�q����<[���'fo������f?xƕ>��J��zwv�˷�5��+�ϐ��+>��m��`��؄�9m��O ߴ���u����[�SDɨ�\�!��A��+o���o|25�]���|�r"��hD&D�����ʆ�H�XS�HO�c���T�Y<�s�J,��̹�MjZ/�����B��Px���3�.ر���AZ.Vܧ���Q;���lWs�Xp�z��P飱Z:s�~auLum:�}^8hC6'�Ɵ{�,G��Lj�V���(���������"8+z�LxW�
~�
(�!^��`N�)���mp��$�Y�[�t\�3w�MG��2Ng��BF���C'	"���GȤ����#�kp�7:p��jx[X4C�F��7� 1zU�-2qʗ(:�9gW��J�p;kg��	���m��(%��̠���
WI3zҞ_ű�HC�gߏ,�V̭.B��H�(e�,��B��;z]	��C���G�NY���KP�eRm3:���ַA=���.	�!Fy��b������29(�=�6^����R�}��V!-���U�
�:���9q{��-�E9W^t3���q!/����䕎OkC�y��pF���+I��+	���I]޵������IZ
�p4Y��Vm*�:U����'������S�$�E�$� �v-���.��1��P���2ʰ�7������a�5'�XMO���ZG��|*q�쐿�� �3�sK���r���m��p�<#�*��1oFB�ŷu�l� �2���iK�Q#��N�
1�ԿMy�ԅ-��f���}����'! ����y$i�2�����B��=^�g�1��A�=$0��؍;{�!����\-{#���2�lQ�L���x�4�	��w��L�G@CWڎ��-{�s�+6%`���Q�ؗ>~�y�|�{B����/�����6�_\�ƕ9���9����wx+����A#Q�F��	H �MX22��P{Խgh`"����o݃�)߿�%ku��RۡԬǃ�V�q#�aQ����ܥ�Y�:�p\��@��Ψ�w��=��ϡŢ/�_-d������=����z�6���6��%Ub?.�4���P�T����<���K[�v��I_Ң��z�gȖl��Xt�ԙ�.���
�Z�}�Y��/5�c��Y�~���"V�]��� ��8C{�P������'~4Pk5Lj�tf��U��ZQ�oP����2�ƕ*q_-����z�l�ɷq� 9�G�˧
\�|�;�w���>x�l\��YCR���������yO[�]�~k!��;O��Ĝ�?�d�5��pI�y$Z5b~h�`��ZCw�څ�3Gh*�rQ�G���q=��TĥkMs�9#�L�k� ����ܔ$_��g��ս�C�jc��̸K���,�J�IS��0p"I�����@~�`�zj�f�C�m��+�L�N�`E'\*t�0��g.U:�����ZI��J�����R�%*�3�7M�a�b�s)�M��%�՝{��b���<9TM6�N~���:�cr���3�������_l� 	W�%Jn�tR�[�(ٍ8Ao��-�vR�	y�x>rQ�jh_AAS��Z|n��=�s���
�@�e����[j���}�T�8��2T�^z�XP��
�iܬ�����G���޴d*h���8a�ϩ�m�!;!� ��:&���Ht9�����d�2�9��� _�_ׄ+f�L�ɐ�?�H�d�Y5�m�6�n�^�}-�h��i;��|/,���2O�@���\%�9;���@J�f����:Z?�.e�1��'a=G���	NB���)
�>0�@���K&-��,l��q��
�>�/d�*��J2��� 3I�* O����k�a�)bNaf/��q���D	2�"�Ļ�NPڕ��O��2�Tﭛ�ݞ����� )@c� �y�K
Mg��+U1�;��s�[��*L�M㧆�p�D����f��.�EKu�F	ä�뤎�1Ru�%�"�O�&1�m47� �.�S�+ GD`{U�E짵lv�]?+h�EzȌ��"����w�%���ۏTꈶ�)�k���0��+�~��\z�W=�%�.n��K&�\����KK���Oĸj,c/��?��JmJ �6f�ԥN'��\�(B�4n|�_G|pɋ҅k���w"I�5#�b���ex����"�E��)�+���űGWoL��7�Xa-L���1B���7�me{K���yCV�����V*'(� ��c�ܒ$�b�Jv��~6�����u���Y�,�cҹV���4��p�g���?/�|��g�7s&���I��Z�r��u�(� ���.�
��9�:�<��<�a��3��=Xt�q�Jyi0u%��;w�a0r�-���rM���F�q@�D��	82d=�w�i���QU*����%�eDu2�ߎ��e��}]@��H~�9��ʹҌ[�B�م�����FQr�f[���7G""���b�ˡz��F�Coh(q^&�xZ�n������,MH���уۇ$�h�m����'z<�A�#:���!�lء���S#7�Y�|a��0�{b5�K��8�A����D��oqi���2�}O�p�A*<Lk!��\�%�8��!��x�b��!,-_Őib�)��pD��_���$ ?!���#r���ְ�V�:������jvO��#�;V8�O0�W.?�{y�p�n0U'Н�$�w-K��1Nz���I�C�×HiL�Y=x�7����)�\W$�~�G�MI&��e���}E�^��,+[,��� c�@����Pi�oF����7�5�{�Ȼ��qs���`�a��H4� �1�G]@�u�x�����2yEO'ba)/�0��~?.�d�1.���}�%D�3r�nƎ�B��q?�{@2܀�G���/� �����SD'ѼD#�_=��}�����P3)�yKf}��	�;���?�aiٗ��__}�^
�T�=Õv�R�34�<�4�[}#�* ��G�<]Ƞ�5�t�͂--��󼂩�}�z
D/@��U�+].��޲x%5���`�q8��%��D)zC���+�����	�ʿ���LM�X`@��4�G
G�և�\�i]��Y(w9��Ϋ���.�������a���ʬ�sh�y]Ӎh��T�&k�1��v�����WE.�IY�/1O�r.�5_�Ȫ�ǅ(~Ǣ1Sm<��]��t�)R���M�?�W��h�q�8v̴�I�tFY#��뷖(ӧ$��K����IA}<w2<��H��q�)��b�n��p�~K���a�ώ[�1	��[�VwT�t<ݪ1�	��������hX�b������Jl��CDs��j򺲩|2�Jf�[#!8-�&�A@%P����t *0��7z8%IV6��1�rm�0a&
a����L�e�X!��i1�1�%��Nd0u��hĉ�Y"��m�R�Y���`zK���1�����[ӎ�)��9%$}r�YՔe9qd���\rP#OiG��z��?�?m��T�zA����ܷ�ŕ��,�ȉ=*d�AmG��E*���$������?D|�v�������Ѡ�a̯�e7j@֜��J$��c��	pO?�,�Q��b��Ă��u1��N���W���2��A���;�B�qfBOj�jѯ�� �9�[ɜ��D7̼�axX�!n���_�C�+d�T�����	��@�N�L���[{ߦk�|y�'�
����ٗq�d�n5�t�E�H��� ^@�� S��Q���*�ئ#ML5��!Q��C;Zȵ�"Sϓ9�o1}D����}`p�[�J���^^K�?R��͚��M�+�]��][_��1�?[�N��9�$��m���J����=l+k
���Nk't�4�C��\�{ �2ů���qB��-
yZC�6��ψ���g*Ș��:'��I��*%<Zܸ��x�)�\1vXj���F�։
�ޥ^�l���N�X.��e/�x�C����IT�S��tޯ�~#�F��&B�Wͻ[�ٝ�@һ�N0s���z�h���P]&�b��	�{*�oM�&C��Mo�9(`��|q��h�p>2����>%�ڸ3�hZ� �8,��t�2��'88A�Z��V1���<~`1�}H��E�'�Q�ـ�.K~r�C��%�|Ȑ��+t�R���������D�k�B��x�n���Qk̪�>�4�N*c��������������H��l:�)]Q�.�����5Zy����^��k��}T!(��"��(��}L�i&f��Q���6	��hv(���g�H'/�c��Sm'=�.�P^�l�շ�n��K�G��"�z"��J�P�O=A'ct	��i=��-Sց&�H� ��y�L��ә�����:��+Pd��jK[uyD5��DAX�M}.�L!��6ȷS�#i&����O�-��!X.:�)-�uՙ�~`/?[/4��%�V!,H7S�~i��g�d%�����6 	&'�E���8��e��כQuY�p��ް]/%����>�G�|���j�^X��klf:���EO��YŦ�lc5���mހ�䐓6�����֪/�~ �_���+N_$]09�p�|�J5�����9�R�YY�'Ϲ9��Kg�]Ԁ��A����_e��W�4���^!��:!e���<�p.����N7F_4��}8�DC�nh�Y)TJ���C
�Dl_�r!��.n�YmR��%ӈ�3�W�y�Ģ��A�3���l��
�.V����|�W����W�Ҝ� �X<�e�%$v+Q�����?ӟ"��e��,P�b�n�X�Xx��Y�]R�O'�O~�����d����F>c��s�����D����iL�\�y?.ʐ�H}����Fz������f.�):9��(?��9��g��W����|��'�MUu�G_J$�:�ԃ@�y�����[�䣇f�������s�>�dY�ȯ#v��^�ӵҜ2&C�/����2�"]��3^���i�<yQ�q�1C|��}��/c��H���2��g����Q
S���MNZ	�I�l ��>��!8�'�X���N�h�8O�^C
�&E�c��a�d��"���x��ׄ��q[�wϹ�;���=L�i���C7*��K�~�������}�^�ܭ1�����ea�3���H�D�#lؐ__�R��`��� ��)1L��zW�pt.�<|FP����/M��[���瀖�W�=T�+�'5��?7�!�2�|��9�`�͟�̛�`�Ո��B�m��������gVJgܐ�{��
�A!5�3��2��2�|N����	}��!�M��E ����2h�x	�`�y��'r�h��f����m�{�k�]�ͧ�����`��ZJ��D��N����ׇG^;��ʰ*L3m��-�Z�SJll��t�QuḔ>a(f���5�`;r��YE�I�����=�Z|���1��E�3?����5��rZ�*Rې�����0?b���gB#?��՗��g��i���M�|O�Rg�|WF�K!Zlö�L�_�;�`��:�:�ivfw���k�g{34�m2Xp��!�����qzy�4[>M
6����l�2x�׆8��ܢ���3)H�#��Y���BA���QuBc����S@��S0��4D��[�51��c�9�f�)}��`Ý���AyOq��Y9i�؁�.��>�"`3��`.VYB"��aQ%�@��-US
yq�\\ԨĚz�Z��v�G�G��P �a�/_�|�S3κ:<���@z���(0N[I�t��l��|zY*�؜@A���y��E���E���t3W���h�'4
����:N�K�yw�o��4<!DL��^��E$2Y�Uz�Iwz��R�;�|ȷH��w���EE<⮣S@m�h��c���т��F�}v­����k1Bڄ�ɋ"�&�!��9�����45e�C{2��xn髉Wֺ�VE��,�<�48�2�b6��煂��1e؍��3�О�l%�L�pM�ˀ���� �w��K���u ��&�A�� ���,;����M渵� ��-ndѮ��Ei��Yo3R��1R�~9��C�
/H����:��
�;NѮy�|�X��(�����t�dգ�c~����?�0���hl� df��8f͏l�i8�B
����u��ر�j�ߨj�Ǹ�.���rә����չx�"��]!����1���������z�<��#���65�7�a�W@A��@y*�J_,ؖ��H��_�{�`6�Ūe��xG�۟B͕]�)(ۭh��V�!�׼��b��8(�}����;�!h�6FW�@��H|�e�:@�sM`�%$��(����"�E =%�7�IK1na�g�3��� �1W�iN"n�x����j�#S*T���'&�s�Fa��6z�_N�,������Qڃ�m56��@ΠS��v� �b�a�`����Sy��{�/G�9y��(TˮT��a91 �h)�Ѻ)��U�Q�m��dڹ}�B�M$5E�w���:�^�5��i�r@� $�+�_Җ$�hZ�9_��`JwB� z7&�ַ�[��.Dn�2 U��c��ܟY^h[�D}�!��B�)Ur�^� �"T2�\�}�~���͈K���$�zWD�7y`O�R���7M���'�=��c~ROQE���W�5��kg �]3�>�z�}�G�Ȯ6�\Ni���x�OY��r�^�5�4���S��*b�S 3� >W֮�v����Ӥ����J���j?T4*�S|�<('�1��V�/�҄�C�6p� ��׸:Ճ���唪�<mc�p㏮�����t�y�+j����3Gap=j�T����M�F(N�������~��������_�y�/�_N�]�37�S�{T���䀦���O�)|/�j��-ϐ��>�*�g��B�T8��0- ���=#φy��{�*��7�����
�M��0�8�%Z��f�{\ґ��5\0i����CK"}s#_�4w�NXϗ��e�U���	�(��ʍ�:�!kⰞ<@�;μc��=}�:ʨ��h�=]�^���Z�8��OJ��<�b8y=Q�Q#�?u
k�L:��גꟉ��ʫ�7�Ǧ��'�r���#�QT�s���1�d�0�x;w8$W�w�nk�P�y��m9Cd� a�=,�K�)/���&�� ������5�ƞ�����ό��'�w�������}b�bs��ǋ��d��N/�]�� H��$�T����iim�h,����<C���19��$��}mh]�<� ��԰_CB��h��}'�����q4��4�RD���}�a�T�����|	D���3�n�+���N�F�Ea$7"�msݒR@F����E�X���/u�'$w3��ӚY�\-����/�	G���
v�J��Gt�=u��,'`N�ښ
R�#��S�lMK^���ϼ]ŹOJ�z��RP�uˌwT�Uj��acD枾���V@sI����9`7���8�/6�S������ȸ�Xn��a��q�p� I�R*�߭aU��Wt��i���q��!��b%�3r��2K\łm!��;b��s��Q)�	�c���c!��f�|���d-i���iH�z�z'�BE��);{��B�Y|뷲x��37��`Ua3�"��1�V�nQ�d'a&�+k�g~�f�R��M�X��+Y�MB�I�kl�~�(?��uy�7P�Q?Qjk�N�l�SY��hεl7{]���H��3lI<��ˠpj�p��g�`���i6�!hr=}�@n�#�n[͈��Y�g�C��S$�3B�&�b�"�n1;X~�j��� �j��s�Cļ���6����["S�;��F'P{����o��m%�T��)r�Z	#�"s{ !�f����go�#�+Xe�1B܀\:J�)���`*N4Ϛ��ޡ.��Ns��d�H�"~$���l�[ز&ُ�ى�V��f�ѯ�^���pX��!;�U��U~��d�w��La�\�e�p���W�S4��K$ߙ9%�{���	O��v4�= �PH�4��da��j@:�)+#i�o�J��؄�PZ�`��	�j�E�P"��X>�D���C[;ڶ��9��@6-�fYb�y�/y�xǹQ�����uS��U,%��w��X�[�"��aPG�q�^���nY�7��u濾��ϭ�'��$��0�#�p��-�sH&����g�Cu�y��=���J����)ݭ�v 7�N�δ4dr�s-�eE�n��|�z��[��$��>��&��n˺!ԃ�?>�1^7����|ˌz ����`NȺ� \����t |�1τM9i�+�lv���3B��pNn������C~���&�&�^�Hː}�9Y�˕ؑ�UY�M�*���?J1{/��y��]+sh�!(__a��ڼt�W������1�v1��?��9����C��v�s�����LAwq\|f�t0k�R�b�,��';�/9�̄1����p������V�+��%���&<��,=��󅾾�JB����yF�����10B�Y�"�p��$E�zv��!!�4�1���D��C�e�w.����V&7�0U����7��x�!��4�0����*�o ��ψ���ԴF�z��}(|#�/vA ��X�;�Bg|����Ҍ��c+S��.�J�HW�L�:��t<�(�'���H݌Y�&Q�=��}�6o*��Y�m�q�?��9d�����J�^d2���|�n���ALH2KۮYR�F[T�Y���#�&�߷�7�[_�q$e5��Q�F��Pv���ײ�P��<TTO�	�#YN:��w��O�����s�]d��?���'�����"-P�I��6SG�C���K��E��(N���:b�&> l䈹��!s��z}W�ި������/��V��`�>?����@1���H1��	���<~}��uj?��D`��\�U]
	��v}��X|�j/��~O��Qo�\���[a��x@Y�ЃJ{G��<�B{L�JH&˃=�Ln���%	ob�{#h�Ւi��
?��iL��LAE�Rk�oB(?o��>qaBd��٪W�0�V-����2�|1�ؔT��	_ә�a3�-��}Z����l�� |��<
�؛p8����_�E�����s��"�O�"��\�����;���� ���I(D�5�ڸ~!}EQ�f?`�H�钻u�e�M��)л����>d<hB�t�M����a�~b{A0D���*��B�)ٞ�Z�PO\䣯.���Q@�0�R�
̪j^���}�r6 F!�{l���S���e;��w��I�����뚎W	l�n���'F��ȻV��1�.�Sѵ>�Z��x�4�ԃu�a���s��,��D���eh�֌�w��'�1p�+��6?�%��&�I�] ����߯����*5���l���*tzWE�̤@���ne� b���Q6��R�X?�&����]1�ˋK�=!��nGb�6��)�ܔ�������!��\q?�\�_��v4���c/p��N�xf� ��$bc��U�G��1�O��1�gA�=\�@����	Oė� ���Fg`V;Z�57%�km�Ւ��> <|��i:�k��K���SVn�5�j�Mj�S��`@�}�Ŋ����~���5b��$�F�O�-��r�hm�o���kTCY&pgP'����g�����>�+`����mD|V��b�Ӌ"OY{�B���G�K�����Y���
�c�}<��W	L��KH�fl���,W���o���C���{��ve�x�c�v)En��Ec[��?V��w,�|���
0FC��X�@Ś�j^r��� �&�^z�sʫ�Bw��aFp+XQ�Le3N�kU�w) ��i��F�O=��!bD�Kd?xm&`��� 6��1�P������h_�l���nݴl�Ft�S@>��� G�:�zk�l��]R����0�_C�4�63��Ꝼy"���?J�R�R;}����mP��VF�O��U�V�)���r���pפ�ݾN<�2�r��Z��h��^o��s*esL���V`���#�{+���<$Qm�;V�fp�����)�\���ϧI6�E;.?��=���G
��jk��*�U��<&qۑ�u''��6�}$�N[ntQ��z�5g�1�.����L	�'h=���i�4j�����u��b�,4��S� �����C;v!��ɨ߽b!�i�6bZ܍�]gZK�36����:��;��K�:�Gyo��������ž�;���u:@dF{`cֹBE����v�Yg�p�g��=s{ �z�Z#�-��l�{�N��mi~����!I�`���@3ҥz�4G�e�H�E�Me�gT��"��aV�ٹ��ݦBE���3��J⭖r�e�k���Ӯ���V�{KG?xLAa�� �bf�~�Wմwhk��8��]� �~1�hV ƚ��p���	K"B�-D��`�(�����u*{ת�*�����(À_�
�a�Ue��u�AI�~����]�q�(���DX��Z~�i��^���j�9d���`%�S�"�?��Lî����\�4����O�d}���x�5�X��� �m��r��
�A4"^	F֚a�l���6��u�h�ם����߾O#15y�s�	�Du3'��D@����F��U	=�{�&�G�	G������i�>�⾙�c�_b_;�V8;�<��.���"	�����d���J�V}��w(����%�J�-��'�ˡ�	�NC̔U�a�|Q�>�91��v���&�Ѻx�Ga4�9#��uPx3�)�Ȅ����p=UZC�m�A�CAe��J��6��� qH����A!Ų�g�%�}K�����틐��R���;	�c�ϣrB̗"pO��3�僞5J���狫������R�sm'��)��\l�su�3�I��[�z��[{憤�U������絕ط�LDާ�x/��|��SF3q���,&͌Y��
�ޯ��Φx��+=���������7h�P��C�D��ľnd.�mZ���L?6�+j�;ܾǓ6����>��dm���F��*�2��/ �X/v<-Q��d^y߇bN��T��v��{ܻ5�C��)�lE��Dr�*�KGt�,ϯ����ifK[M3h�0.�X�o��9�x/bl��T�te���������K�[��@<@����&�:��P[|Oy�>���	����[��WW��^��}���F�B@1���"�+RN�O_�V@�ی��/�\ޔ�[q�bWx¼�KX����+1��V��;���ߢ��4�vʊb��e�9c� ��)�Ѣ�$�jL9ZÉvޣ�F@��	[A��F��S�uP������-�Vg���2 I(�=���4�`�jM�:������3��9x�Bw�Ym�nfA��|0K8O��	9�Ԣ+Aq��閇MHc�g/\�C}�C�I��D��6I:ǅj�vv���*�]�ѽ&���E�vkW�'���� ԏ=(*(���?=���է.�s����ġOL����Y�t���R���O�	��g�cnl�C��{1��1@��� �s!ȼF���X�zy��ɿo�8oTd�ڱ��4�S5-���fH��P>ctd���;�lLB?��}���Ö"R�@R��3�ͮ��;z���I�����S�9q�.U��F{�_�urdm�{6R�~�e��=E�{)|4��&�%���;+��g�/��3Me��f|o�b!�_�����d�)��T|{�Ǘ}����)�R|Y/����Ai�&�	��ZO����A��{�?�53`�������1�"]pOv���p$�������]�7��%<�=l\r:�o�ժNeB����}�~ud�*t�������N��"��i� <�,����p�S�B_N4#��7��f4%��Z�+��+ޠ%��LL���2BȦ���$�qY�Bi?�䄞�X8*([U�z��)��An���J��Y7�ރd��$�XJ�A����W��!5XN�ShQ�/�b�ܨ�.�(9�u�*�g���齱��G����?�\T�ɐ��$U��<	Qo���yy��g�.�u^p��q���|;2�,�k;�U�V�H�ebyp��o�̒���~o��t�gy���&D�39s���X����}�Ur8޸��ŉل	�ݍHG�
#�"�:�>���$�nqUuL�O&������M ?)����$��d(�<W�� �y(I՗��YA����w��?z;�e|��x��͇8���3����5��N���q��3<\�-7�!�$�D��kY�ɹ<�q�2/�K-*{��kf��0)q�ٕ1��ط�c���@J���Z}y7��	0L�r)������<f�DCT�
J����B�) ��M�dq��[n..��$�(G}�:��d�8KW������cY�i���LVϸ�o��[`B�}�Ң�K��a@H�[���R�b)c:��}d-���
�:ƈBz5(#���'�t��Ɛ���Ĝb��_/(h�9rN+�Qa��Q7c�xԅ���Lq�(�NiAd�}�"P�}�J��Z�f��b�λ��ӈa�i6m�|H�0�~�N�ٳ("w��q:�LÀ;	>� ��BS�#�.�oٞ��+��=��y~����Yf��+������,-yfuE�:�=:Q�1p�MjoNǛ���jh`�7�����+�	a��X��A��gZޣ��=䖕G���YH�V_�Ī��"O�B~�O�*�[@ѣ��+�7�S���jzs�稀�|����q����O��|��I��] ��ԝtoyF3���=3>�j5��W���j��Jٴ��i9$�A�f.��ȶ�c;o!�%��0�I��s�N5]�\R�+�_3�4`�PY5��d0δr� ;Q����^盀a��
�z2B9��̇ea�E���q�G�my!u쥸,I@҇4Z����;���BIX@�	i���`����T	Z4����L��4�I��P������I�������kA�y�Y�8�Afn���0a��Y�I7���u`�F���a�mt�M����RX���bs�#(���
����\����)|��$�<7})QK�s��}h�����_��Rt����MU��WY��P�(3N��Pm��kF�U���s\�j�
�l�Ie�����Hi��s�F2ȸ�V��!�W˝k�Ѱ{��0���@G�z5����	Q���(cT��A7�ʤ{�le{�F�I�v���qHܭ-_�Q��Pa�X!	�7�0d�o���J�<ڎ��=���Ј�At6�1hw�ndSE�S��mV8��(!����K���"olV�20�Ar��=5կ'�?�.�L4������J~���2I��'X���� �(^b`]׺��4̞4Fo_xgw�/!	������QMǟ{�@uh?�r�2���n�1X�`��~�	�Uj,Rn���W�<ɆWJ��݀��2�����Xr��?i ��p'2	��|Ԉ[,锩@)���0�x����������&�9�_"q��g,����+UB�c�J��!JYvՊfi�j�ۂL^�D�X[�)-F]�i3ʮ�%	�ɂΦjAE�`n@�F���9nv�=�kp�{��w�{-b��Z�Ȕ�:+m�X��Bhp?&�zOi?^%r�y��تVBkG��������%�7Љ'��E��N�1������l/���:]����wۖ����j���"�hC7P���rJĂ���Չ%m&�����ϋ��3�P�}�nS�n��I���Ed��&��:���Cny�e�O�ߥ���ݞ�E�r*���0%�l�*A�G菿7���o<�d�8v0�����
�����Ү⸲�1��Y�����T5�M)X�uѳQ1d�����%�䕪���C�/B�gǧi�����0k���7�gaϹ���S����[c��L${���	��f���ˋo��y�)����@�).�x^�fA�(:�n�"*���2�����ls
��� b���*����^�����M�ɟ./�J} � =�>�\�1_[�V�=L��)�����s�L�Ոy+�S������/F�pC���w�-�P�U##j���u͚�f7Y��GDՇߵ^�U��K
u
���+��RG�Q�g��yp�?TX%Tr&V��d^�!��O�;��	
Zg�}T�r�"`iޯ��U�B��<��6l��
=]����`���/J��W�y_��\J8qQ��0C�Z��n^��Mɳr�<�I���5td��0Ė�j#5���V�����.T2j�>> ���d�Vb� D)m~�L�>���v��q.Ɏ�'N�-E�``nD����u$�����+��)h����1�5P&
W��4 ���L�J�L�*8*ݝ�*�D7�g��(�0����%�#�-[VP�?~{�ѯ[�Q`޴ܦ娳<@����0 ~s+*��z�_���m.b֗U�����W�^l�m.a��fNl'p���fb�͟�K���g�������ʺ�ґ<�β<�\�_��)�q@������W�s���?�\�>j �/D�|Aخo�h`P���n���ꭲ�)�ć�#?��S�ԭ��z�NP �
��_A���6^hn�v�AV�p'<��������c#ݒ�W�\��ݾ�%l�m�T#*maSr8o3"z��-@�KgN� %��0޾ !G�ُTy���fhx�`�谥��bݠ�t���g�x�(v7��	YtH�F�йj��f9�U��>��B�p%"ڳ��qQ9��[��W�:'=�<��oθ��Ӳفz�$�ay�
���U#��c�E�#�m�m��Η�>9g�]��<ka-��^+��'���3�&��1�%�mP���L\�>���-n�nל��+XL�����j�K;�����L�'>agG���]��Rt&F�dvÁ�I�|p�|�>�2)���+1﵄���G>���S�!eJ�	��`��2g��C���.�^(��$�.E�fD�#�v�6��x��M4lt%`���0�b��Z�P�L���oV�� �t/�w��wE�M�2G��j�(=�G{�1�5s�ʜN��ZN�$���R# ��pa�)/����B�y!�w����r�ĳ9;�AC.}Ї�JJkm����ж�SZM����I��>���A �%%���dT��՘b(�}�JVJ�3��m��gr��J��o\!�����J�����|���B$��HΩS�Z7U�ҙ�l?�X�Hqs`Qi[e��)79���/ǅ]��jr(a�H��0��8:Zl��l�ߴW����R(;��P�:尘C (�ZYGa�����Ĵ�^�=8�sb:��׹`5/�)����ik@!��5��ݫ�:�$��y����-ͮ�3���7���3PI��a���
���sGաwX� n�z�(&��)�ǎ�J�i���^�c�<��=z�	� ��y��j�T��*0���M�tXɰ[�����W �v���L���\Qhٝ����#�F;�]x��ü��07���%�Mng>��2��29���ț�^�Ur����n�}
x����&	�5}Цu��am��>K��W,�ǘ6���~�WT�Ֆk�0> /g<���o�������ty�uE���Yi�3�Pw /4z�H�T
�haw���f�0.���Ʈ 9�F8�DzB>HVϔo_7�	�}�k�x�1�.�%W�5��9驗7�u�ǂ���M�m��c�Ϯ삍Y8}��70�F�3|�aOu-�b��Z�9P���G�+rT���(.DE(��o؍X߸ oNV���K�`��Wow�/j�����O�=�=;&�l�ӳ\v��Ѷ[Y��}���4?���?7;��}"��(��Ξ6���XK�>�$��u�Q*�.'P^�f�I	@��q�	?�D)��d�}�)r8(\n��eȉ�ڪ}�%�-�bor�ń�;)�Zz�cl \9Vők9˜�X�F\`G����p�K/g��2T��&2�j�����$�qG�oX�t�c�]�Y��~�x��:�y�/��'F�}VG�k�5(���Lb�-e�������F�JS^��RrǏ�3�(#�fp]�L'@	 R`iU� �!������M�Jn<`ˎTg��ny���HII�:�|�*�A����HH�3���Ő�ߏ���00��'�v���/u1+��޷�H'qb�x^��,��upK�38΍p�b��g'�ӆ��0���,��Wo�a/�13�����،�����_m��P�?k4W���k�9/�X���~a-ʚ��@���K�@�A~��
/����u����V���Hűp�{���9Cŗ䢻'5��YO-#�T�3����X7\�&�S=9�31�T/�cA�m���������Iru��J�B��Fh4�8���w܌��ux m�c+�G���N|5���\!׎޺p��+�{�~ބ>�ґ�h?h��:AV��}�~����V�������utt�5?�K5 ����)�K���d[�f>L}�pyf�r%��z���JqH%[	u���@vbqH���7�1�KB�
�$��]���(F�;9K�^X���zL���m��XF5�U�7�V�b�0��ĺ4w�9����yY@f�R�&�}�|8��"u��9���@$�;��5 �x��6팋����f��l�)�技P*�y&���z2L�%`:�:�����X�"0ɼ���&���Y�r�^hUvf�t/���8R�O|T�og[��s��}d?�!L3��q���L���v�U�! Raץ�Qb�6��ےz�4f��4|j���f��2���;�Bi:��d��Ĥ�t'��z(���cU�E�8zmt v������>cW�t;��ؖ=�w��L�8���~��4G( ��HyO������5oul
�Y̤���}�v��Zߩ/�X���ZG4�4�ۗ2� ��o[�)B�v0��>#s>��ٔ;��8��FJ�?c�>�.��D�>�{�J+nJ�vxܻNb�r�V'21&�F����p_���<��D�3�T���_����,M������6�%s�3Q�/��fsaU���b�oǇ�w[�����4_����1�zI=�5)��#] �-�q�ƚ���>�����K�T�+"��BJ�p�M}F��J���Ў �ن�^6�9��#���v��h��RM7򵻩�q	+d>�C;;�
˿�������V+-?g���fn�/���̃�=9]����n�����P*(�\K�Tw5��/!fm�F�/؀f#�V���Q�;;3� 
���j��_��jj��(�����`�̓V�O�˨��V��fon�C ������-Gu8ڝ�c7�Bf�Aa�*fq��)�%уL���ud��k��4��i���&x�;M�R�:��	�l���!2EJ5���<�˜sӕg��1򆬣q���	 a�:R��r�r`X�B�,	�ּݞ��;2�
AOɠ�ḙH bL4�j����m�s4��4��N��pߒX��P��ʟ!���5�|S�����Q�=[=��ZUG��V����gUWg��"�>�GAO�j�UՋ����%�D������,��Axk@$]��'�u�K��u��i�R{A�t�E(*����4��0�������}z���Fl�▮S[��l�'���N����)I�	��p�OdTɦS�*�圫*e�����k��jy]y"���U�����g����Dr�`�e�#]�Z���,��8���j�@��I.�Z� ���䭖$Y.�%"ܜ�
p��(P�.��2=ULUo@r���-���T�<t#}�����j������I��Y_}�#p
��mQ�̵�U�0�¥����B9�R���_,n��g�K=�TM��|��}-S��.MB*�ץ��N{�����D)�ĕR�x)�{��:"�v��8�܀�]>�1>���d����/�uLn#��z�:{��/pW6�#��m6Ar��G������՟�#�*/�L'΀��CY�?�{���kz����3�U8ga�S�����}9�DD��=e�M�/�G���z�t0��|a?�ib�<E�O������,��>�:=螸���K��N��ŏ�U~�V1��3bǇ�Ӗ1~�0C5X�8�6R{n/�i�ĉ 웂_��Q��TIEC�����ƭQ�I#�խ��3*zˉ�����IX���)�G���Ƹ�B����7�v�1���u{%�tH�WU!�	���0�PxD�|��p�06P)0���M�T6N��?U��Y�������Rہ�� D��nճ@2�C%�W�"�r���� ����Zct�C�DU9�7�i��@��8���H�,��d���{�H[���f~��v����ƛxEH;�%{YB�t���(ϱ�Yy�\�(��[p�6ݓ0�P&4h�7�r�"\ W�H�W����g[�k�w[�Tc]�����?Gc����d��[���{\c���(�[���d�ώ�$,ݍU����5�z���˝ƙ1����=�3�u�?6���[��t���2b����Q\��<⣋XN�ؙ1�38��z����Azٿ)����!i*�?����"����D�G�������Y�_��L�ө�}���
+6!�3��U����+��n/�'C)�좦����7c������l4i|�����u�m1U�	'X�U�ʀ�h|E�R�r̮�k��h�C�CW(@b�wu�R�b.ٰ!�l�+v��0�UD=QY�ܰ����,��Y)xZY�@��Vu^R�1@���݌�z�ѡ�c:�*�y"*�~s� �acT�ET�\d >�LG�n��1�{�c���n������m��qG:�ƭ~RmG�qu��Dȅ������[!�S�X[u@��C�{^^��p����Z#�����x�'"ޚ��Ll���	&��h�����������+�eF8;T| �N?K�]"5����y~8s���]����q�Z�fm������>�D���67.��:�z������v8^��J��
]ݙ %FY���A#n̊����k2.]�Ids��F���=	��ӓp�����沂����L��c�ǜ/�S&9C�G�D�'�gj��@K�k�P���>h>k�)�hI��4$6i���o�˄���	�ת�U��pn<X?Xe~�P�
D	�<�ޝ�t���I��ų�/q��I �@�xsd����j0��m;�cN�>xޥG�H�]hDc�=\F�5���:�}�"+�tq<Vg��&̜1�C�a�=���+�Y��Ð����� y��9(��I�ԔȖ���+�G�Q>��:ȣ�^��UHT𭦽�h��l��qٞ����[��Z��͂�{������Z�S
�{�Ef����2���2d�7�}L��YF莅3T��� ��1��Lo����aȆ�Z_1&�4'��0�tMd����gv�����Lv�De61o��R\ډ�tJ�<Î�$9s\����sT�}r	��Sڏ]`(�\Z_t)ʻɰ�r<�U<P?a��㷬��#˧\�)�eCj	O��Oo��˩�D=����,�!��LM����[�!��M�z�+Z_]Q�5[��RM7���4)$�Uc<���=_w �$w۳gQK�kT��<�~�6��[3��\!�3�R����ݞ���A�ͤ���%.�1�R�x��	�\�� �� �����xa� +@��Jos/E@T/����=D}[�qs>�#2X����V��y�U�<�#��nə�� ǋ�m!��Iw��
3��Ir%��U-������a�j��;�P"}�!FE9 T�,0Ȓ���2�~>J9�V	� |�f� ���I��o��\׍"���h��v�2���ֲ^ǟ�( h�]>�r�g���=��N(@�M9eˁ��
~�qӤY�7�OQjv���HK�v@;�E�6���}�&��b�?{�� �*i3�b�0T�϶f:�c����,��.Y��ыwpn;��Dve��$����T�ή2B�H���s̑y$#�F,�����n����
�[ҷ���u3���̧�FD�l�)���EAl�U������|.0��N:3��
j�b\\�[iqE��=���jo��8;=y{1�Z����?�/�,��4�Ւ�+�ybt�qza�_v�9;�x���q����5�bfv̹:�tF���-����0�Ah7��JT�� �*�h�1 ���!uX#V��}�t �-g���՞Fd�6��8|.��v5��(��v��$|R�;K��F�!bm��hJ�]���J�L���]b� tY�����i\��q�	J )5��7(lc#�fϋ	]��� i�4�5�CT���>�M���M��t�Xk30� z���Й]o��%�HT�o7�}M���������Dg'������%�H^��C3�P�Pr�4כ�V���;��5�7�ƒ����m�)Q+Kw��9<ϲ{%ړc����|�BH_Rc�������eN2@	����4my����0��D/Kz)
��7�[�`���Tu�T�(.~�tբ�e!
�.o�'r�?����"4���-���LEG�tД�����;[R�50��h�S��,�n�L��[���o��Q�Atmq}g�u	�z�h%Q ���g;�\9gq36�)��a�亦��xN�'4����?�6�.�S�p�4K}i�A!�4�.~z���n�0&]�W ��nW��b��F��%�q�2��*A�^� k)*�M����-�/c�*�]7�a�Qųk�ـ2�Է��i���X�*��ݿ�"A��rt�m�����I�u-(BF=�h[��b�-Բ~2e��P?��/��	��&�<�#�k�zZ2r��}��N[.����s"��3z����gz%�~׭1)T����H���f8�8zyT��y4�5f��=��K,选���ۘ�Ճ.N����$���N�",A.��,|����?�)!�e��������@ {�_�k��5GT݉�z�ި���+���,^��>�Ӫ�6��j~�T�|�jc	uM�G�{��h��y�>��š���n�g�$S��,�&0�j���Z���l.����9�a���gd;��5}�_/qf-��u���8}&N��ߤ��f��%�k��#Ш)K�7��u2Z^B��v`�7& T+A`�V�ж�d�9���{�$�ʃ飰�"��xx�L�t�¢@H��3�F���y�c�FX����=.�L���^��RW/-RX]c�=9�h��zY
�Z�O�2�M|������5\�%�+�c[���V$B;F�n|?�B���uy�Lc�ڥ��@�/�[��&�2 O|k�J�{�!O�~�8&o켦-+N�L��yTNTE��V.��p\xz?>�W��:��u�n�̯�� ¢=M}�6���p��EW �h>������W���~�
�F�,�C>B(&%F ����'�j�U}��v�$�M��m~=^��:?+��ݚ�.������ִu���t�A(�qϟѺ�-�F���%���7��2��"�N(������)r�\���������Uw�WM���ڜ��r�m�7&}�@DJ��_�o��{D��P��	��Q}hK����&���Q�0���	;�D�����-C5����:ˀ�tK���-�I��$P"+�����S��+n@��m�˧���ٷ�T�5�2h2ˋguN�"�+�~(n�F��b��tdlf���Ҁ��I���g���W0]�s�0��������~(��n�MK������[j9�p����ɛ*-Kh�%X��TAQ=Po4v�t��3���:�����\��#�23�1�5 ;ڡ*#�jUa?�:�u���(��̤�(2�ma;�!>���ׄ�D��dH�-�N��e1�]![w��XM���l<�1�an�
��st���	0(u�E�!Ľj�x���S5.�v�)ĕNf��~��~�d�8zC*�HO�G�o���v�4p#����|��;H�nc˦�'g�nG)��{C������?�� ��E���wQ�o3U�Y�L{E�e5M�RM���)�0u�u6ۅq��7CqLCy"[V���r(Q?2A�����l�����e"�yNUF�Y;��ȥ`/�U��代҃�u �Ӯ5R�D�	b�@�����zUpO���%�H��|�\P��ۨ��]jGɨk�I�EBH�u��3ڝ9D��>;��Dz����;��V'-ŕ��V�V@��h,�)!xGC*�}.{�U.�'0�L��;��{Gx��.�u���`�pj�>���)��Q��z*���$ݎ��J�P⼼cPL�]�������=G��i����!���e��g�s�ȩ�<���;�p�?}���U�(��Q�"�t�����:�Q�t��H���&I�����C��eX7� ��fO5օ�����@�őy�2�9����+����`�r��g��k��8��lLwv����څ���S�3W+��hiA���4om��i&�LOPr�,�g�{��4����K�h�"ww(�#U��\���:d�K��7mY|z?�5S��W~A�〼��12U�*�}͙�΃2Ýؗ���Y���ߝD;0����L|(r2�HD����7�xp��?�������4-��ş���=�tSߨ)��&=���glh'�TR�n\�~!ZǗM�g�c����E��&Y�3��e�<�5�3pcӁb���R���J��a5�W���>,)�JlJ�E�o;��BTr���dO��xPɗ�ä����=�?���P�B��g`z�`J�"���#���Mҋ�LrP�ë�N���ؗ����@.i�l���]�:�,��i���fC��nF#TQ��C���yR����-T]��?��呥�\�*���lca��0d��HUJ�݂��r��U�^�(�Zr,����/�C֒���qA
�� 
dyB{g�`��L�����B�3Z�&v��u��sO���E�F.�!ԙn~��c��C�u��^��&�)ր�h��uh��eY�9Y�9�
r�p3ܾ�N��Y �e����d�G�H��o�~Vmş�1�X��y��|��.����E�M�W���I����܉������%���y��:`�.��������k�9��� �Yk5�Y��ī�%;v����PH� �FO�uL��5�mD���� cu<��Al! �AL<�;��l5J]1��lW�y�$*3 ޿�9�0	l��J����ٛ�I����W8�NuQ�P��,n2X��vw;p����):�OP������=\��FK{j"�0񎈑��a�m�4J(ԌI|N��ᚔ�����2aާ�q����X��9|�/�3��'H$��j�M�PG�����A&Q-���.����M�o�f���.�	 � �'������n@j��.w�2l�"�
��8~����'^D��8�SFt`?�ϤFN��]"�6������7�/�a�$�h}&�����OF)� 4�ƣHL�G
��ěJ��_���W�e��pI�*���j�]{d���+,��o�aT��2��(���*,z{��0(E̢x��,��4�`(�=�9<FX#x}^J�{d�9��G�Ӟ͇�׵d���N��i+�0j�f5�����|@H�/�²m��[�:�}ni��<Fw&�x>Ag�NKw���N�;�oUX�Vm	��L��mT_e6���*�L.a��&_�����*cN�F�;E�b����>"(Dq\�L���I4��#��At��R��*,��.H������v�|��7C)�	E�1�dB�߷��x�b����%���3��ER-{���sԤ$��
~4�9�HS���ܠ�cϵ	�3�Tv�����3t���jB��֢�(�

�&���<#NOZ�Tj�r��H��2(�=���ܹ4�3�%�	4.�q����[׽�q�
Di�		
�6G�*��vF��������i�Y�ؗvt�_���f�&������1���>Һ��v<���,(�\����5d�z~���� �]dXPde͆T/f�Ӱ�8��)��������UcG��,�M�j5��Ē���`,e��x泚��@�1�]��������{ް��ۋI�Q��K�)!t��x��*x����f�/�!$�!���A(!��D0
�z֟6���z����g��	���Wxx g."#�=P��2�E����э��U�=�%��
L��"e�Mp�b�3Y(qϻH�\B���zl�����p�6�6h�ԃ�o';�IW<����Ÿ!U����f��|�[��T7��������P� �a�W?0y-\��qB6<��J��^����`��� 8f�3W�����Lz ��t�7{���*�ߛ��8���F�O�2z�S�u�O\���R���y��Q����L[�	K0���{Fb(%��m��_�u�L!�hGC��eo0���pR{yBJ�`����4^��vW8wZ5X�(D����g��tɪ��L�V�{�T���������~��݈�q~kR�"G���ߩ�Q��>���I����d.��r�R<�/����ᤔ������^e���z*��X!n)_ ��D����{�9��Ժ�a��)�~(��-ս�Ђ�9�(V�@sB�ӱ"r��D�K���.\���
��Fs�	ɬ�}��-�s\^cd<1�Ga��m݆ȬP�#�Y��ל:�C��q�P���	���ha��;�T�.���,y���j��DNHy�3z��$����@l媲ϐ�;�-��a�pF&ԕ\e,�"�a����0����l���xl��n�=l����ˮ(����˒���)�v	(��m$��[�<?lX9���=$�Z꘳����y��7YS!q��n��G����rb>���\"��?�}m���m-��
�^��m��"�������aw�2���j���4�cBbI�q'\= 0&��6�F;��z��"5o.=㱫�w,��m�����X�L~`W�w|���'L�0k������Ĭ 9�Cm�����D���������TB�v�Cs���y���>(lǈ�`�fw�m�pt�'��
�3��+��3|��ˬ��"�T�l�{���"
�z��63,lG�+c5�\�L����hHx<�Z����fyт��m�	���O{�!�:����G�*>_�����6��T�^�A9bt�1Z�vE�/�=զ�<3e�q��k�
�h �k,P�c����n�P2�� 96J3)��14�Ȑ��Jޫڼ.�W���Gi-�ܝ(����O�C��˒�?�(	�^ͮ���/6{1>�~Ot�(�8g��9v#'Z�g@7�d�~��Y�f��KĂ�W�n"�>�v�Ο�;�����RYjA�y���ʣ����C�i��0Y	�~�o��I�WKn1����)[řĊ�_z�kO[��3o9�z�3�z������C,N�٘��F�]����d��^���Nsx��G���lm����'/�KCJb���>�(�B��T��U���ۏ\WpIZ�t�|\��57�bb��>�$�R��H'�ފw��q����g�/tdxe����bq��>p��]�MHwf|�c�&���q,���$z�֪ϲ��?Auڟ��Ƅy߽v�((�Z�J�������w�����ڸ��V1�mD�X4�cNJ��6�K*��'	���u~it����kpꕬ�8;	��A
)٭uw���̦�����A�1��y���Ggd���X��ՆF�K���ߊ���L��^�#1�Ly+��emW���J��)OhD
GD�*�Z,���U	�m�m?h��(���\�[N ������<#�iΫ���<2��UHkN�7v����mQ)K{�VZ>�G/n�)�R��/tn�`�$Y�����߻*-���Ѫ�t�@C �o��۞�[w�#ʜ�X��2<����.��]�M�/R�ucM��$���O�Jl�}����x��޴U�y��M@,����c��]C�hD a���*L�q��Ⱦ�� o�/b�#��F��q���(� J�=%Fa呠��+ Ϸ�iY�n�:wՈ6����BP)�(�b�gi�~��]���˲���:�ʔ��rѵo����u��A������E`P`�z����ʾ������,z{e�����Z�a��V��N����/�^�0����M(i:�b&����E�n�������2�Bۤ	��W�c�s[-h���&Az���`.$�)l"ͥ.��+�(.@+/JW�/����A�>L#G-��4?�;=��Śn��0Ӭ������)����۽�b��b>�o}_��T�+�Z= g�����%�Rs`S�3-j�=5H�H�8-v���ܼC<(�D���V9�UMu����R[��sa��M�H�ɵx#����J�ޑ�G�r��3'�$2�z�L�W�V�5���k�a����r�j�t��e���x
[��q:m�����^��USiR+�$�����-$�Q���;(����*A�&k�4��;�4�V/;Dt��G�ٸ��Z�晐�s�q.FA����U�7'k?E�|�&��G��a��3���ږ���E�g=y�SؓO�B��ӧ��gq8QQT�A�3��Ԝ�Ց�� /������I���m.��# \įk����>FZE������<~�Y�T�f7jqg��Z�-�
�(U�������:�&� ��G�Ri�i�&-�7������YQ���pyz�	��V�)��R���h.�N��ޅ.�S�p�l������=�Bz�%�ʌ�,/A��
S*�zؐ��G�)n��/��qk�����cH#����"��[D��M�\U���٫R��MƄ�y@�n��L��so	���q�|=}$:/��M�w�V�aW-�س�p9LH՞�ʖ^���2��]b�H��l�;��/��[f��^24��2�7s��0�:�q_)P�C�ė��$�5Elz����wO��t	��o�C�{>3�����i�bJ^#ԡ3Gɞ��S��\�9:�g�J #Y��">����b��Eg��8W_�7:�KN�
ִ�A����@� �	Hu�T}'��M�y�4�ob�u'���cw�����k��kKqTBx$fu����o-@I���L���t%�c��KҖ�J*2(9
Ĉ`4A?�X�@RUO}�������Ԇ;��Q;G2��X�6�i���Z��yF�z�rH��aU�K"�!�&�y�?��q��K>?#�\[h W�Z��Yʏ�\)&���eЉ� �3�H}�R@�p�G$�蔨أJLY;8g�4V���ԝ	�0���Z�h���}YG��Z/�C�3�ѭ�� �&[�?%��vل�E>�c%뎋�Z�R;o��]�|��"�7.;��n�/�M�J)+~��*�-��S ��V69���xhX��T~N&��w%���u����؟���@�q˷F��'I�w6½�ᤘA=4�$ъH%��a�Y!h��e��b�g��|���Q"�I�)f�Z�3P�6k^~q���\D3��ܳ��k����g���o�U���,��y�˖?�T:@�ÿ�T@<��c�xs���\��Eh���sd8��V�mS��a!f����Pv?fo�kE o~xf���e�,�5��C�,$�n���W�'Ɣ�I� #���Ǹ)=�k��;��tϋX��В�4�S,7O��Ԯ��Џ��+T2ȩ@h`_*O��n�f%�ڵ�L���c*���=�ɓﱚ��K�T�wg�
�IH�jt�x#ǣB�v�K��k��h˦l�Dti�޻�J� ����h&u�,j�R $�w�y�Ǜ52<E�&��1��9�#���:y��q���=�H_΋w$�4#�{�(S��>�{�=�������K�S�(�<Aǃ�Ff����dr��͝J�G��!�,R0��SR`Ҥ�*�S)C���,��R�X��ʘT�����l���b�+�@7��¬X7G;�,a�\�,��#���C;�&��`1�#En�^�XOrV�^���⻱$տ�!��W�gW��jB���,�S#a���ߘY���O6=?2;;�騱40�n2iT�8���y�Ôy˓���&�� � �;�j�e�h�a�K�l��'R1=�I��A��R�`TR��	&~ĭ��������k���� ~~z|FQ�N>;�h�`o �G,�݉�L���g\K�j�6z�+�Z�7��s�1)�[ ��eW!��D���G{8�􋑢������}2KR�X���Q��l��X���.C�#��Au�s�К�n��V�M�^����"Ob�߉G"��dP���l}Y뗵숟���*���*DG�\�67�3��^R�n*�y����,[����]p���
�֊ŏCA9L��1M'��c{��ZׄM3�2M-M�!=P�+����IG#�+����G�f��o�] �R/��َ�ŋ]d�CU�ծ�ߜ���#g���䩉i_��јYB-�E� L�����QA��J��V�����f�E�nS<��\�{��:�9��ҟ��+��g�2ȲN �-��^Iò<ψ�t���pܾmO�{I`JS�[,�@؍r8��rٳ�y=_<���j!���?3�`ȑ������D8����ъ$8
\�]P�ҋ�+��_����-<������M�s�5���L�V>l����^'�nݘZ�I�a�ģ��h�{Is�h�cl5�a�$.4�c�2��A3Tm��A�iq=���`'>�t�t��x�(��l�����o���"Z�[�꙼�f5Y��^S���D����K�^f�0��/��kG��!t�
��*���s8ߊm�W�
���})�O�h<m�Ų牏�UP��,�w�~ֈ��Q��v�(l9�|�"/�K	�d'8Q����Լ�����.J�UB������M�U%�a�����!�i��������Q揜!��3,
�<��Z$V��$ƭ,���m�<ޟ�FƩKn�n�YuX���$�cv�ՠ��E�8z��<�)��D�q���	��h�ߕbXC����U��Ou�r��=��{�ϩ;$� ԍ��r�
�U����5'J��I't����Ŧd1_m��]��	2�� :`gO����p%z�S�ت+�3=�Dh�+���ʴd��o�d�hʷ���}j\4Nu�?	������uv��J
��Ms~��y'�(��o�|��X�ِJa��p?qǵ�W�����m���!�`'���i6�Cd�;�H���&��%�F����&u#��_"��9�?M�F�G����F���U,�xz��s�hUB�?���uj���������B%·�`j��?n����\��yo�F�$!��3�����J^��!ͭ���� H\1�JɿeH�	�[���G�Y��z,ȣA�.���OD�0\�l�I5�Dp\]��������KO ��^҅/rN��{�������!ps����:����UW�����M��U}�����C��E-�Y��v�V὎'g�	S�%2iINa1t�����VC���٭!kf���s}���5�(�4 ��� ����_�������c(�!F�11]�/��U�����41�Y��]��ϕ�G2�DD�aIޘ9jb�_�pG��I^VtB��mW ��݊LG^�0bɵo���0%����r�f#R�j��#n���O��0`�=�5��Z��B���3?3��~�B6�@U�j"֠ )�F|?y�QI��"��>���x��S�A�C:Д��2������:(�=�*Dp@JO�$.:^���`;v]ȀA.-t`Ұ	�u��&���$0�)e |���ʫ���M\�_���Ǵ�b$asb͇G̢
�KA4E�R�zm��NA����Fۏ����VLOخ�v}�dl���M�՜9�ixy%Oχ�&�N�w�D[�\�*}�z@C�'�8�������� �{�^V����!]C��r�^��������R��|�w�E�f�U�s>}��x͏�Dt/X����1~��N���9��Yk��M&{4�D���&���0�a����~��/>�bO���F|7t���21�Q$��/�kuMb��C`�$_�	wCel��B2wԽ�]���|���- �$����Q�����N�.�TnO�8C!�'�+���/�nm%'� ����o!=��
�����?��Y:o������`k�˒/Пc@�L��OߖwE'W����^�Fw7�D���p�������$@�>9�&��kƦm%oXs v��ψ�Ǚ��%~��Q���H������� �@]�tтcgE[�ڪb���Ue��zLPœ�z�>��Y׹��1Ɲj�`�l�8{�q��wq>ț�<�%����q�I<��i�_)��y�0	I?I�г�I��&�}�,0��}!e���\%�[��S���J{yWWk��I	'���W�JD���$nl��] ���aK2��@Gi��	��\0��li���_����A�g��S�����7�q��w������64Nh>������>����aK���3�V�7ϵc��@�͎�l���i�.���I�C�(����sCV�`n	��TX�ߝ�h�5��9Ȕ��őp�G����HU�)��WC�wr�o�(-m
)�� 4aC���R��Ȯ�V_F$���b4Hz"�FdT�A�܄�KZ�Kl��Z� ɋA,��E�CȪ���N��IҊ9}�̉]�PJ"}�C���@���{���ڛ	%��I�L��b�Ǻ��`��ǖ�̯���t��K��O,�ځ�Bm�j��G{7������3���S
�*�[ա����s�l�7�٠�k���-�����Y���H�h+R�*m�������v>�u�Т�;8�@������b�6��ҲA�t��͝�0A3�8���	�P���s���� uRj�a�o����I�J��<�00�.�FPL`��AF�X f"����6�~jDGy���`��R:�0����l-�+�Zԯ"��Bx"xܳ���:��$P6%�J/�M`��x�	��~u�20�*��@sX�(b�
:qhonୣ��(I�*��!�z���R&�M�שO֬gh��}1��!����a�2n�fI
����~��Ri�(�2lz.�e`�d�("��<���غq������0��QK��� �l����-`�v��k�SZ�t���;xi������jM8�?��?��
7or�J֩M"�e�m������������W%��p��&��
4W_��:�	d9�	m��5�d'4����s SV�G�(��~�n�M�����՜Et�N���<r���/([�'���ѓ��)�$�W\�{Q"ac�7Yz ���F��c:z%ݯ�3`}���Y�}��k �N�Lx���]�j�<��y�8����ۏR�����@����;�s���g �1��_� �9�U�i�����t�,���,3m��e�F�k�Fb��*��1��	�{Z޳�͑�_���M$ i��S9���-�]�xǔk������%\�"��B'8c��&��W�D��FR����!�|K7S��/�Ogh��(���?u�@�ޑ'V}f���v�N�D��k�V�&��j2,}{�ًoVd�.u�%��F�uͪ�mU�l
��Ə���㖗��n�o���.�����t5�;�;������w'�O�u�H����\�G�e���e��<��/�)��P\�E��}����(�;[4*� ���I�H�SOp��2@b�QNG����CHr��H��H�@pa���?ЏBL[;�(�`���A���6)��M�s���6�)���(�Knkx�+�uւ��a��1��M� G�䆥����=�e��É���J�;�~V"��o��=�3=�=�D@��Z�c�1�@��
����$A� �V�>�|�A����|�>�~3.G% 
�A_;�(4�m����1xǨ����;�M�^����� �l���-���Ԥ7=�k����x�e���r;�ٲ�����QJ�>=��l�y�v�#��a��0�v-�O�tk�a�nM�v^(����&�Z���Y��Q䘒y?@@�6�A:����<����E��g�#���x��SU�ю���9�h���MYSI��cr�C٦a�YVG��l�5��zW�/A���r+�����XCCC����÷�@"$��V�Mhp�H��}���"n봟�ȣ�kPn���tH�>��E�&"5��IY���^���\��p����4Ƞ�W[ }��E��1�,�r+�%����֪m
KM�~aD=� �k�S�gq�]�#�C�@�7'��)���
ԴM��K����I%�IYL�/�ŷYiV��;?o���}��
�J��t1��((�,ebQ����m҉�j�Sd����j0���Z��+���l=�Z/��4b+
�h��e���+W���� �������7 {X�3��J��[���җ/����"?�f'z��7q�����c�
���N 
���; ����X[s"?����W��^t�eGw����i�"�Ӯ8+��ڌB� �!Ԕ����ȹA�	�?2��"-'����x��u1><��J��J�Q�Z_���:2���R�R�2K��)w8vg���%k�R,Q��ktf� ǻh�����8e\1�m>���D_1Τ.ޗ���d��ª $�PNw��B�V�k�螀L�<�M�����	����l��t�U���8�X�w�>Hb�bs��[Sw��;��/��sP�`��C#�.��>�������+����b^xԎ��9�'E��U K����~�1�!�4����{_Y���r�W*�1�c��C?�$�+�k=+~���Mhh����P�~6�5i`��Հ�R�u��������_�s�su�n�G�=~�u��?��_:S��O������g3����Z��"��#���7Z� #��[k����A���1m�~'	a�S���m��Kldjo�d��Jtɷ��O�e0E�h���~6w\��6G܇//K1ʉ��2"� 7�Ju5ai�	�ѫA�]���	�D�=)иJӚʉ�T���{�� Av��|8[y�0|�����:����
�&���6W� >���x<���gL�7Cп�O��P�Aն}h��v�,f�&|�i�a�,�"�Ac�����\��ǁ�	�F���=����,l��Ү��H� �fge	ٗ�q�J�'z�u���Q"J�9��d�B[���D��X�a���A6u��Σ���{i�r�W�Y�WF̈́��d�[�*�{�+�����-i�n皂�"':�J4C���Q_jT ��z���AI��@?� �4M�������hc��٤�o�7_�Q�rS�~^-1�N$�A���XFh�i	X[1�9��@ym�#�
�I*l�/H��..<)	Q��b�gT�V��CA>��~iR!����O$T���M��;�d߮���3�F,��l�������(���I�S=i�Hb��n8�m�m����G��^��rd0�=4զ�~ڵ��vX[��-υL�S�`��}ekM����z���y��-r6OW,�b��(Mu�(Ȣ��F�/ڍ�G��)�]�6�ެ�j"]�k:��"��N<��O���b*�����v��u��I�3 `T�$V�K����'C��x�5�9j_3�i���� ���2�ֽ[�ji��G[�M�Y�1��At�)A")�E]���/�xv�fj�R<9��heuJY�g7������[q�Сoov=�4�y_Qd��~�tG��)�{���0�QF���σ]�\�V�Ǒ��/��8Z�J�]}������6�~��*&L�ٰ-�Rg��������n;"�	>ZK;G�AK���������r!����n�
[p>�Ҙ)���19��`�d�zćB��y�����͸z�p5;n��0�J+�9�D= ͽ�_F/��?)�#��/�k�y4�i��t��F8b�*��(�K��vesԲ�E���k��ʡ7��Y��,����.�J�vQ�_���ؼ�y��^�2� ���gH�[����yW3��^w���P5[|4κף���d�
�qd4#����\�S�熀����󗐕ࡶ�K�\/�fI���R��W���N��8���}qv�7QF�/g*	Y���e��`=N�G���P�-��PF������r��|����(;;6�c�ѓ��]X�xr�ڟ]���  ZԐ>ZҚu\A��pA�~&@B�G��a�r���^�Bψ �r�B�f��NV�gw�=H�jE�J���$����Q�4,{ňb<<�m��3�'�;��5b13�F���PO ���48�mv��7qkU��+�V���_C�����UIc��Q���ٺ�CQ���yO��X����<ʢ�Bt"�H=nʽ�����m`{�37���i�ja}uAd���I��D��+���9c �<J������$�A�=�M�pm�_���et���b6p����h���'5h8���N"T�_إn���v��(�ы��kƕ��y����I���ȟƎG��������a��k/ރX.��)���`i�$���T���&y�]���E��E���P�)��`��p�ˍ��h�����<�;�Qj#��ڮ�:����qm;��A��T��I<����\P��D����(`���/� 2|�İ�}zy�p���|[�-R�l�����'%V����?m�����H2 ���6fx�5�G¢?�ϴD�=lf��s����*C7p�Sz�f�H�J���B��o��p�t�C�pm�{���Ʒ'��qT���n%��Bj\�D$��qĵ���]m5v�~b�d�-�B@d�=�X� ��<�暧�:d�F�P���U����kѨ�xb��7/��*�,�?E
/*�(�u.�K�Jt���ߤqLW#a��|1��H���<��*��ꥪg{�L(D����nNA��a�蛓�������dT��l���1�I��!�k�f��N�9���g'��I��(����B�n|�yUa��4p`K�q̢�
�_����W����3�Uٸ��J�E��4T����&w2�����J�ZI� ��F�9���O�s*fP'Tv� ����˄*�bN��K�����2@kd��E2(�(؀"�<��t�e,P��S�g/⣓����F]Z(�xw��eYz.����,(Y�6�<P��I�L�v�{�`u�Ht�?�n̵r��:+�1���"��u=c94�Mn	�1������K�G��B��@<0�hܛ�<J$��;-����EoAq�(��W[�̚gճI�B���P���1��4A�w#�Q�f��IHih3Dm9�03#O�D��=@WwX>��_�)l9&�Y��xv�x	;g�����f-��X��T]Ul�eʤ����ܫ�e�Ȃ��n�;wh�!��|�#��iޓC�*��ڨ��̊�W��@ʺ�eB�Q��q��]��� ��J�`�-#�#5sh<��~z���V���-큯z���v����_:��ї�5!H��c�IH��wCEdX�}l��Ŕ)���Bң��H��G�Z�u�W�eE�x�Z�h��_$�+�Eh߾��i,����e������	U&�x�D�L;�.A�ࠃ���H�����d�CD����W�1�k|UC�W'�'�?0�Q3l��w�
��IT����{��mM��Wq�ۛ�".4�xa���?PU��dY���:��ta�OLa�³�.%�S@k̢sQ�k�+���I��dr�0ߗge>�iS�ǌ��.�Lnps�^@w�z賐@��M����g��C
�	��[� v��;#��^��n�P���ڹdF]0��8�A��?z�yp}�)r�WCǧ9
_. ������I�>�W��ㄿ��l9g�?����1����LK�K��4Ϸ/��A�b���v#�z�1 ��J��"���B+��*5e�
���c�@i��Wע����;s����3z� �;$w��>c6ǰڳ�O8�}��7"����Ӥ��u�>�Nt�n�_�jRN�2�&"�c2>ώ ��4��[�����	���7��E/���mO	��*���S���`�=�FB�d[�!��Ν��_��⑟����M�^T��-Z��r?0�߆+ME�}܇�J�@�0�U���P������T]v�^@�Yz������+uB��4P���黋��}��g��ʂ�f5S�(�c��׻3����!裘�xw<s�����ms)ɦ��q�:&���]�}���u�K�e8�Ԥ�(��?y�%b ƫ�4.���^0��8�)�G#�5�PV��]�QI�UͥN ���G~����.�;L����&�Z�d0e@�rHgT*����p��n����$��ARŰle�n���.4f�+:����,�Fk<�kĮ��Aڜ�ߏe�?��#�w�g=���TYV
�����?����tBI@�i�G�y '�&[��kD��