��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u���/�m��,_�v��kH&��bwH�p�ZC�P��ٙ}�.�J�@��*Eu*Uc~�ߏд���Kږ�����H�X�d���U�����f�Y�f��ts�Q 1�<p�
�Q�����n=��7�+;P���l=<v;�ߣ�:GD:Ή�mq���I�s:�j9_��U��N��	A �#XZ��
H�e��� f�ZYP,����0���k�)�ߺ���df,������4�>�H�+�$�!>�����戽�3�rC`9�=�;B�^(����m�Y��z�(ߊ�L�h�� ��5�2���B��K��R[����&�)�^��VV"Oafk�E��B���:rk����cB���\�! �Dpl7��0�0�����[�#����	�r=r�ok�{��
�`�*���
݂(��"��ϯv*a֑���l��	tMų��.��7���UK8�����Ш����!@A�B�`�Ĺ,�|q#ŶX�%�h��%�{ֈ�%/;>/�#ׄ~b@�ą&ڏh�a�����a�s��a7x�Iڷsz =��,n��# X96o�A7�%�nR�)��$Ki�d5�8<=x��6<�U-�����J<_�Óvx0����;�$�%�m~s�$��0��V,ʹ�{^��y�]i��{u��p¯Ȱv�$�\:�D��8�ٺ��̊��6z����:�. ��Q�����PE�8���&�6o�̈́���P>Y�Uc�6~5앒.f��J0�b��`x���d���Wcc�G�u����0�<���1B��u��\�6e`.�-{v
��i��F=j�����sS�b�mz8�����ά:��o�H�e�b�r���e��|I>f�bV�����G҇Y��0Ǎ���|&o�'"s��[ԾXC/�i�2;���'"��@�b3�X�D���c��lñ\�D�!i��t�z=Y�ae�I,(z�H5j+�n�}v�C�"&����l�ۮSbe���v�5��Z��:roWq!�J+�������t�mfc�.y�sG|K>�0�З�x|
ߝZ�؆(��_5�"��mԟ�mk_��qx�Q^�b��@SCJּٞH�[�-�i��p���<G3�C����`y�K }�E\Z!�3D�r²��EcE����n�EU�<4�Lǹ����A�t��s={�|R	-3�Wox�	�e淺������OK�a�Rf${��8[���ѝC�H��N�����=�� J��K��?��#�p�pj �t�X�Ē{����h8��<BuM~�a(7��;⾚L;,�������`o��޵1�[Fr�a����4��:��rJI>����� ��N �6��$�-C
g�齊���,��@����OH�1<i����
�!����1���#��~X�Ʀ��Zrx��h�#�ޗ
N���w�OZ��H5���X�Rю���
���X	��G��z�^Հ��:��:��0(���z����'z��R�]�zŞT��0گ:��kԁ& E0lY�q�L{+U��)Lt�u �8�!1�vZ�萟􂴐7�f'�9T��Z���ON4������=}o)
�?/��8Գ�vxLZ
�#�d(a�)C�y���!L��c�G8�>;ڸO�S����:��iW_J��dH����9SҌj�w��O�N#)6�d�� Ab�}F9�{�0	tk#ױڠ&h���Y��x��p�|���v��j�K��!�����ʙoE؅�����=� @�˕�X�u����Җ)���]j��;���wc�)��)�  -s\�����x��(��͘�l+�Q�T���3` .w�ō�w�~��gN�Ѿ�X�u�P���T�������<V�AN���W!_�UĲ�} ��ߗ�yn��%�C"�Smq�R�~�Tڣ���Aa!��{i������L��*Gd��=��UF�G>�7��,�EE�i+�=���#�,��Rj��P{���+���]R�s�8��ϧ���*1U�H��W��Q�Т���zB���5^D�s�2Yb��m �su��GGBFe����g������\�4�i@1}�V����x�i�G�N��h��T���1xv�$��$�,�_᢮Rת��Y���7�n�(�?l�<u�U�B����.�'��r^�W��?jFP��m�_~�O''� �g��΄�F��N���]G� Ӫ/$ ��b=X/Uk�U���1+t'�e��{c����	ݷU'	�)�w��@Z��J_�%�g�B��d�.�ih�g�������^#�;�$�/:��s/�t��oY^��>��;9�)*�ֶWEv�j���¯P^fy�`W*��ڧƵ�҃rW~�Rqį**n����A_*X��6w\�yi�8o��3P�8o��)������ua��C�+��0�	A������~���ߟ���ޘ�msr�������h���G��[Fw�n)#<��?�=��wy&�}��Z#)����ߪ�^�o�,��7K��3�:~D�6�����?}.�W�آ&K�wƞq�$K��2j�҉�
sߝ**Q���!F�B��!g�W��x�2������BG�0@�ۄ#ʏd��d�����oEzAІz�QR���a
Z@��C�J^�{���6m?���l�n�ى\B�-� �אJw#TC[����&�O��>p4%5�e#�E9`�*Zjܤ�M{m#�l��Ƹ��WdQ?�����v7=՝` @����(�ߒ�R>�\Xd��2<��sӽ�O՚|w�U������v!H����A�O��|�X�K��ނ}�;A�BG�����=|ܵHo/���&
���G��1���|��p��.&)�O�/F:p:���=��ak�
�Y����3C��o�n����ek2�]�@��
�Ok{&�l�=����x��Ȓ�1��;*h@T��[-:)h�i^{X��K��)BL�q��� 㲻������F �|	�pM�Ԙ�K�2?������d�#	�V�I	�7���������%�i� �e��t`��+,��b�)�����e7��ne"ZIb�}��#��k��X�� ��x��EFO�ĩ�
���e"����c�Q�IiČ)O��a��bD?�ax�J�:s�F��>�άN��m�	�!6��,d�GA�x�1�?�lA����`b>������OlK��s�a������xF�A1��@Az|��ĥ/C�?�N�|��
FW-.c���
�����0p �7��FlM����Ys�UW��t��!7�'�ޙ�Q(h���{�]����O$䑎�p�#U˴�٪���~��F36F�c��2�}�5���V��~����r�Y�MqJG9�R�����8��L��s��