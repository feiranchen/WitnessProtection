��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX�K��w{�E<�h���沣 �B�yP�?L�j6k�؍$�G�Q���<y�s�q7�Χ���A�@�7+2�B�8:���H�DS�^� ���7E�3���.(��I&�b������ɚH�������eq�;=�8���4���*�����0��x������/^�d^��+�~a��I�c��[ۍM��ƶ2�>C����G~y�A\���iuO裑�b5�|�sŉ8�kb0:�����eFTb�g�jT����Ԑ[cP��pZQ�T�@���G�;�y���W�!���"n,�����ޚ������h�%�aux"�Ƕ�H�v8�A�30��gH
6�A�ilh"'�b���,��B�U��S����P���mX��2�e�,���j[?5��W*E����TP��>�FUY��\�9tR�ME.�9�HvE���c��SC�g�p�D��]�ﺹ��ᅎٟ@l�L�}�����]RM��ใ��������]f��� �}���tҋ'	I��NhEk��6�&aߡ#�d��G,y�l��IVz�?��0�o
��07�s�D���p���s��6�_�#�ƈ�c�=t�>��9�B�v.��P�p`=�ԲT��ԃU����]�5����"f7�n�!VU64���H��[�� Gp���B���v�~�
|{��u u�}�D�z�Do�!��������=�� i�I��"�VÍ�v?��|�u����J��!�^����鯐�Xn �Nٔo�/9L\�pWD6^���m^"z�����yc�N����ZZ����+cB3dௗCK�
N���@�U~E�t6+�!�.0�����?�9�F���c�5*�GQ�iC-��&�022E��Iqx>�w9k��n��42�=,��n���+���t��)��U0���T���O�v���*hT���ˋ����ֽ�	�E�}����QO/����dzjD��5	1�`aNyG-߰{�9*�o�6AJ GF�կ
���Gq������K����.Vv��6]���J��@���n=�lͶ�Q��ذ%u *�k��9��JrI�F�t��٩���4s�+@�@���o�b��/����C��u��(Jb�.�����=��n�M4�!���IYu�]�S�{t��(`���,�"�����LAeu9�9��ƚ���q���W� ���s�I� 
"U��Ü����[���4	�+�p�d�v.��h`�*2��X
(����9w{Z�7/���Q������oJm�&�<s��ف��W�����<��mB��vcY �l8�>/��o�+�ǅ�}s�Uh����J���� W���~���Y�w�x ����e`BE<<o�o
a��Ư>U��	��l(0���|�zGU�}6r��8[�u{
~g(�4�A��qO�(܁R=?���庝ۛ׹���r���w���K��Q�?˗��C}-�1�������qb}O 1�a.�m��h��M~R ��#����;��a�$ҡ��xO"
[%��kId;��
 C�w*�:>�*VHp��QX��p��-��I�qX�`�jq�p��dJ��=�5�&�	ET&ܫ��%	�%&aS�v�-�$S��!��ilRt����B��E<T-����v�k:�ϒc�&�7�7a�4�Ԋx���e +X%3�h*r,*� &%�K˛hr4��3�a�;񉛒'<�@���n��ࢨ�#��h�G�+qH�{�A09�������a=�9�Hzf�S�����}�zW��t#v��5x:&�q��P(-�ц�9�����Gj'�X�@�;�0�����@����l�3����������.�9E��C2ZS��
7�x_l�F�\��E����X��䃀�ݣ��x�ZD���-��O�1#�����B��q�r
�BN�7rx�g-�,J5vmyY���IW5�t�,��|�J��[�<�A0����|$����F*�>c���9�CF8����L ���" ����>�YZ��׆�p8��0Ꚇ����[���$6��m����؎3dوYrમ�}"R1dl�{�?����r�<<F�>�/>��f��׽d /�9�7<aH��|�)nʲk�k��a���>	T��p�}�]�L���YSx)kU.�"���̯.*�<Qº�Q��㺢G���s1���`_P>�G��r�e�^.��fe�.άg�j���;��}cY>Y�*���,�n-��� 
���N���"�؃�'��f��<�X�����~(�K�.(UQlK���Y[*3�������x_�e)���(ՉI�[��x2�]�I��b-��,'��0/��Q��S(L4P���SH����/D#Zr���v+"�j2�p�ߔG�X���4�z*S�����4�$Ǡ}���iqs=r|{�>;��<�eR@����?�QwinxP�:��_��T��"���������%�p�����1_`H��ʭ`i1Q�FVc���wT�3?ɾ��t�1uY��Zd�F,U�6ߪ�����P@�܆�������)�ݔ�d�f������n��X�T��B�K�ͯ���~a�[`���>byMT�K*�q�D,���g$���׽�ɪ�߳��6�6�\���0>֫�s[&^����Õ&u��w.�n���6�Ơrx,��wA]�U� �?�yֽ���U#Y���.�*P���MT���U���s&5:o����-�s������iy��*�ۀ�Sk뎑Z��*4�#��җ�^/VT8��*���	��&�۲-xQ1��/h��i�|>����bMe����3>ǭG6�Fp����=^���a&)��y�SX{�$��Gu�]Q ���S�Ѥ���J��
�q���et�O~�t$w[ѥ��O�l�V�T���jsf����-S� ��g�n�L���B�
!^A��"��IFg[^^�P�:Տ�Y0�p�+]Z(�ӯ�����Jko�ko=�k��CE�!�� Oo.C�#���p3:�]���pK�Z7"O��P�I5n��h���K��>Y8b6�=O��3���բ��K�J]�5d� �z�U�	�Y���kytL�>b	�q������f�)���B�J�z9�Qd�Y f�t�$�z!A۶�f:Mt�Ԥ��pȸ�:Uy����w�84��;jК�*�V��W��K��>Y�+��<Y����u��.�/�m�O��I̠�_���3r���]y��Ř>I�vcȘ}�yv�-C���ӏ6߽Hs��f�Ѵ�r�NGB~��v���T�����<�v5�~[��ܬ�R��۽�������FIs��]�� >��q9��i���]<[7��o@���㼉��F?u�6Q}00�E�]M7���
����G�~�׽�;X\;�R�Qb��p� ㈃j�j�<ӣп!�D�� ��;���y�>����PP�A=�gjb��oK��3���}��g@����+IFEńu��.��e���4:y4����n�x�^z���z��10�Sʙ_�Q��-*�ƻ�v�����J����f/��A����{g	-Sߌ"�����t5H�����$w��~�0<Y{*=�r/5��n�hkq�)�a �<dδf�����b 	9����[G�I�u3+�̕T8Z��^k����$SV`*��5u��S؛އ	�+��l�ա���j?�E`��\m���m�\�$x����wG�B�z�ݰ��E��\������t��
0v�569��j�n��gѡ�F��;D{�\���׎_���G�r�Eӿ��X<Ҋ�n���"ha��2c9�Ʃg�ԑ�ٕP����N�R���+A����<A:�54���(��6
[\�S���2W�h���7���&���؀ݑ��"Vp�#z�1��l03M(&�2�k����l�`��tM�����lf�!�bpST$�,J�����zB�X��-�ǯ��kϠ� �$3�7������`u�H ���&/a�ǝ�;�j����ٯ[1my��.V6n1bb����R�f|
{밋�.����!cC���%\_�1CҸ�[R�;��������tK�?�]WFH������ڋd�S�h�e<�d�+7���cU7��f���<����S�l[Au	]��A�oc?�|����?y�99�&0�����/7���.�'C��Y��ݣIMoE D���ўc�K��ThDc+�"�v]���K���B�y�Ohb��vL�Gs��	�l�T�,�^ɈY��<�OYjF�%��f�@_�+�}@O[ޮ���qey�a�� �$W��Ay!�w�}��,�Oq7&�OG��}AK�%Ն.I=�yZ���3)/y\j����Go���I<o������s��J`ܬ'��U*tol$�a��=���1|9!FW��(��q�r_��y�wB�E�����+%ï�D*�㶳�_�H3����[JT�����y5���Pp��*䭠��',�Sv��K��J�Ų#$(6�+Ԡ^DֳX������1�u�`�$��Y9��/��X�7t���Q�L���w2�������E\rY��\oW�xx�H�Hʒ�rr\�>�^�j&�x{#��|E����jy�k�P|8�	�G j�q���Z���?0=[���۬l���)E�xf~&�и�T����d�20��;*L��eA��y+�P�j�b�vܴ� j>�%�/���ܞ��WB<�����f�A���-f!�&S���ǡ>�HPD�`-Е2���Hw�$�$?r�|�r,@e���V�Ù�e&~��H�������!��@��y���X��G~��j��]4i�j��da3p�3����B�ܑ/����Ƈ���e!K"yFn�&.�o��(
f�olސ*C|���UR �9���N< �}(w�H8S�Sǵ%Ae�O��:]Z"�<
�z^	x���`2VK^G�j�Hn�����sUʧ�s�QwT�n���Z���[a[� ţ�U9�1}�O���Oã�Y*�6R�{&����g��w�p�R�VE2�V d���+�b�����GQ�Y�N*�d��pB�2y��(ZY� ��S'�P�1�۶ę-�[�KՕ@����(��Tw���B���w��@P�I��$j*vw��ڨ���n�"����h���Q��[��$�H�od�$�D��%�K�
ȡ���,�6W��?:�� �`�Jmn��:�� 7ҙ��3vc�P��h�dY:_;�X��YI&���*N��J��ԼRX��XGRF�@�������v�e��)Y��=0Tx"�#_�����>HÔ�9��]���/�wI_�.=�jAlPO�ĥ�pC�F�wՉ�í�6�8�!�*V���b�a�{���&�ӵ�|FX��CՖ���O�N\>�"��۽޿%�U��=����nc�<�ޣ�jLH������s"���]�|�B�~�"w���_��I��x�N}��t:bd����0ؐ5	�V���I��z��!��a���'���c���,e3%D>�L����0U�}���>�"���:HАK��.rOQ��*'�X����BM{�N�.�'�n��P���<տ	�`�~lM/��p]!=�����:�W�ȥyhLP)OqЭAj��
���]�Z�K&u�T�U8,"�����Я�>�������{����眄�� ��so��fI���j y���2��8cAÓ5�2�u����,�Y���w�^�r��֯Q�S6T�*B2ls��\L��J ����&�|Pq���`����M���o��5Sj1x�9;k�����T� �a����-t�.��άϵ���$y��\C3�z5 �4��Q4 ��1��s�O迖
v�R`;	���N�(/m�+�#e�(�$�AS&��9z�D�XC� �י\��X��vz�l�T� 7?x>qL���K��)�tϳ�N�`�!� +��A��E.כ�1�d�"�H%���*�]^M��kdQ�w�܌��4��&�:�/8���@࡞� �r��>o�O��{e6��Ge�bd�#�
�j�+���;q�ш@��ܕ]a��jL`�\� �懸����1h<�C?��v��F��iGҍ^�q��6	Q2�aY��g֤�=�&)m"��E��?�7Ǆ$�3R%����V��9q~�p��Ğ�#���+d� �1�C���\�c�L�a�\-Hӡ�8���
aRvb��Pr��F�o��8.2&z'(�`���Ykp��{�=@1��R����L�tو6��r�r[4��CY�9��mJ���9y���\
�ł��Q$BC~��ۦ�5�Yy9(ѕ� ��ï�9�d|���m`	���a������7��l ���3���tEaU���]n#��_��j"�e�c�03.ʠ,�|Aa�3��%9���i�`�@B�yL<_��s� __�$�Ƒ�3m�a?b�G �բ��&������0:ņ%m��^��&���p1�^� �	����D��hبH]��I��>��q� ��JQ�����5����H�M�Y��7���)��O����#~ܿx���S>�J� �,�\r���������6�2pC\
sdd c�p�R�F���>�EpJ�`mh��@�X��ִrc|`]N�ן�0[����֢�&�������2�_l:��f�haɵ��t��	����ܢ���VzA�7}S�Mx$g�ͧ����:��d�U#�vp�L��f�s�����+���P�� º`s�G�9n���e���W3;��!c�	sU����	�u
�A�Ѽav{�����ߖ�J���}b��|Y$�A�e��Pa��Z�@W�^7L�M�A��2e��}m�VO2��C�;e � �7�o�k�K<���ޔ)`�0�^��`�_��rP�tQ��P3~^�C������0����W�k���f&`��>�/��msQ�}J�'�n9*�Mj${g�93bam��a9�]����鵙W�3�H�m�۔�1N�d��n�c�ĺ�1U���zI��N�UR��v��8��xtAބ�L�z�X�>��	)6��-ځ��mS��`=���%F��١��.�Ñy�L���'�c���wN3\BX<C�N��<�mB\U�e��d`��T�R[N<�]g�u�oM/ǘ�a]SO��ί��Z��+k�؜����q޷�6�ؒ&��o���0\��g9֧'�*Y/3��?��cv�ъ�������!m<h$���`~���ߚ�H��Do;��W;�R�\t?��ģ��fz[C��X�\ܢvM�gxЃ�o=be�	�	)�͋�4����H$�<ɾ�z�YK��=�wp�J����ѭ��os���M���>m�H T��h��"��=Bm�d�
�*r��H�	7�v��Ub�Q�f~Rx��ܩ� YQ2"���b�������L����p4'f��!�{k�� gD��?$�:���CS����1|��_��.(�7�¾�a�0̺��Me{��š�/.��-���լg�b��֛�d�Gm]���e|��i���bC���CK�Dz�sS�R C�c�Z�t
Ƽ������E�Ń�1T�g։�V�>�m�\?pҔ�XDQԘq�g���/����]��2��5�X��L�6?0.u]�0�#e�d3JʬAm��i����k�-��\���S�U�P<�ɒ]#yq�,���@�E��{�$���pG���,Պ(!�^Gi�͹3�64����X/?�nW��B��K��S�F�#!-D��~`�͊��H��.H�A����upHS�ߒ�w�Ѿ�ւI�q�~��7-� y��S�]A�a�D�� .��.>Ϣ"tU͒%| ���%�ƕ����ҋ�� �7�+8�h.���6�,��VL���v%8q�)��P�a�˅�j`v�3�ɖ��o2�=�z(�"ŅC%I�(�{e��y�!G�1�p��=\D���J�r��ϻpf���$#��}.�wt���%;b�|{j�)���;��蜌;k���[���Z�=@��f���YQ���6�[.-���W�.��w�CN��r՚}u����q(+��k�Ba�_�Y�W';�Q.��dC�7�6룷������  ة�J�
ӎ|��c�b>�0�kL�U�s̖4`�Ug�\�ʸ���j1�Y�
��+9�th�x��G�Ll�ram)��De4��$Q�#�'�r���q0�~:c��lP���2n��v�h�1��Q���,�}'��`�!����W��j��7��(�<W�`�\RJX���[�%�}�̽��3�����#]�{`�aU����C^e�^p����莇�N�*e<���V0o��v�|���/����T/v�F�� �e�<�^}Q5����'f=��ak��Ãyn��� �c΄j��V�/5�|)FY���.�:���0G�x7с?��g�
��|`#�؏��t	�üL��E��j+����z;[���� A�3N<10�D���h;c��Ǜr'�ź)��'�룫	{�v�}W)^��1󞛄Z.�W0��f����� ��6��d-|��:�⟃�~�� _�A_?w7?�r^DoyXl�v�c��sS;m/���D�!�NSF�_��a������A�˰Pѕ\ГJs���W�hy��^y����<|�f�|���T�F�U:
`��.d�4��c6t>��F*`��6���6*$��W�X���סa��o9���[>G���m�h�'��M"�=�A�>F�Y�I0����`KT�X.�[�rk.ę�&�T�	��Q�hf�):E�x���2$���^�A�u�.���� D��;Eٌ?��,Kmc�_�H��07 Tn���2� [�D�]xc������~Lk�#�[��I 4���r�5�V�0�8��K�������(bqf�s�ʯ��,[+�:�9|,Z`�}:�IƟ=� 82��4r٧��ˎ���=�ʹY���!̾H�ٷ�as[��}����|e�����W��YӉ�~�����)=DSU����KpA��p�z�jV9�Ta=��[i47�i��Xj�_�U��� ���)f0X�ri��ѦU����
��S����gɐW���9fM���wҜ����H_��o������}�|�@���1� і�B#��Y-��}6g������,�9`/)��Ǩ�k��5W ��q�ʯ�K�2��zꡏ�G���5�:�Ѥ!��\Z�xm{=D�X��⁹BԼ���n��coW�Q��	u�at3����=z���Q"�y<�Ư=�����&~:�?dɛ��GQ}����&u�T+�o�~X3�w��-~V>�� 73��#�!,��U�^9o����rcҿ�kvG3,S�i��};��s�4�J62g�Ly>>����i.2�0V�A��0
É� ���!�.�dYO�;��=(��������P�����f�S���C{�h#�Ws_��_X����7ʼ�op��Xb���t��ȋ7�\ZP��d[!Kc��qu���WJM/�L��DܭUg����<n��2�:f!�)1��-B��E�~(:�D�0��$o��6�.��-0��Ep���t~"�M�t jX����[w���,̬�J��$���lxV��A)��c�_��Z��mtT=���]�5Mf2�n:���� ��4:A���\be"0��/���6��9��W���*.{����(&�q�ѝ�z����<M�_i�ӹm��P@���vW3*�{A�l�Q%1�V�m�(=��r���$���bEhCB�D��K�[!*�Wrt�>��1���Dd;��X�[������\d!���.P�0�xX�9�N	NUPx��s`0*��	[�kb;]J��〉��"S�tIڵ�o�ݠ#|�#�3T�t�֍��Rlm3���Q9Mb=����t��"��_Ͽ�x�.���
77V���e(��ƗW�a�/���)�/_)ut�#CĹU��1V����g����p֜�]|#���X"z�^ȕ���U�9ɭ���KS9y���9���JYv�u��'���J�;^|υ"�$���z��cvs҉},d�F��V�������Wd6��R Cj.�l�/���g�$_�Y_#���(��p걅ݎ��!z¼�k�Ɂ>S���ɔB��SmKx67��}p�Q����sl�ǲ�z+v�9� ��WL���R���('I���d.]_G�޲��\|�#���%[w�۠��4��J>��ƍx����]E7~K����5������d���]�X�{^&�얎v�x�<��W��l��喼�e�����~�_�t�4A �<@_,��?�����9�p7��&"|�\�<  ��ԕ�Or�T� �����Öe����o��ǚc���=�]ë@&=��j�੄��������9�^f�ڼ��vr�Z>Q��l��*��$�o^p���I?���p��H�q<Z��H E2�Z�o�iJ���Y}lk���$Ђ>��h�9%,_�%�~6`�~ZKH�-�,p���L�A���:�[`�u,�� �;��gבh�uI�k{?�����o]���; B����#*_p�-@'��V�iCT�"2'�=R ���|��˒�=o�:�w�Њ@h+0J����!�ilm��ii}��y�*�\��A%��K.���4[�^&��Q�eEho���1��y�(#��~�y!^����JFx"��"�3�Ʋ�rMo7mo[�{��S/�o���!Zًo��^gMT�=�p��yU�Gϔ�a��G�&���:��,�Lij����,4���"�u,�T�� �����lx�
�|�u,Cݵ9��0GU3W�$=s�������!�D-h�܊o�մN�v�Xy��w{w�,x�HX!����<��IJ��Q{�S�7]$&�L^��Wn�$?��ܫoH�l�y��Z����A�d�^6�_j�����>l�z�