��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f�\�G~m�7>�#'r:LS�^���{m���#�kE!q�e\�A/r:�e��.�I�td�*�Ć��@*j���	]13��%��[�L�����p�n
2!ӋOV�dM��)��������t7����^����B�H�FD��U��!�<��N��	NW;�K��G'n0��e;�N঺�4�3����b�qu����&Lh=�I!�W���z��P��o�}4�Vq���\�K�l{{_ ��؏d?o����^U��;�".�jH�g�Bq���ǒ>��S&�i[�v�������ؤ�r���dܿ0+w�)�� Gfg�C��G��� ��m���]Q8f�1pnXo�&ǖh|VcMBv�.��ef���Q�i�y^�-�?D�����]F�s�#ry���c� ��>��o}����̡��[��p6&��#�zLZ�d�-�}��dCn�-m6
ɂ�øx`<u�>ʹ��z�8@;F��. �+a��t~�V '8�_r�9y�^���m�,!r;���g��;Le��tQ����G�*��X!���G�@�Z�sM}l��b.L�&y��I�V�7����9a�FoJ��P����A����,�yCLFv�H��c�\�������\Xؾ�:r�Zn
�˥m�����f	>e 2���2�h`e-��%�]^����GEf�KF�6��jkr�A�|�x����p����d\d%����n��c�*��=QZNRA=���9�dc�b|��a;�T���]T���S�6��U�LI�؀~�6�V�$rx��FBӼ2R`!j��	�ˠ(p��O�a����x^��a�&�O���֠��x�O�@�1��T��Q?�K{Y�j�[m �.#r��*���yO��k�B�8�k�?�pRM���c�p6�V3�U�͗��ts��ĝtWB
o�� �`Kcu0����t�W����Sp�_��L�>�v�$aؓ�L�R��֢���$���ө�Ϛ^�v=���W�3�.�8a��2( �j�2e��q �n�@p���:�^��"�2����z�?>�B�^�p'�)�0��bu�q>A2�L]���6��	�����y<<@��Y����˨zF�&��|@ɻh%A�@����F����h��j-���'-3�L7�7�*�^�E����šA���+E/�fb��/�5��S��h�b�~*���/9H
/G��YA��@>S[���P��'
����aC	S$��*�Ήe!�*-H��~x�&��I��͚П��H�b-ָ�������@JӭU��
��j��יZ"�V��ԟ&�ܓa}'.�ך��@���f)Z1�b
�%�M\|��_��R���l㾙�:cMS��%o�<��)�������ex�s�*x��,�</�H��W��v��:RP:v��B�����+X�[1�t�h���kp��]�������j�bP���oG3�j;�0�'/���n(+�X�]�s���'�N��=���Zٜx�
~��$֓2M�`��%-�h`��TX���u�O��"�`��*�i`*y+�����˸�##���Mk[�m4ݨg�ʭ�* ]�U �_�������a���O��σx��n�^���W�ݶ4�����B0X���ʡ�D�]�� hݘ[��a��V'Dvhs�4i����y��fH%�ŅH�Jk/#\.X�3����Û��({�z�a�J{;h�P��Zs>�4[K/�9B��q�'�u���h�Q�ԛuJls�J���d8���m�L�c�O�4n&FMV�{��������_��q$�	V�B�^`\�{��kF��;ì\�QM����[�,?�/D�ݏ !ؤ���A1{���`��U��O��*n��/%-��j+;z�+Ng��Ms:l��������#��喂`�h��IF��0��82E�Ręנ�C$0M&�3��9���z>���׌� ��{�1��OF���,D�+��*���g0믆/�R'�Dw����(�������s.7S`&�V�?:6쬝� ��?n^����c�BE�s02���$熂��*k�Ž�&Ji��1�B�C� 4�!�|P<��Ul�8Ȑ߹��p0N�ٔbY�Ӣ��r;ıy�BQ��;�Sᘬ�?	�u�
��h���]��"�_��v[B0_��COK@`��W����n�t�_{��ӣTl=�H����U��\V�hh�ק��;i�Oo�B�+Q�7��v��������ϣs;�x�
����Vy�!��]P��g���W�=�S��H�K���l�J�,�䗖Ԗ���Y��dd����|tf��K�A�0 �?3��~�� 3��f톲u��Z�:��W��g��7�p�.f��F}�S#53ٖy4�(o�c��4\��Բ��]�y��a�Y�(�U���x��wl@gĸ~�z�5<���3pgO#�V{�a��s�Y������2L�,�����V�e�N4]<R��D�֤&,2!�J��T��pO��ը�O��c&�[�vkh�ja�2�YJ�zD(�-QϠ�GL~1�n��~Y&F�"�]�d}�C!�J6);�
HvZ��_;Aq�1\q���;�����U��*Z|���A2(�)H(A]�1F!��w�\۝.���f�T���I���a��$�8ޞ��|�F��o9������7�eh��*�rΧt�e�#�=�NM� >}á��wKd@��x�Y�T�E1GI;/�'��1 ���{'�-c����9-�Y�tVe�����*DK�f���G@����UB� ���~�. ~s��敏b0�7׻�~�c�X	7�	%Vn+�#��X;���R/�;��]�v�\�Z���L.���ԓ.�n�����B{
���yըnu�x����|�z�2
Y��H��T��q��� >�a	��Ξ�*�*��WH��e�B�D�z��w��`�~PJ_��S=f�v��*yn`�����pƸ�qkԏKu3;�?���P���&f̏n& }h��]y'?v^_��)k��qn�������6�։O�1?q�c"�ș�D%�����|~"sz�j
*��н<t��Z��S9�P���A��}��8��:�f��*�e�ǀ������[{+��/:$ ��i���7�5�p *�6mڂk�����NI�!*�Eu�ԷC���;�"�qk:�#
Z~$k���S�̬:�ڻq��;���${�p�#��VU��5���.Kb�c����oE�2��$�c�f�Na�N��d#��gZ��M)��p��*�]�/��l�1�z�!��z+(/e�T\�������쩷t�v�d.���T-���qQ�I�\��x�¦�d>��mEM����.��6n4�j�`��u���ޭ?�ń_,>��ilt����έv��u+[۰wZ�2�oKC�q�F��{��e�Vv�R"�,�4�9H	=Y�W.2�pf��|�=�8C��
HZ�?��L$+��k�-���aGJF�m��l!R�3�n��Uo�'�|�Jb6���V'�j#'���`�S�"��ٷ��Cѣ!��4(�j��\Ŗwo��*���AH�MHM�����3K�b��(Sv-�1"缨ep����h����y��%� -�&G\+,.
6f���_T��>r�&�+g7
{"��c/@D���j��eX�P�@��j}H p�~���?�ʫ`��A�s�;3;{�4K�����ru5ɾ�e}*ƾ�',)�z���3V�i�(K�������:At�����A��BQ����A�����\��KUyA�D�:�[�����>eV�,�� ��k�.���E$72�)�hLOh��X�,��JLqL7np��ڙk��yꗚ� �:/���P�$k3�A�NoSJ����7���U��
��r�]xh� �- sA�5�2S��"�� ?�������u�ɑD�� r� +w�fIf������6����g�l�NAWۥ!fNA�4�ѽ�W�4�{!+�"���$�[��8��#���\�S�ܲ�Ҏ�Kxd��2�*���q�Պff�E*L�mM6�	Tks�i&̪E��p�?ݸ�X��{ĺŹ������1)����=i��b�
 ���	��� ��|$�m����鄊R�^@��E��I�n۔���FM���̌b��;�2TL	���´��4�D�J8�2U��)�4ێW���擠����,��3��s\��%�X33��&N�#Fw͐�"Vt�=���i�������:�7��/0 :��1!���L8��)�q�aR����h=�.'N����j��Z�W!�*���m����5�&H��cgl�!�e��C+���_.@���ǥ��v.y�J���!?9lw\Z�3��0U9�>.Xlfʦ�����}A�����#<Y��%��2���Վ�02���(��g��<�	�i���b��BY 
z�n�������g�	@�ʱo�v�v);�"��K��F ȸ��߇S�������nM{��0�K���是�����zL�L�qs�!!�$�smHj��)�v�'���n��3RoH/!Zf%b5 ~cy;,U>���D̋��@�ׇ֝Z�y�*�t J����L�5�䧄j��y����������c����߀�z]�)�k�NKg���	���������b���^1����V����Ћʯx`w\�g��c���N��[�$p�3�*?k����-��;�z�[{�j��?���d؏�&1�E��`&�s|!N�⪎���8��^(;]�+ G�ti�[�����I���#\�`�m���A%�� ^dR�Kp����w�G�a�!ɖ�A�ʻ�L0r�W���7�n$��~��'�e�y���δ��g�s��s}��Z�����=�s�t�g��л٠���Pw�L�t�ǝ�yD�m�[� ��o �j=�<�I���^��B�i���GJ).y�ڝ�)r�8��bX��R�[jY䱚��P�T�7�-��n��yV�S/��a�A�F0��@��*͒��d����f������.��#}Q�@s�^�I���zF藄լ�A��\p�B�F>�Ւ�29��Ȳ�=q��j�+.�ᵽ��^1��3����V-��h�B�TlQ ȭ�!81�	��DOS�-H��W:�@{H�!wR�2�o7�<�S�nO���R����U5FCIZ%=��;n�;���2��6VK^�PŏGE�\���R��X���o]�3��@�ރ:�5n�e�[m"�].夵1�i��Kt�����b�Q��9E#g��pW���;���j�$>�Tx���x_�)�]%0�S���%Q�U5�q��0abkj��Nԉ{�`�O������qFk�a$Zh:pVz���4:�UU]�IK5���;��r6�p1����L	���2�?;�ǫ)��K�h�#&��$3���*�o*}?>�� %���1��#h�F��<�.�	}���sv�ʹO䤄�G;�`����~hp���V��]�r�_NlW]�ra�9'"h=%��4 �hCHQ�ZH���y����h!a���3�{�ν~|k\~���1�:}k�װ�����7ǽ4<�%�ˡp�ḃ����n�Zlb�IuO�apu<+:J����'
�7[�0m�Da8?z�����	a<�m����:=Ŏ�HaHbi �%��U�9��L&����S��i`�[�5.xx;��(����.���.R�%a��}�p{]#��X��Q�_�W�%&T��	�V۝��_������]�<*Ѡ~5�3v��JN)��%үugi�����d(��Hl�f#C]�����)��t%'�N�[�����U	�����öthj�ӗ*h� )�rO�����������-�y����#���^�}��׏TQ��H�+L�c	"��cf�۬�+���H�n�+ �����qn}�9T,��;ʊ����ƌ��O(�!�͵M�l�JIj�sO�E�򫓌/o�OD��qDT_<��$#[��hbr�yV�q����Ͷ1��������S�d2���U�$W�4�?�yG`V�e��E�kn�5���!�����b2�Y^���z2>����+��I�@�F���'��t���a��烴��S跂�X��x�_G#�@���ў#�BV)FR �aq`���>�E��'�w�o�*�C� Dg����z��e��w~͜�8��+�%S��>NTo�����s�5]Ӛ�����?�Kq�z�;��(�O.��$!�D�c��#�3LZ9�əA���MW-�+;��*�Zm�c�'�|�D��9���(���*|�������-���U��o��[h��jڰP$]�~C����B�w�R�T���MaUˤ�$`�{�G� 2��nSQ�O�Y;�5���:����2���v}���^�XW�?�Oi��X1�x�������:"���A�~N;��0�W9�_==�(I^� �5y�NſVA�?-�������gջ!#^���)<7	�~F��ƻ�C��ib�ן�$�����@j�|춠|�m�q�����GAOy4�N�������*��@YM�cyx�^����ӦtA�W�[K��i�t�m�&��_�����Ӆ4��=9�3�5`�0���C�4���No
�\^I,��}��3v�]b���!S["��k�2�S�Z��w��G_Ml���hH�9�A|�8�*|�|-�<�����\�U�*ρ6N&G6a9N	)o�qz"�/1c�VNi��<q��S���I�Z��`thk�n�O�@�뭮iӼ�ɢ��.ٶzh|�E�E�F��A�є9�!��T����R��h��k�����3%��ŧ�F��E!r�L���>��#{��PIy6X �a�4���$A�������4	Z��m� �����7�
��7�̽��]O��X�P�&oCF\��qFl�'�lH3� ;�<)��\5
����/�FDvYC��\������ce����:����wB�zg_��a��a�/�tQF ��a�B�2���F�@JI�n�ŊH�X��W(7�����ԡ�P�y���G��k~G�v�3�?���7^#����#�*«��dY0o!���,A�r��� �~d��*�d�5MOݏdT���T���M3��p/��h���N8-��9�VD�-��_�P�)&�|����[���ζ�5�N���_޷�/�)�#�jY�i���V>߃�מ#�sL:�^��W�wm�c_F2��\5��.����=䶭,�(%�v�*7M��#7f��G�����8���A]U�����9l������M�	Q�	`��r��<�Th �i�OA�.8'����a|sj�ꐩ��,��F���P���ѱ?I��ʚ�!����!������b�Q�v�Oq�.��K,'�L����;�'�t��u�!����ǉ�`�I�_��G���k���C�#d%Z�ȝ�*�|���^jvk�{ ��g�PY����+��Zrqe�!�����<{(��:$J��['W�xh�~�X��S� ��� ��qu�F���Fg�dR��	*��I�[����g���w���?��1d��C��,�`]I��>1�h}���B!51���
��r�O��]�ͻoAi���Zs~.̡�\��<�W�E�ه/-3�_Z���f/3�U�75YM�E6UX�����B󷘃5��EXy}dzj��y��A�y�v\�v¬D5i�G�o+C�_��x [��O�^������BS����Zb���)2^�//��lV/:[u��k�m����c��͗ydǧIWQߖ��^�n�E��-�fC;�u*�|V���.��}$�y�3����Z�0i\@��x��D����rS�"�L���^�w�s=�������:'�\�6�vsbP�u�<=sؿL�=#�N�V�e^��w�5~z�ݜ��w�eښ�Q�M�QL��K�$ْ�aE�E�{�%�K:�(�����ma����W���+����?�L ��u�AW�3u\��%�f��F��E�@�qT-H1���-f���My���^zk3R�&܊<4�R�j����T�d��VP(�77\&�@�̖�h^{[����K��_Ǘ��2L� T�Zc$f>�f��P��(_�G����؛𪹑��y���1SC7�	�SO��"^Gë�k�1;�Sj��@���o2T����_<p�G+_�E��UXu�ʽ�Ls����.ǂ���+���������:��|%
�^v��O1�l�Uu�%�z�
�>�r.�L�V4&����.
�Լ��VW����n��Z����za���)���j����4uXa���p��v^����ay�;��g�k�\P�o<@)�F�{�����s����Nz&�;�U�����M�`��k���9����|us��qZ$<�t���VG��)���e�Ś�3^�O�4����7c��Z�q|.
7� �� �!
wu� �����3���rf9�2������㰶'mv�l5�`��&�Z����dz}�2)&xcJ�fXN���w��&u�Cq.���f1K\���ŤPqy��{dPU�]���S�0�{�Wj�T��:c[�ո�ML����T��q� �ˬ�"b���?��\��� ��-�u���?ۀ<�t�g��1�f�닽�FyN֚�ϘݷC�<dί��E2TV��M?#S��9"�]���A]G�\$>}�?�Ѻ��Wx� B�uj�����OM\~RM����5|���n��@бz��d�;�ŗ�<u��ā���	?z���&����5s9P��^S0t3��j��	&Ţ�3�G�R�Jr�D�.nrU��
$�o���9�L\�� �5*[B>c������8�V���@�n��nZ�n�.�C	8���9�-5k���O�\]-��3} �8�����mT��6�d*Y�����T�B}I�!�ry9;G�[�a�%HJ�p|�����{6�o�!�݈�H�L������asݱx]箦�P�M���e��cr������l�t�� ���Z=ʲ�	~Hr"�	r�>�d���~����y($��[	�yn <�H��aP*g�#��J����iH����q�I5�T�?��g�['���rZ2����a��g�Ͳמ~n�Ж���R��e�C�p77we��4;�pd ����˩n%{h/��/�9;q��e���w�s��p��., �Hez2c'��G�aϕ{�PkeN��
���-u䛋���38��5�u�!�xH�ۭ�"���H��o�����I�����\�w���(�����`�|�O3l�¡��42�x�8窘����JV]����WQ,����t��2�}��OJ4�rpx��w?�>���U��A<2�E��AF`ir!�4�'8�]�0�X�gkHf���-��{��M�E���)3��d��ky��k��^�d�@k���S��r�gj�C� �c�a��g�e�Y��ũo�a�@����{�G�. ���G^6n)�f��'Ux�g���APQ'�9��;�I֨�P������O�ݐ�1p8K�5 a���p%��h7K���1�`�y!���ߐ�ŏ���x�>ex������u��o3b��T��-P[�� �rs��8yzs��t
����!6V=v��)3�[N����zR�E�&�$=�#�/�k-~U-uuCl�!4����sRO��v7�(��l�.�0�\��^e=(�dѵ!J�	<!��U���/�(���-�Y#/���<�Ź:J��N�J�ٛ$���զo�V)1�M��8�S[#]V�����lc<�3�s��?���=�#�9� ��\X�M�	;i.�P�!�%���h�A��[�SH���-7	�ܭ�.6V�������味��c��M� 6Q"������E���lU�SU��	�:�Q�>Oޛq@s�3;R�܍J'}1wq�e����Љ����w�ՙ|�vYX?TZc譍xzQ�&����dɂ�(�ӟF�-6?}��@��v!l���$����V�5Ц�eU��<�#U���U)�ca5�*�P�������H�ކN�5�0%���C'��vh!Q����<[̂��֓_��LqE��ף8F�gGc���6�aΜ�|�lb�l�$��o�˃/��K~�G�&�x8�4��#�V�)Ϫ��_(k�K�8�i-�4T��1�j"ˑ�>����|��-�Oݖ�(��o�m�%��īW�ƚ���Џ$N�+�瘏$�q��J(���jp�^}�O����-v;�v߯+�Y���%	�[�H��!I����J/mP�/�<h3��lxMNC�#�wL�:�Zç�^My#^���F��ϊ�%����W��keZ��Lh���63�Q�ʖ�T���A���*E�1�G���:k����TǤQ�S�w.���X�^�Rn����J��G�Ź��YXP�W���X)Y����Y��+`����U�f_dO��ն'r��T��I*M��p�_^�	�yk���_�'�'�Cv߯�C�,љ��'坥��Bs���h9�U�o��Eli�x���
����K����0�g�p�٢K(�|u�ܑ��;��J1^��Dz��&�i���Q�7V���~�j�|X�"���ŝ��A���-O���eC]��8=�c��1� �Ou�/�����-�k�@���H�4Cb�u��� `!�7?"���P(�h`7۠K�xY���nW��Pƣ&Zl��!�%?��x2Z�;3��tQ�2K� ��̱���{�Rpi3h��/Z�ɉ��>���z*Z�� �N�b�k��p ����,@Fz���E(
�F��)؋��+�;fp�ڍǱ�|�8�ܛ@zݏvW0�m��M$('(RL����( CX�zw5�Uy���?���H�c���j���b$�r�6�B�
q�P2��F|�����p3+�� X�Sœ�Zϒ$8���	6�E��ܬ��MA�þ
�����(�h���5S~���YT�B���-��w�T����3+�'��5n�s@���}yT��7-a�w�DY�a��T�\	��5�AYə�������*���t���&W�]��ojI��|�z�T��# �t���*���n��1Qy�Nߣ><���\���2ܙHc[*��)�����1Cf���02��A�0���ϰ����`����A躪hӒ��հ{�g����WV�3�_a�~�F �aߖG�#��^�-mA*����� ��~u��t��j��Å8ŷ��T�M��p�:� r0����V��sK ��ۚ�Ύ�94$l�_C�X�g=�q�*�)u&���4u;��	�b�������j9<�2��;���z<ۄ��e9މi� �M�Ǝ��/b��T��F��s"���v(*�l�>a`-�"�őok[�]]�*��:�<|� ��:aue��܅�Lc�y`�Щ-9��ڗ��n���n�`Ū$A����3������螑>G1��k�Vd���<�zUz��ӟ�Q1O��K���D[�)1�vM�,+?Q�>w�G��m7@颦�� �Z�&�	d1���j�3| �?����y��-��������"���h�>�2rhao#���F:�/H)�.�CY_�@.��l����r�F+KӼ��[�x�ҦK�Q����4�Y��1rK�Wg�Ԍo��T�b��[�����a���*}kuR�M�C�Jl�����9�^�+&�۬��*2}n���>v��iʶ��O��V!GQx�NM���$�J�ˢ����Z�&���9�yY����o ���F�^�)��yb#keo���äj��cd�]���� �1Ոf��w4tXz��!$�
��i���ƴkwZ�a��@�� 	e΂n�b����,&�7�<�թ��LE��7�����*� ND��y�E����22	G���RD��v�K���uab��l]������/BL�-��5�ͥ�`��������at�Y˶l����D���)2��&my:�yi�����h�5� u����#$Sf/�"��)��~U�v��\5՘ٽP�q�w�a��R-��S�Pp-�_�-ς|i�]��A��)�:��z���O���5�K}�4��/����}5z@��MM���S�ӧ �������x�Z��0�p-r�%�v9Y��>J
�-Xg.���{��ĖO++��%j��?.X�b�R�)��ȵz���W�g*��gӍzp�x���?9�"�$�֮B��v�	0����_��aތ]��v���6������d5����нw�B���0oj��;�[}� �pv酆��y���;�10���i��|�§�	Px�1��&*�À�X�?Ex��h��'��i���,HJV=���	 �6��v�d.���p�ġS�1�t�,J&��Bu z2����G�Ɂ��� J�-F��*ss��C׆�s��>|���l:����488>�Ai�ذÔ^��3ET�6y�����Á`쮂���P��b%��r;�>�jT��H��2|�tJ�V1�ǃ�rY@Tn���vNۯ��:�RO'^���K�ʼ 0^��3��O+�M�o�/-{�{��p�R��,�W�{�a���p�9`����o@M�K���Vpq��3oU{P��W�V�����w��&j�9�����Dy�����l� �V��L��e�_\�(��;��]��]�r�G�۸���S��������Tι���e4��0�d���i�^�
�"D
]ˢ�:��U(]I,�d��[#U\����g��E��U�%���H�lq$w6�}�Js;Z�L���*,
��MS�s+6S�	'�j�� xv XWeo�5A��y��G����q�.�Ad_�編����AnXf��f7�Uw�4�ԟ%.�,b�ƕ�79�1X����k���.!(��,�����o���KH���������s�U��Li����n�+Ku�r�TkbC�.r|��:d	��0wA�Z�}�e�\֣�L����a�EM��5mIA���ژdG�E��u�$9Z�ǣvK��ٛ^1���<E?����j���[%*�|��UA���yF5mUA⁙�&�	���F2��a����d�R7�8�ȹwӅ��䘷��U�t�[�^9�Z��t�':wWx�V��Z�9S�h<v�ܜ㶪וf����*D��p�\"�>�f���3%8>�qd̄�lT?�z!A|���Ã
�h�����x])4v֛N/z=IO�# ��j�����	�N���=�;�%=8���
��5u�:b0��dV�_�4��	�E��B���ˈM�P�����!.�R?�)6��V����Yr&ݽ#�I��6A�JV_��|�(�(tG�(��iR(g�b��*��[� ��k\ό�|zm��~Tù�Zޯ׃��Y� Y�_g��:��Qe�t6qhn�s�Rl��y��$֙X�a�t�k�U;�Ͱ��A�Q�1� %��B�+���P`��8�뉉�����r� 5z�VP�S�q�M���K`z�TJ�7�y�HM�)���	*T\�#�2Q0��R�6���N�P�ڡ-�H6���y�����������T����ؓ�hAĊ�J|��k��3t���hWq�_�]
��t�k�``n�7P2�!XhJ�� m����|\�� ����g���S�9�a�yd�K�E�B�!��"��5�SmiF ����ҕ
�7t�,��K=7[���~�lk�@�Rp�R��_6���pz��ᄜ�F=hu�|�ל/�M�/ �E��lQ�0��z�ϡ�j:Q���y���#�N&�D�aM��S뷎>�*��=�d���ԯm�\z�*��-��2��t��)/�N8��\��{ �y�ô{�%,i���w���-��,b�Fs����zc�������X��=�.�(�����K�����/ͻ�KF��BƳ\@]Rl��7Q7�>ѵL�VO,_��E�!��^&X��˷�c���$m�؋M�f�kA��!�\�h!��;�rz9]fj�߫F�ʠ�i�#u\'dD2���TrгC3�f��j�&�n:)� (�4��EQu՛���.Ա��>W?afE1/�KǦ���#�
Ë�!�/��KG�$�� }u�#үy+�[�w]�Db� ���G��(q͐E������%�R�t�y��`A�QlDq�X���W����"{��78x��8�*����� @Ϣ�D�ő"W�YaS^��]�$f�u�]����v�?�īN��s����O|�C���[�^ʝ7���W���b�c�e����XU��IC<�e��"ޘ�?�l�y�X�4jc�K�H-�~�0ʮP�ii��A�y�N�Д�� J�Hu����v�RHJ���%L�9��D>����T�+{oGqF9�K�%���Ux�k�ҴheʍxJ��zv��Q1��\�B+)�7g��L�����&��@rAT�^��`Z�$N0�Y�.�G+�juh9�^�^j�u��g�
L?Z؇�2y�}��k��-u��P%I��/h,ځ}��B�"�XP7�;^0���P��	�8-��ݱ�
6�ZP��ټl�������!����Ү������Yۧ1�:k:���� �&i[
���khbDMϒ��RFZ��.��x�֮Gf��E�{� *u��aK��Q��5_���7�t!�{�����h����2%�J0��s����$8N-"�ɩW��"*�A�)�JČ�!�0`��&>Ϡ:�}��0N��	�0��(
v���_s�z�f"�΀��O�3R��7�.���C��9+ڻ�T&�bWJ��r��*���ǵ���_�x	�N8����H[�x��Sܾ��Po��\�|h������T�V��(��q���0�+�"��iB$
<�{ʮyM�{�A�<S�e��+�̒wh��:#!�.�5;Z�b{�)����c�J��ӭrw��k�L�Mbb'	7��fvv �^�J��,����qČ�����Jo��@#�]�5@�6�|Z�Uǡt<�:���ra�┮t�V�8\.�9��z0·�O�+�ɿi#`O�a�O��K���$	���E��ֆ�����M��_=���-Z�[�`����9���mw	4$	��BF�$أިAp��j�4x"��-h���v�ޭ� m^����P����<�pgR���5�|T^�-
�(�{��i�!�Cg�P���������f�#����*oLx]��BUҲ�R�1:��oZ����X_�j���1����>%�����#�`鈛���~����/��a�X�y�~WoQ���dj[Va�|���|�| (5&`�Q���|2T�a�%h-0�mRц�!�➬y.���r�v���R�&q��&�(a�Ј�*��F��#���6Sc(�}��
:gn���a���+�{���tl#F�ѧ���� =�#'4��`����������i��W07򅴇P�>�M30�h
:�l��΁�/���`z��$++�#6A��_�%�ҁ-&'�#���ui��Ԗ1Ծx�>���>T��(�����qg� �t����u�,]	�#����f��ڧǏ[د,�bCNYP��CP� ����.��T�I�YX"̗��MQ��j؁��1߶�z�5�ur�x�H�-c����~�B������7�)nh/d՜��|��HhCf���b흦��T'�@�)�V����Hɯ�b�L:	�� 0)�W u�c{ܻ�r�W}r���17�����U��:{Ս���bi��{Yy���5�z�ǯ#��_�����ă�h	�q�%ǢR*���aӘ���Vg�dW�q	��n�σ��@o�| .�+���(g#pj��HZ��"��<� & &|0LV�R�~f'4Ūy�3�t��4��}נ����F�&{Ю�^h��L�L�Z�zebgL78����֠��E�2�߄`�0}�!hic�c������IN�X6~҆{�%�.���Μ�s�m�Zb�}��kt��Z�~����}xA���V:�*��R���jЩ@0\�6s�hn���S�C�4�����Ec��X�Eh�OE�9������ߡxn��m��U>�4wX�`A�0�1ש���F�)��]�D䕃/���7�o�Q�s���Uo�"�1sm�������EV�^
����p P��6@.�#�=�x��8�q�7�=*8P����I$dU��Ib=�i���%�͚�J~KB����nC�:�>��U2����-'ú�I�r���ݳ�"���0Iр��%>��t�V>ΤXZ��@��0֮QU��첂���9�Da.I?����{v����Z>�/f	h:��F�����]j�7=��_O\���.<�m����N��_��4� ibl�ؖ�li>���Q�����As?�ᓼz�8&g���86�m/� �?�a�S���6@z˕K�F�g��T���&����2B]��}%�0=&��M�%qy���~?���q	�F)�@5 �%��ih�; ���S;���u
/N�b���u��o�3󇣗n^,̭C���C�p����9��[0�?�[/���Sϯ�5?��0->N$��8Q�]@%I�Qz�L���/��p��'x��EH�J�:���t�<�0�5�y��ɠU���/�M!n���Ցy6�V|��cd9'��tW�9/�r��4��2m��h�&
�q/�3�cȵ���M��!ً̀������qZ�Mį����M�8����۵�����7v5`Nd�7��{���;�zO�[-{�%�[�/���^�Y��,�n�u�CfH�/?�����3+��v���T�u6%�$�}Ѧ�� sL�{�x
9��zY��
�m}͉�y݁��M�F���Z;��?��NJ�WS�i:�M	"?�qIz2lOKa�s�!��3~Q�X�B�p&9X_9cx��(Y|9���J�~.'L�ߑ�R�1s�����ca�ɭ)�M�"�V^�BD� �! ���ZBN��D�=yy��2re�[!y�p3�]�D�/��H���sc0�SK��L�F@��	�p�� �Z���F���ѢyL�c])66��R
h�E��G��Pڍ��XS"y2�*�|.c��d$?�/g@��T����4WB�WXnӁ�����?��c_�:�g�m1zʙ.T��S��v�i�`���}I��!낪%M�/�
��0	�ʮE;��R��XLF�3�5.���wƾNM��p�*1(�-Q��,T=8EYg��W�}�c���7G;��A��4[ �s�*�bQ*�zKҙ~=�= =lZf��T�?^X�iBd�y���л��9�%�!����ۙv��"�f�kh+�'y�<�癍\��RĎ퍎��T͗����>á��Gk��ⶱ�9��>u�& �ߛϝ�&�.�}�Rxan��:�O�e�GnY����*ǳ��<�i������ƒ��@8�B2�7��:����5���s�Ea/���Ǹ�q^�q����:�spFy�����嶻�;��Ym0�r
�pJ�Y���-��r`n�ҍĔ���g��>eC�=Z��g���D�搾E�U�)��� z��4�KΊ ��=�t5R��Ӽ����:'. ��>���0��'����Ȅ�~��?FЄ �Ew#.���0y��Ur;:�B%�H�7)�VF>᯿8��08��󡶰�7kMI\����O׶�4�5�h��Y_IF�)�J�~Tλ�^���K�o�G�M/ڨ;�SJ/�G_ �H�U���$�l��
K��j��c�jt�f���ܔW{������%0�й*N��܄�vI:�9��"0�	�*J�۫r��g7ED�	�1���v�\D�BvW�J�BQ	��	�B��q\���5��|��xn�������/��~���?��-�F��M���P��0rF��-����1�͢�-G����K?�Y�y���F���v���{1Ssw�tn���h�}� �zD%�Y�0aI���	���P{L�o2&���:����g�.И���yn�6�ᠣA�dH���2��k="?�[�)�z�u┺�ґ�<���1!e�Y���Ŷ���@�������C`���׌�q����	-�1m��#���ыx��^,���N�)z1
�����ux�����CS��f�&X�� �뀂�O���$D�M�O0�7]*8��%o,���C%��<(�e�z{T��S֤M[3EF��S��b��抿�v9���G�\y��|�q�WQ����C{u�7��E{p��ywA�ΐ;&#P[�y~�1�HyA`���`u���ͅ�rɑ���>,@�X9���@���eg���g~\�_e߷W2㖵�y�P+����a�u�2�>��s�~�}}8'��ܺ 7L�ݹ��W+)��0ݑku�k݊ߢ*n� j����N�/����Ndj�1�T?� P	���x���[��W�"F�����Y����_�'��
ϐt�����W���*b��;17��]�\;�6E����Ɵ��"�F�8���o)m�yAQ3mg��-	���g>
(sPc6;�)�^��ՉV�^B�����h(^,��'f��,E|��3I�\��-��+u�/_56h�_�b(��/��Fzi����H�6C��:���)�zq��T�5+R`�m��2w���H�/E6.��i9#`�=���k�
v|�O��<a ��ɟ]��J�f�:�6|�)���$c0�`"z�v�U�k+��9�v�A�%kӫQ����^%]�i�eB�� A�[W�/㟁U�/����}3��m�^��@�{���2/��o_zbbS�'�h7��x7;�>��A�&ר�3�.r���24>����G���w;�>W0�O�Pߤ:�Y2x�Y��E�H���k\�u��;t��!���H�x���$�D�R��ɂ"<�l���
v3g�W|4���v��Q�e����I��3$����\��  fIf1<QL����,��c��a���F�V��T<���˕n��);�PM#97��;�F��ژ�����������g��2���d��2<�P��?���"�Ot8@�����Cz��#��qIL7K����N��c��0�Ql��r�)f��;�~#���C�k(��!3<ؿ� 3��Y}R�
��N9�L����e۷�iSz`���f!�+U��~���`m{F`�v�߉,89��k�7̹Rm<���[�h���(�"i������c�U�%�-.`�������lw���K�2_~ �;w�b���K�f�Y��OO���r��2@����~��36\�>��X0Z���d�j�]T����., ��J������!�B���?�D/.U�n���B2��[CcaBkj�Y����K�>�]�HA7��XS��o��;�pq>����[㿐�,5����@>U<_*��G>��#���WdX�"�}�[aNUI��x�����3��J��M�(m�#ԸJ�Kn��L�b��Y@�v/f��>
�-�A*K!`��c��C�=W6����5�|����(���Q�S<��F�>�	w�Q74�h�(��k���3����%��y���-i�ʴ���]�\ϙ�o�
�֣�Q��渆A5���6g9M��U4�C�*�����7D �3�ż7�y-�&�[	����&|�r�1"���IXI� ��~Z�p����2�[��m���qi%rp���h�r+"X���N����3ʠaDbG�gɬ8<�S��i�Ő����ĩN��6[�Gn�_��#��jL�c�۰�=�E��tNЏJE�#�u<	�M~a��߂y(w��>����T,˝�>T��>r��iǖxq}��kq�5�����OE�l�����U�W�	�5���E�#��c�L�S��[�B�jQ���u��*� ?�eI~��m��-3���߷���^%�CNųJ����&���H����'۠IS���;��dM5�\׾�(���� ��^�A��G��i�������Ʒ_L@L&'�W
c�H7fǈʃ��db�R��dB�7�҇6d;�>>+T�.�eL�{��n1�S#��OmX�� /��`9*w{vާB�sn����h`���M�W�W�+|��8)#�LP�U<�?K�Ӓ�yϡ���zH ���U�Ob֏\��Ņ�"��آ!ʖg4���4�+	^��B����1S��Ϥ���@�H�8a)-�Ƽ��aכ*��V��?�h�|kzT�6�'���(Y;ſ��Υ?Ibs_uA*B�KXϐ��v<��ݞz�3��W����.����
����!؇�'�hl!<����0��/$�����W��;�=�����%�bn�j�;5`eK��w�0C��6�i��� ��s)����{mW#g�K���0��{�?�Zt�9����s���ށ5���D��nk2
�d�,�
�\�=@��� YԼ�O��/L�3Mְz�����t��ޙOX�f����\��&��;��'����eĜk�^����r"��2�YT_�拇4��d��KZ,���|[���l��p8=���`�?�0�?A(�4�M�ٰ� 5ȡqCi{��s�֭���"c��;��̡1"����AW�<pƉq�A7I8��8�u����_�"����7���u���6��=*�"�.�>���+�Z�����g�B�	e�7���ϋ��KO3����O���I.&4�q��Ƿ������+Se������t`0G�Zx��4��Tʉ���:7Ms���V��s|��h=K���?m��T���FÚ��t������Ω�܄o�z�z�ᖮ�A@��d��;\3K�} �{ފ�� ���Ð)󥏷8ͬ�2���e(��:���)b����SV;�c(D�+� ��n���x��0!�e5hL���}BM{�������V��{̹�	�#�Q<��;δVn�
)�u�( ��3qIO � @l[��u����9�Xϣ���ε��叭��'�i�I5
�6YDc�)�b�=�P[���-���@��ł}
�!RR�}{���fZ_7�1Jd�|ř$�ʪ()��6�f��ъ6x��GY�Q8i]��Y�J�y'm }��K��@X6#7�}��/�Y�/Ւh�Ԯ϶4h|2qގv��>�B���r������� �H �yY1.�7��t�J�����r��{~J�/�IY�v�"ښ���#ТX�%�7��M�/�0BS�ce�|lt3���!�u$���rW$B�$Z��	�2k����.��������>H�_yρ����#`&����
�,�H�
�R[�\�ؠ�hs�n(�YJ�0*%>���]G愘�Wj����*��;I���I��/���M��Ͽ��rZ�F�Ή���,uE�%������'�w ���\��r�To�̥���O�h�e��X�27�"ʕ�J兞�>�@�t�$�C�+�q36�NM>Pb�_�(z#��k����\�ٮ��4�pվ������s����{��D0�. at��e�����t����ͨ �|��/�P�O�Զ	���b����a��6=���;s��`��W�!��ۣ
�B�ar����O1�A�;��7>�"�D�����k�W���y�S<o2l�F_�f��𞀓\l����Ez*ֆ�Z�aE�W:4ID�����u�Rݮ� ���\�F��hF�eU��$~�k�Hj�:��K�lm����qc;�#�`K6����|yrZ�����V���YY��n��k�XrIxe>��@n�!��o�~ޓ#���p�� k\[ƦS�bJ%���^�@�����Fa��M0f�9r�%;��W̸�1��3��ؙ���Z:���&:.�G�Z��C��F������G�����\��^oKo�+[)��6��~7��ѵ5/^z���vn���c>��I�8�˃��%���c����Ϣ{�k@,_�/�L�t��&��g*AnH���Q?Y��	�Dј�i�)��&/��7��k�v��3����;I�=�%�B-Ð�)��D�3��Ϻ���+ȥI}�^��P��K�y�9 f����V�(N�''}���!����C��͹���;�K��p%�ڴ�D�c���m�G���l�ׯ��D߃�z�w�%�%���{y���=�:7���*��VNa�o��;��)�����m��h�#L��"��L�b�v�Dd�K7�C=����WdI�YY7��F����.e�!׿�>J/���C�x?��A�v����5�����b��I��8;&��X$-l�w���m�?]��c�P�J�+1��/���P����o��)alK��C+u2����U��8�j����ɝ���� _��ȣ����}���**3�Vε�V\�3�Ǡ1�"j�,�)�vۙ[˓��4C�`�I:�/���_��{Z�����L`��V���2v��ʓ���6Z�ݽ�eO"����Z$�M}��7a������T&�s���$�R��>�Sl��
=J/@��RfH?�Ҕí��t��K���V����4��a�A��x�O�|֖� �`��K)�]�-p����]4���2�1nD�����B���͐�YQ����V��'��y��:����1�OSFrf�m (㲿Y�
p�8�l"ő�d��꽩� ��\��P,��D�
�iAqC���3H5���qL��;JV21U��u�z�m���h*�_?��� ��6�Q\=���	U��c��s���[���~�=��x�+$K��ٔ@[T��)ƣX�`ҏ�����u|�,X���Ƭ&8ȕ���y�H�S7��`��k��n�ƽM��B�ȍ�S��z}n�?B�9�s����f���,�6�곋�5�O�-���DM��❑�v���@B}�@�@,%����g{��P�뷂�KC���1��P�ꐸ����}�[�����C��)��%���T.�qq�4��JPR��߃y$h%�2�F�q�;-�ȶ���e1C�:���j�$��d�"���:I��Ш�[�&Է�-C~�/m���gnG4�F?��́�֗+�m6�79�়�K�ȅ,��ۆ$[<4����<����G�b!�z����(#RϦ��]u	!�6��([cQ�sm�O&�4�ϺWm����u �"t������1�L�"�Z�e�it�Kg��%7EC0'o���D~x�1�[,R��xP�D0�:�yf��u���T��<�$,�	P��Ի2ǽE'�]�5�}ʋ��g�1f�������[��]�W��>0�!`�j(�8����Ж��ljP��>n�])�&e���@��ov{d6l�k���{<|<�b��>]w�yO�F���ђ�/�.�ػD=�����[e���9L]�u����s���7R&��?�����cgKꏧ���a�)b=������v����Q�N�Z,E�׵�_�C�ĄmSJ-ʸ}�jE���3�-��b�	�_�����6��H��Y|q3B�5`x�OK���K	m|���m����g�,��5��'ɨ�^Rv4:��JZ��>��D�1�z�<k���e��zT�Nݕ8���}�'����nr�g�����w�6�F��ee�Ō(�m��Xʎ�S�Zҵ}��f�3�j���y]{w�o�6*���ǫH#���7ݯ��=�&,�k������z96?-;j�`�%~z�C�
hk�|�/2��pH�{v�)T��!�M��{��N�J�53c���%/�M_i�6<��cV�mʟAUy����I!�r�/H	���M�A��;��J���ʮzAY�6���w���y�%�������$�ԍe3�	�|B��}�#2Ln#3L��. �>��R䇒����w��l`��#��߿/D5��sD�D�H�!�*�����Հ�*\w*��@����	g05ۤ��nBL�'��T<����61XtK��6����h�aKm����g��S&|�����֧�qm\���C}��J(U���T����!���dXy�
V����Rw�Aq��ȵ!~?�T#�J�՛h�C����5f~"}��z����哤pʘMZ��#�{Tx��N�L~�@����Q�kmz�`l�$.(M��FC�H�-a�e9N�;����F�#)����Xò�f*��	�f8�%�^�7����Cٴ���O-����wˀ�ju�s}+%�-��S��|�����ޙ�ٿ��uTo�����:��N����0�D�:�iǚ�<��!�~A1�'=����}��/��[X�0�%��U�w���S���U�t p��?�P���C��e��gĲ�T�C�s��c��D׹8!��p����<xbU�v�ل�س��s\6$��^&e;G�	�d3�yc��Hb�%�3��!�ho��:su{�RY���	�c��	 jAC��l�NZa��f.�M�}�m	D@��G1���Ԛ�0Ӊ~���ϙ�Ð#z�E�4��'�k������};�6x���~��l��^�����$=N��{�,ë��#H�~�?�@Vt�W,CS п�m����o7kc��N]���|���SF�r�����K���%����=�+�U:��
�~Y�B\��\�N��ސ��4L�>���*�P)�ro�rReŦ��
�ξ}m�kd@��=|M	j0�q\w�6�]j���"-ޯ�s`1����RV�����8��u/t6�%����\������<�՛�c��(��jr���!!�7P�����v1�$-�6����2	\vJX2
�5�Y>!Oړ��s7B���Z�w7r��˿�^h�f��Hܼ;�GM�8>h��
w�a��B�J.i�z�cP�5�$�P �L��힦h����*P{t��i�I��I��Z���7�U�JRݗ�t�\s�냪<-�Au�;$�%9���(c�m@�F�?��P^>�@�c�_F,>��[�6u'�k���Ϗ���c��=�t��J~��=ё����	kDњb�C��f������P��#l�����r�g�@��܅����KKxi��<�x�Ү��W#
O,��!�M���#ꆰ_�b1ӕ�8*Yo[%������9�`�у��]x�汇�+l�$_����Z�W�cQ����5��B�U��֮�����Tz��Y_fŬ��.�)ǎ_�Ŭ�L�I�q��/X���xu-S)�bJǒ�	�*�۴�ø�2���Qv��H�,���R:*�������4�>\}kx�E[ҏ�#Q�̉^��m�z=7������q6��
�C��/a�A_K}"��>�o�$�v��Egv�g7��Y7�L�N�R�a#�� �P���I,�q1%�	n	�Cd���|G�v�ˑ�Å�&`a3��G]����D�n��19�ܩ<��,/Ǥ7h�����U�cҭ�>�"�Bَ�R��M5r8˙}�OYw��\:�/�DIj�T/��E[�J�'�5�G�ah���w�;ӀF $��؆�wT1\����3�'� ��}�hlU�a?��=��K¡\� �/�O�[Æ�\��fBSQ8��bE�B:b�1�-����pG)����/6�C��E�y.�f'sڅ�۳�ܧ��`&O wE~V��"���P+Y���mn�"W��lű�p!E�����m����X�q���xe�n�L1m�ٱ��I�}�Q�J۪�~�[�d���1�m��h+�
�s�������Q�����G}�Hb���P܂�3Wْ:�@�0��@B�N_+��*7�ЌM
v�댬P_�~������g�[�t�2��mw��r��[����6�[b4���Vg\A�����]�(���&V(�c��AL�"8���~�`���ŔB����̲1q��6Vq���`�L��*���0S1��m�&�w�ROK
{ۍ�2�s1����ז���x4wTm�M7�yٔe!�§��ZU�fE��=_���}�g�f\��/����{�D_�C����Y�37�4���fT����C#�?��"9�Q�<w�k�!���F-N���^]�[f8 ��)V�D�:�\�_\�r�G�����!��a}gм�[��RyW+����N��b�d*�W�b��M�{�;���.z��ˌ��ś�r �������<�z�Rhs�Std����m�-���qU��1j�5������AF?���F*}M��N�j;
W�	���ـ�Q���fr�׷�-3��v?-[��J�=��S�'1�ot��q �'�c~��I��T��Y�Y-���t_�vp��&0���c�����J7 i�C����$��DK�א!��SL"]y����I.��J-O�.O�\�mx�\�����fFO��^�Z�Ȼ�<��G7����z>��J�BhY����'�Vӯ�t�U�_U�+�(e]�u[�	�p�"�ƻqF���������G��K�@��3��	���A�����xsǧa%�XI�T��ߧ˻aZ�+\qڏ��YiI�����'�z6����≻Tc�w�\3\�\(��^x"C�w4G*���P��ũYb���O��J��0�0�~�M�&��#n���!���� f�^�o�ڵ�sfI5�̆Y�
B��#QV��;�-��Ce�*��w�_������7y���WP7
+'�w��e
b��]ʤ�L�����K K�� ���Xrb�`%.��o�G*m:�s� B*b*�;�jk�g��D<
���3�>�Nf�I�%��{#�K��d�:򲴁Lp�5X��z·Jrbjͮ��ߑ�f���P<�̒R��Bc������p5���;/�}kp�}����8K�C�@O)�r7���/F�$}�Ó]A�fh�oh�����oo\��q�a=~�P�	v_�T����雬x���Ő-���0B]��.D�c�6xj�A��M��Ư��P^�%
�^|ܪDJ9�����1mU��GGbXk�a���(6B;y;��r���D!�����׶����!��W�'��{O}�O\�w�S�S�ZYV��E��	׷F���I�}��ەN	X)^s* �%)?/෍a>Î|��iz����-����EzO����B��']�k5��� =d����R��rVX�|���.af +��<��:;���s3��M�)P��������'�.iQ�j�K"�f�|��l��%��
�����A9Ҭ��L|�#��Z�X���ؚH���`�k�<��A.�NRwB��R�������RN�����>�����;���F2�z2��$�bL�+���	'EyK�d�~=0�pQw�����c">p��EI[$p&ơ� ���S#����s���y@8~@'vm5���+�l��yS�RԞo8���K$ʂ�Y)d.���2=w?Û?�N�M���5���b����܀nt�U
�N��r��t������x��+2JQ������M!@��d99���NU7�Pf�m)�n��Q�s���1�t��Y5�7lŪ�N\�^X���|����0�������7p�m��.��͒�i�/����3�,���#?oy�~9�I��v��CN�����$&�$�K^ɕ�0/��e�B8���
ĒB1@d��=BzYTc�����ܱ �S柟���D��,�����z�_+�z��"`�J��v���m}%�ܟ���{٣�BS��b�)XP��[nK`��kk�E��u`V����k�6��5�h�,�J#XuM�,�8��-)&��~��6	&&'���r5��	 �?=a<��4������j0s���Z ���eH���$O��w���0eWj���˺J�v��c>���7C�ŰCt&&=���F�c�&
dV�a���"��Ϲd�	|0�[��ԍ,<<W�$Q���URJ��dK�@4�`�$#�_5����z��}U����O��V�S�Z��3�Q�ۜ�����"JG	hH��0ֆ.թGU�[�n｀�YI���%Q��=��|�����}Dy�N��;��Yk	㖇�����R��g0M����P�:>Θ%[��B��!����[�WOߴKn����|E��c@Qb�7�" Zg�k��Z�����	6����ەP����s��s���xI\\���3]�5?g�ח���'�3�<#���U-"�>�O<z;�v}�X�DHR0���M�}P��%)`ËF���U)��=�<�gN(�Dh����7h�x��xT�{����l*Ͻ^�][���Jp�(���\(�,�LP�!L������9��\t5�`c��Q�;Eb��wӚ��ē�6���R}�����9|��lަ#\����*H��}D�KU�C��$ d6���������4��>����Q>�h�s=�j��1<�3'��#���+2��lV2�!�� �ͯ�)�z��k�bD�_�	T�l<��6�w�CM��T��T/k&�&�$���0�.��u㎈ob��	��K��;F"��v��K�ʏ���a`"�u }\2�Mj=�~�E�@��	!�$Gz}t�Q^EfL�����v���M���PJ�U�m���V������(>J���{�	ۺ�MQ�O����)���Ϳ�P�f� �h����oTBM��L����e����p�f%L��#�N�Z4������I�,y�ڣ^j>��Ob�$(Fs�����K���n"��ǷЗŽT��^�y��/R����qG�����U��W�YS�>Iw��W���f����b��t���8솆i�D�������ж����B�7S����\�[�x����������[���&�����W���
�)���+e�����*�lK���񥉞أ�&$�*�Qm�n-��įXP�Q&X޺t���x���kҡ�;߭��o�d���t��CZVK��LD/��_m�����O�=8����x�Y{T�H)��pA�U�� *Lh]C
L����=�	�C~lʌ��Z<KW�����8%0���M櫋�e��~��l���U�}��%� Ĥ7ĥ=XN4xT��zND��S��m"Sr7�
�ǅ�ye!����Y���ǌ]nE��q�:Yc<��x��SȚNC�_6 ᎅ]��Ӗ�|L!N�<?�0 ��s#O���U<<7��P��w�FB����~��W5&�
2�x��6�h�7�}�)��J�ǀ�r��Y���b/�����n��p9��k�����f��	�g	=�+��oh���߬.��R�$����뙨^�E��g�.����ny�لo�HV��I<��Gż���[��jśu1 h�i;���]m�i��+ϖZ~ ��7��{b��D�mV��dv�A�X��Mb����fn�lD&��=ق;����U���Uu �\�~=�DX*�]�gmq�ֈ���D�^�ț�>�%-���w:/k��� fQ����h/hFB��x�{��=��M�Op1�U]0'	@�a��c�/ �v��!��G:�H��5� �!�/z�b��x�!��9����}�+hE������T��� �%�������ń����dbᚳ3	� �q�l\�?Ju/k�-�6^<M:�%���R&��J�G��oPug��!�t�}q.������<Xy�?��.�Ț�I[P�߁
�B�wݠi�Cx �0s��@�kƓ?�"�4�y�	(YP�G%�3��?C<��j1H3 ��'��y�t#����=�5z���Z A�]�������*<R���R����	i)���V�kռ��E �^��W�Ȑ`��p=-�e�A��Px���<��ZSx��V,b)	J��<ڤP'�@57�����2���Z�Ғ�}Խ2�\c2�yAj�c���$�W�Rͦ�,���L��c|��s��o,�0���9���	+�G�ԗɛ�a�����-a�1t<�:FŤEQ�K�+���܈�`��o�W�w?��~���CȘ�D�9���õx^�<���E�	k=ěI�D]�kɹ����佌�y���Q��EY�2r�w�4(e*�4C�������X���}b�r��tc"���M�B���GR���j�)���� ��?�GD7��bE��گF�ޘ�C�0�r+�0��HS�b�	�Px�OF?qo	'a�����:^�Z���9�����(���� ��r=�e<���{�(���o��Z�"V/LfΙ��<"heV����g�f<F4;]9��T�cJ�/�2����v6�Y��}bK���f�t��H+L��:TΙ/�V�}Dٟz!Z�g��.�/s�2��^�*��@4�]�α�]�~�~_]�)0�2b0q�?VA��p���)4�Ą�
����-�݊����׺�@���q�M���W�����݅�S���q	5�;g[e�\G�D�{m(����Ѭ��Ƿ=��ɷ\�����6j����cH�"��>]|hM�/,�_�~P�#�EX��]�������É���]�QfC�CX��B��α�p��6ή��#��ҷ}Y���/>O����{c��}}��F\NU�U�b8�Uϔm�HEV�Y�(D��$FU�@�t��/�@�܅����WC�ry�d��c������W�f������@��Y��9#�3q�S|���?��?�B������'��$u��	0X�)'+�$x2�AZ�+|��Ӽ8c"{SN��zKL<����F��%�o2��l?R�zʄ�|�fF�I�=�.�g\Iǃ|f*mbP,���%UV�#����L�@����H��J����0�k����#� �,暠�h�_HkՁ��I.�"ʙ�,5��9��n��(?���Ybx`�}K�� X��d��0;�k�$�i�����>�P��w2�+�=QN~܀�Wu��[	�~O���������͂G<{&�3���'��V�X�?&��n}��[.��:&B���so�����f){)�'g����f[�� ͌�RQF��&����8o�!+����rk>2��?��$������-�$�s���Ǖ���1�����nB��$μ�s����x�%
�Y�_FI
c"��XJ7Vpd`��h�6z�3��9q�}R�_C�^0�Y�b����F��@��|a���=%<(u�oF��|0��wp.f�J.*��y�"��طl�����!��=������5>gcS���^Jj�a`z��̍���܃|_�S��9���~�����}���H�kQ�B�	�_�l'��'��1oi�[D69��̅+g�#�\o?̣�|�\Ye��0r��qa62%lfbCe�Y�>�et�߯[!c}R� ��;VS�a��yŨ!X�����I	ޛ�Z2"�!"�x����ʬͿ�2L.s�+��%�
#ă<Nݫ�@�M4c�����
����#,g,�U�q<+Kg�Y��`������X�>��e���
-wt�6��v%�.~A�!q�E�����?1OO�p��_�I��z�_U&/0���D���	��g@��z����8����	;��C�Ȯ o5�bD�Mǟ�Nޛk^.������]C��y�ߣ�u�@��	`�F��R�1Vײ[,.M�2I�(�|�V�w'��1偩D�7c��.l�����Q���2���nq���(��Rx��7����kB��s<���uO��Aw�-�m+�U������=�2z��qχє� mh �u��z	��v��3�� �� ��T�`�̓{j�]����a�,^���`���b�1$.0LU\�(��(��[f!��}��h�K�w�7�x�4�����f*:¶���倇b�2��������`#�<o�m��گذ~=;w)�k��u�Ŕߍr�^F����u��.�X�C&��Oq>�ɱ60��D>1��x����ӣ�/��R�a�Ӄ���8陈dZ�3ۇ�[0~�/�ҨJ�ګ��p���Y<Y�VU{\��#D�3���P���e�Kro�N����X��5f,Rʚ�9Ѕ��b���z1�`F'ր�'�H�*H'��CAx
�}�T�_�Hɲ�dkm���<&N�SX�RN૖�2 $��kgf.���3e�����+�?�eǇʇPI��a��AM|p��9���[�ރ�������]��z� f��D�l[{��?�n�ݡ,%B%`����@�}��`g̐�i&îJH�v�{��u�u��^I�<�e&e�Nv@�ݼ?�&G�µ �cH����BᚕD­�ڿ}�Ϻ���-V̟R�v},m�ax$e��A�'����{.��Jg�ݡB����R�S��O�~QV�w�W���?~i
�o���.�76�TY����):�/kh"�-}��|�;#�f���	o9�M��$,�{�B#*c��y��_�~�C�i�����K>8ݯ��xI
�T8�6Q����"��*t��-|G_����g�G�o��x_nP�b}�Y�F hp�e�H�0���ā#֭L�lc�rߚ���B�[?�u��S�ǆ�������~Wu�Vtې ~`la��)��L��0om���� /9pq�����zdl�����#�Qذ����R�E>�/�G2�|���$��R8����_-|TH_-b�.,\K�@k;c���,�,��J����U�^��℩,+��֮8���R,��$�RF�!��CyU*��4�h�򥓶��=~��+��Pخ©�\���[�G���!�����j�h��*Iׁ"�S+�bV�� &
�?��?X]na��K�R�d8��c$%�'q�)1�b�d�*C�:r���Y��5�gJ�����+������KGXc��|�t���[��乊ޭ�S�t]͆��gp[~�Y)����݆9�U��0�K���}�]OR���,`s��kdr�}�tj����W!O����0�F�Om�NF\i�-])��cP��A���@�p��>(�KN_Љ�E�N̼l�WI@�j�Z��&D���B��d�����BS�����xZ SbѮ":����'����E�w?�i��_�'|b�P�K���p��%�U��7`-�
��)د�R��J����,v�\M�"6�[%Bp���u�����5�t���#>�KVg�\�D	J�=��]��V8�J��;�nγ�1�����(�6�����>����	"������|��D#e��T���{V���6D���!�U�*c��ƴ�d��l�� �O�-��
if�3��@�� gO��	���'�U%$+oĳ���'�l���V�ꘔ�.��<T,#%]��R �x�!C%�'_TÂ�Q�z�W��ݻEӤa�C��9�2r����`	q��F�xh�P���#Z����0=����Q��k��A�cr
֤�w��g@E���r+H����ͯ�(��J���Nc%��ߎ ���:k�/�l���B`%����D�ZkU�b`O��z7�w��Dw�ym�?4,k�x�eA�m����#�ǭ�����.V���������7�kP�[NzDw^�,kU?(����pM��/
2���z9U�c��8'��ې�~}oq��Q�Ћ;uK(�� b[7|��p�ta���(�6hF戥�-�˫���/I�7T^3rSOb2K��:����dy.�ќ�[��˅�F�3�lj*��k�	XH����>s�ˏM����;$������Y�5�p��T���jV�qN�U]sK��Fg�R<��<����BfF�����<�O�|̿����h�;�
y���}���]��'f$m|t�ԪJ�Iu���g��u��A"���gG41̊��ݽ���cF��-���2���u�d�"�'���<���";d4��G���0�H��#{��f�^�v���rc��Z��,�����f�Y�,y{R�Ԛ��uZ�IXH)ǺL��'u�.�A���0�����|�������p����XW��.K|���p	b]&T�kh��{
�K�=�gEW�C�ֶc�5('�.���3y����EnG�o=�>�]����f��'�7͝h�uq�5��l�Y�.�j�]���eI0����+��MtK�_Is�|=��VZ���{�!�D����� LaI|�EEy�Jԭ3����А�vB��G/�%��ve(7(*To�N	�&��ˀ�U�⹯0��+o'��'2���|m#�r'H�����ƫl:�|�/S3S�OJI������ ����|�ﲘ?���Tx쾰��S
>����*b�,��g��F�a��?5_�AX�IZ;���+�.�&p��Z���)�R�4L^��p�Qm�*7��	1f��qt�@���-&�,���U�q�X �,��ů��V��6�;��dF���H��&2�W�*���h����V���Sώ����>.�?Nr�7*��-�MSL��5�!��s��S�3�����@Os�tI%B~R��$M��%��~��Q��qg�uYK���R?K�i>\�?��hEI`�aFP]���(X1����)���'#=�.�C��ʓ�r�c!�DG�5��q��{%7~?^���ݟ�Ԡ����y�S�Q**�6��]���V�3��4�����%|o���v���|����x���pi�����c���e=��>��ARey���|�6�3,0�Mz  �)���꿬qDCQ�����?d��	�s$������Ċ��D�ϣ���{��[<����غ 5�������;T^ ><��̐�t���Iq<�g�@:��R�וѦ{�<l�烿��ԎJ�"5Y(oo"h�w��|��9�@!��
��;%�iT��A߅9N0@����i!7�S��f&Ё�CM,����	��4u��1��bR�����j�E��%Ё�uv��PT�fr�*��v�����@������̼����eK%b�V��a��K��R��<P�Hˁ��A�±���#*1�����M�ȫZ1t���o����R�Y���[H����t����"�l�C�������@K0͕�Sf�3��o�3K��E#|<1���d�p���1t��+(68�N)1�ݬ����u������/(8s����3��\�����@��F����w��tXO�6�/������wF���8���	�͌��������dL�o����g�T��������Pa-q�l��I�C�q��W�es����t���!)�h2�*N�h!.߉�;�n�� N����e|���}3;�}�=P�"�#��wd1%Z� �"��(a���	t���)���@|Nē�E؃�NS�u7A��t9�8Yr������1f~�Q��^E���A�e�q�R��<e2�>1?�N��%f����r#�O���qh?�1��r�x�ל�d���C�Ė	_��o,͔��s�����X��zg�tŧ�����7�tt��oq!�ܵ_ޱ,ξ���4Q�LJ��|�#�Z�|��?mC'��P�6CIծ��g>���7�yT1T�B���?+�l�&3i�dZ��#�P�G��[����0�<h���|��e����<1�y��UA[��P�]��sٶ�V�*1��AR�8Np���W������{�7���}�63���E)!>��͓���dr
\i��o��n%{���p�\�!$���L˛�:]�} �'f��=� �g��G{�_M���l��*Rc�]�����~u�}��aE�aqv���Mm��c��r�f��SY��iFxdoE��ԮӀ�����z)���s�c:Y�jW�NM���d����ߵ� ����Ӡqgd��~1C�p���J�XY���� �~S �0�?�X)��oW��E�3E.LJi%4-�����'�>P��u�6�:��n����N�����)P�H,jH=3��<={:����ڇ�;�����ΰ���<��E!~Ѐ��u��:��3�]�&]A�e�����[;X����Z�;G����ɩ:m3%�V����-�Np:��ҁ�4��]c}�Pt:�NS�T���݌�*=u�՜�\����D�X�HM|57T�������Ǳ�]B��y�`��s�ա��d��A�3������(7�����Ǭ�31��-IL�(�?Rύ��m�8Kш�`��F0��V4��O�!��z �5��o���[���g�'p褫�"�p���#oT<
C����h�����	$G�@%���E	��n���Q:|�S$D7p��YWӎX�[�fƗF���-$�B'IR�e��`�e�k�7u�d2�R�I���	��-V���\r�p�ǻ��?Fvo;.��UWq,�Ɛ��#�jT b�\oe�,��/�GB�(T�d�^�3f���^-(l(KKRzSs�S��m�ġ��SoX�Z�O�מ9BHo#�H��"f�,��%�?5'Ю=.�ҵ�� �L
&���Ûv|��]i9��o���|��'=jP:!q����|��-�#uD3?�p9�f<V��;�]�����Ȅ��-*ksT��[8�~�ire���B��=Nh�8�k�1,�O{P���� ��.�=��W����l �ֵE��)��ß�\2�T"���);���A\[���=�t �n }��ՐA�J�͹�u��
��c�o'pD�<��B�2uk0�"k�Jy�R|6�i9����T���@�NŞۮg�I"aJ��N��t�zX���!�C�~�ٿ'`�s�y�vѩ{���\���֧���6�B�0��̙d��S(�"�5%�X�$ݻ��{
��p�j�hz�]B��>~�Pʥ��[	qHHXIs?�p>��l�e�L��F\E��݈�^�=x:�F|Uw��X`�\����K�bmBH�ێ9�#�ɘ��R$Za��<���"�M���7A�hŋAe��t�GDѳR��NՋan����Լu	��Fq��%�QO'C����v��}&��;$>~n�S]-���+��[���π�)�&�_�0�S�CF2\'�6�Wb��A.���%�f�����/�qP�%�(&�币�H��_d~$�_�J��S:����d�� ���A�SN���c�u|4>Jv�L��������~_�!���Q�"�fH��K�s�L��W��x���`B��̭*D�#�U����IcE�7&���o�-��NM"�b���u]]���sE��.�����	�.Z@��g���I|4j�%&�3��n���:����2]o�'�0,տ�46I��j%P^���IKo:��S��O��ץo�3�Ss����������	���\z���Zǀt.�@(0�T�oP���i���|���z��><��F���7����f̏��b�2�M�H�a��[t�L�'��_cU��OsE����YC��,��f�v�c��z���h^%�P�)�ՄV������|S똳�4���]���@������0I�-�B��t�����F߱%�E�$i��q?˚]�*�y�M{�Xq��b԰�?ZRT���sFJ�]�����쭛܄n{����Si�#z��i��fQ��P9c�rq �����[0��
�m� 
����&/�8�'�fR�Y!��qU�W�0���p5�q(�zi�.��T��e�C��M�����J}K@���ӣ��/���Y����c�E%sld�f�X��9��v�_�=X�֬��5-����*���
��'\����h�g���W]���X���
�˿�J��C��9�K�SZ?}����o���"LG�o��?s�K^�s�%H��Fix�A1|���.��������-�:M�u����e�"����S�d�S����W�+�B,eh��c�lJf�X�"�-�*}�������ژ�� d*������}1�UӆM�,U}!�!N��3��V�f&Jacܶ�;;�!

�;�&�,��7�.lBл�����4D���}����L;6���Wȗ���+2�
X��դ��4��#?�g)tO���T$%��^��`G�#�k�0}D�e������DY�����zk�^��?����$u1Փj��R��(^D�=���}��v?�a��71XӉulܖ�����-����]-
�Q���M�n��QL|��@�Cz�`����0(�#l�I�[�{'G��\`L�۾C=��q@W2M7R��!t-l���j�A
)��	3����<�U�C���h��ܛ�:�a�"��%oѽ-�@p�O�L�y/ t���Z��N7����䡁M�$i�����La��F�����9`P�3���Ef�?�J��Mn:�U� v���F�P*p�u���V���Df�g'��ϕ�S������,]��J׮o�ϵ`-��V��\�1�S���¯B��R�n�6���:���XIOvk�%�����R�lO^ᇟ��˳�W������O)f+���(L�Y�^8�^|e.ej�ɾ�M2nPIq�%�e.2����<�@�J_�']��HLN�ܿw|�,�b�/4��!!��srn�����|v�l�ŋ�c'�$�[�ARzc�v_ݻL-ۿ\���T���k=���J�p���= �o�-��m���*�9x��@�!�{����G��k��Y�"�x�s���/���N�	�'��Z��l�T	8h�|*6�1V�bz ��$'�C�[�'rGx�'�R�o#+�Ϻ�,�= �X�֟r����	�s.h��ШAѯ.��7�8O4�R�[��b���}X�b���X�h�����Oܼ�����bYf�WUEF�`u�6��J* �QmU@�_��[ɺ-)�$��濵Lg����G����g��\Za[v�k)٣9�eG����W+J�?v�'��04�<f���^R����(:9i�����;Ӥ]~6$(B5A�ڟ�+�r��~�/���8��K?�O��\V]R5��>�$)(�	;
��Crz��{��OZ����T`9�����-�0�|�s��P��̾������q�Y�е�a6��`)i��<E@K_������Ғ!��5���~����P� ��hp��C8V^���0��Z�����o?���=�Q �K�Fv���JW��u�8�G�����`}Bգ
�r����5����[���G�+��I��ћ�
���Z��}sk2!���-F����I1'�/�qGҘE�[:������>)�����Q�ϢF���)�O葏iϐ�pk{���i�KB�2��9;f�|n�<ȸ���4Wy:r@j^���Ȩ!,8�Ϳ��k9>��C%�c�X�����.�ib�:1pf����b�qG�L����)���� ����G�O�9`��f���,=oEF4�[p��=�E~8\8
k�~�!�}��^�o��!V�����&8��<��rμ9	���~g���}������#�1Q5*�߬Ԫ���U@{��E�)r��t5q�m`C9'���wYf5s>gGS9g�U�`̄���зU����M]���{��%G��Gj�|[a	���
�89�ɧnbשW�x�q��H������ct�9��f$�\�o��(m�||����a��J�y��d"l�Bk�&76���h���ugCD b*7��,\��^7rـ=�p�ov�6D.�S���. e�����⧖�[5�&�z�D�!yX�IB�d����'J=	uU�r� ~�����o bc���`-���@�,Z�\Z�r����$Ntف�a���p�O���/ރP�z�Dظ�O��	T�߇�O C�K�
^�����W����C�T�K1Z��'䧁�(<��&I3d'|�Ds4��QC��7���߻C���1A��^�ԖȊʯ/XN���%��_B�k���ipY��r �F�zKX��t(i2����1����X��*��t�qĢ	��(5�(�>&�)tQ��9g� t[���<Y�,u"�%$VNu�$��fc�q�� �a+�іż�ֈd��|{�
S���2a��-�_��S��Dف��-�*"{�i�6������h�j�|?��v_i�8+�{��5q����*`�o���}F+�B)Eۮ!��u�=�ߑ��JW�r��!�q1ߝB�'�w��kL�
��̝tVkyΑ`n�)���~UЃ�Q�Z!��@�%gM\����1ع��&�[~�)�&&J@$��/MX���{��UҾ�� sf�<M�-��H��8-6� 	Z"�{䶳�(�
ʣ�a!ܹ���:��0v��η�!6�1cX� ��$��b#\�;u��2
1|���!=�ߍ����X�������0R����~�7���9��;���pp���.K]�kK�O�k<������t�Sr�� zfo�u?J�]��5ɲ�1��W�����ܔ�
�9��U��a�Rb��}l<���Ӟ�N��)�͚1��,�o��f����-��L��)�@wڋ5'�~	)@��1���(^chg�(�˴{�Sh��I�nZ(���	�r�4�u�v��h�Q��գ����3��=f(j��+&&-���s�Y?���+>��q�F{���x��t�]��{}�z�R��$�G��D��;sR�ՉG�g�O��鲫D�#�6���D4uO�apZ�tѥ���:�����Vmԇ�@�%?����)�w�?��p��������t���� ��@z|WK�r&&Vp�X)�E�����)�n�j;�nD�"����+x������>
_�F*q��RD ��ə2Wb����O�}k��V\ܿ�{�t��%⣝�
!�p�54bĀ��$Y��A��h�.���V��)��j�	�e#2Ӊ��R���r��~�Q�[��9];��sr%��Y;��R���qy�I�>4��~�;��������4���������{�L� ��\J���4Ǝ)��Z����[.k����&�<���u�>Mc���$ɫ"\>oA�h��#���S[�u5���Q0�O�ws_`3W��9���ha����~ʹ��UW�::gtYV/��]��3A&�c���v���}�˳�_zJY*m�3�3S��#B5�u�5w�#� L�7#_�<;t�n�y���m7�X괶^�Dd��c�Lec8&��ͨ�"� ݒE��mũ!\�SUn��źo	�^�6�"��-A��2�ޫ���v��wQp�W{@�������S���5�Ll*@M����s�W^6�<·�.#���J�JM���VJ����� >	��cS�r��b�Git�鎄�Y6c=��'4�mv��2���6�bp�����$6ກ8`�?�M��(7��3/� ���x	)GYh�EY�j��O%�J^�i�}k&�슘��j��\��2� �D~��i ���Yc/Oy^S����!#�:��?�r0fe���>��_ ��!u���]lB�xB�B5X�����,.��Cf8�1wM}����Ŕ����t8����m����h����ǖ�HDB$����+}@�vX;�0p�>} rD�w!��I��>�ݫ];?�J}���d	����Vb	�eL��[��}T-�I׵t�h��0`�?!\�w�)�jǔ��:c���i��Y�E%�i�a1(F�}�(�A���E�G��@�'��&Ϛ�/������h��Ƨ���6�a�ŕ���hR/�N]m8H��IEΣ��̉�hv��P���8���,�-%,)� �$��EC�T�,@WsΡl�yl�d�S������.���ϣ�	��z��œ��&E����B8����ZU�e3A�߭T�7�V������5�E��uW���ژ]-���qA@(�t��
��り�EY�	ɳ�ɚr�\�_�S�-��6�EZ��:�y�C����6��SSj�ɶG9V1��ݓ�PĒ)!:#L	�b�Zt$�dW}�!L����e�!�M�/���a���^������$�`�9ϭ��U��=��i��CF�T���tMr���D.8�/fI5��)���$�O���;r�?$�o�Y;��Ϝ��A�g��js&��.c6�4
���d�@�Hҵ��3�F^j.�S*��&�ƝPԕ�X�Ԓ�td%����ݮm��c�l�N��L�;���>I�qj�M��	Bl�w��`R�J��0�]+��o���c�D��(M[��'�;~��p�(�<�,�Ԯ��r�}U?"�$�fv�qjJ��r�4��Y�L
��s0�����{n�8���,��d�V��k��Do1��$U`��^hI�Q���6+S�(�a�c�YTH\e�a����g9�H_�~wx_�
!��A�
�y�&�O(�`G�y��S*�l։m���y�#mW�!1<`8��oX�3U�Q��ƘA\%QB�Ű���-��%�v�>�L0��VV��E��E�6�$���`�k&����9��� 3����W+"-o�^��T-p�}��}�y�;�ZYZ����5]��ҿy���Q����?7�eĂ; ����|{d�.�����a�
91.(�zyD���z�..�lN��C�qp�3�?C�X�Q�}���8%�j�`��c��{���8,}:��Cn?p�����ə�a9V�GJ���_F*��� `��C��Ɛ�P��f��D'ݲ?�˪]뫗�0i%�����℀��y"����x,�����~K@����������FwEI9dL֙@��<|9Hv������a�A]�����V6��z���-<��1��1��(T@d=
��ve��Q�l7r�7�MXY��U�)$Ȑ�'
��m��0�����_@�I\t����Đ�>՟��ODV5��r����I�P�Jߠ��S�.�ꣳ�"]J��,eG%�Ps���1�[��.�(��7�1��`�.�Mecf�J�a[ѝ8Z]�|��1�*/�"
�g�����<�L����@�0�y1���I����� �,�TW�&%@����Sa8��`��H3Ka�{Jן2��C�a�������E�y*�m�4�ӸS�-"��>w�*�׋�R����	B_��2f��f�|�[2�n��dXN��w�� ���cv�
�n��u�ҏoo��,����r烱�/�O���{�����p�w���E=�x�+M(����˼F";�Z��f�m��֎Ŝ�1C}�����B^��}�-Ԏ�����l�+�(M)Յ���mL�oV�ڥ<�MǫPe��[��N��F�]JZ�p���PD�{����cnq4=����[�t�u�_L���9�e{0�W�F,�+���O�:^@8�0T���O�]�p0��|:s�Y�/�1e�,a`���a��2�8�ۼ/K�9��3��,�N��a؀Ml����F9��i��\B�dZ�DL���i�I{�J3I5������ʵc�����_�E"������R��`����O`���µ��X�ԯPzx�Vd΋�e�xB�m��&Dد���a؞=�d��{	ӿ4�*~�{�9H]�T�C��F1����չWrY��V�`6���\����e��Pg��>�NԢ��� S���/#�ߞ�~���A�:6����U̨��N&��V��")���}���i��T�}�J��	�Fu��ג�%R��x�k�	�坫np�F̒N��N�8�K)h�ɱ ���^�����w���# �h���!~1vp�Y�T��T���V�ZF<� ��s��W���� )
�6"�v���T�>ӻA̬��S�k�ČQ�Z��0�ɗ#�%�Q��a���.;�0�$��p�o��-,$�q,2�Y;���:i9+XB9]@��i/<�ZLb�=VF���	�������!β�E��XY@�vU�~�����%TGXM��Q�('���Z�Vr�X��]1���L�#5���������}���3yUD��}H���1�Jv|ܻ[����I�R;	�J�̓D_�d�$�C�{ܶ�$i��V��@y�s��sSkNف%����^����������n&�UY�=��nNuD?{g0��|nf�X��W�f���U0S�E|i�u�YAY|kh�(l������F��7��ZN�6�ƚ�{���j0��w�"��	Qf�taѦ2K'�5F]��z,��"��=�C��p}�K�0���^SB.�G;3�٩<,���L:B+K�F^�@}�
��L�u	�1g���h�t3lQ���f�m,h}�p����$���*��[鸆�*s����?����m-Au�*�׶fWQ<T.�^�f0���Њ���Rhy�����R�i�CEN��%P~tN2�)	ݮ�H��s%�o��u��m�PIQ�w��Xn�f'�y�N�u@y�%!5�y�R���ؔA���ȳ��}Ri��`�m��M�f?PK.�A7�֔��U�J��\%�+:��{컊��ľƣ�ӽ�U��Tv���#I�1�Qm���+)>��g��{ԟ�U��� IA�pt�ϗ��$B�	]_��7��2n��; �����'����Z�#Xu T�
aB��i�k��v����[
���*ł4�B����T��w��cI+K��ORD� ��P��xfί��~#���T�!ZtAhkh8�4}R�C'���cl�XKi򖓹�#0X���iwp&$-�-G>�����w���F(��ˊ��8=��2�{� b��\R}�;	�|�!�5u�r��J�_jf�|�~�\����x�j:����Zb�������Ű_�����'������a�d��n����)f(���-�Ӗ��gX�=3�"�tpg�aL�����/n�����MW���c[f-����N���*�.�S.#�v��8�6��)q[c˘�f�?�E��G�I������	�@s��,���Q��iӛ"u�	n��7e�h&�Qܱ�q�J���v���& a���f�C[��0�ZR���"�{�.�'�P������Er5�'����j�HE�=���A�O��!��&��!T�xp�%�����&Q�8�p��T�_JE^j��s��U )aL�uLwt�9(����=�`�X���(e�ATWɞ�F[�]�:��Z��cZ���&��$.a
k9C�^JwCL���r�`��kbYX���jEZ L(�"�y
���j�|�It���	]�"z��k�/���1t)1���U�d)xr�%��;�R�����czv�+��,^a;[�XA�sԂ���S��W�͸��d	�4���Rz�����)V��3ǯˊ����D-(K����Ø�{��Ik�. Ѓ�X~���?��
a���`>���U7��?��H�d�FA�d?�-���^tM���G��}o��Z�t�y�avu܄%ޤJ0D�!�O�e��R����Z�q}�K]�&���oX��F�R��C�LR�pB����D�j��jc1j��;c.0׻��8�#�	�� �r��O�A=N�b�KFZ]��4��^H°(��Pi�h����魖^���}X���9���DWo��" /���L�43�(��Q
A�p��`{���K@e���r�мZ�2=B��H�`aB<����O�c�4$�70���j�$���Qԁ�M��asӃ=�ȯ�c���|`Pl��B�=07�@������RϧTT�ʰ�x�[Z�Cш��X��k���
�p�=����?T�G�$��;]]��~��q�na~l��¥)9+��S<[W�#�N�#n*��c[
ٽ���a�����"����g°`{��3��- ��v-�K���*�e���G��ֆB]a�ю��5?�pF��F�)|����>y��d��0��U�����%�_����y��H:���B6ib<�G�<��[��_�	9~ģ�����/��,����1z��~	P|��G�-���r�ӒMW�6M��5;_��܉gR����S�_�� �\3�,hnV�a4JM�R�:�O]���k���j?%u)���E����&>�����I��}g�d���-r]x��
a�={s�A����V�e����m����B�䆦����r<���C1s�5����FI�RUkρi�� 6"����Y�ϑ�j뇫]��r�؍آd3�'���+� ����5�!<�!�]�?��Պ�J$�3��3M٧r�f:�ʚ5m�!�ė�9���TK^Y[a<ؒp��8��{�8�t�Ι�VU��5�,V�Gi�!oq(�����4v��D��o�Xi�/��D�wռ��D��s�A���$Sv�����`�o��8����M$9��V���\��[z�Vg���
!��XU�F���92X�0��|�#b�!��#��
�/�	��wM�5�-^[����6�������A̹��p����S'Z�J�e�j���a�:�\!��?h�/s�N8q�K�>@��p*7Ni$7�>�(%l�y�*����a�`�����c����)�� ��5���goa6Q�
o����u	������1�]0l��2���[S[��q8b3�����䛰����93�!pT��[�l+D�+�\')�teVl�R���-�X�\x��`����X�qv�\?L��	���������������V� 
��שּN&��g������������d:r������NY�ȗ��4��O��W��_^��:�0_M�|+�Rr	F=�46�0�59��ĆsINw�~��S,55�W]t���+��=�������[_�b75�Y�d4iJ��8���B�b	�G1s��B��_����x�=9E�l,�O�y%���UT��1��+ߩ�<���Ż�]�SVMv�|������_����A�C+�b���b�=�?L����,�,��7S�~�f1�)#��8� @�n���1r�{�u].nR��Љ�3;�5��}#����U�j.L�ȫ3��=SoC�wd�9���9���~��y��
�N���p��߯�8����ⵆ"dg�[�-X١� ����=~��[�
5N�9����z$�%��r�}�śp�!����W5{�� _�+���ۅ08�A�����E��F���e1����� &�S[�戀^1گ���.���	����(���w�W�2�m�������\��Z=N?���+��뭢�d.���FD�U�/��7���aZ+�u���N�4k��ci�_0�
�zd!����^[���CC����8�?j4;%n�v�*ҏ>IJ� �cU�ֱ!�|!���,�w&OY�� ֎'�ɪ+Y�_jF��u0m��l(�+@A);A�k�L��fh.��R:�x�p�b�=��ݸ�(�]��bQkP��s\���u��S�Ѹ۠�9����9�xY�"8~���L燉)���j�ܤM$�|7e)� º(�B�-F�W ڶ⾦#������;��(P +�g� �z�{
Q0��z��>���>�p�8܇U�	��Mƪ�@�d:,�����!��}���(Z���L*g��R�<�l�7�<
=�/�()_Q���Lf�7�Vt���e��0�"�9��tF#x��k��E���S�l\��9A�I�ӎ&��󉇗g��j��<�s���F儒������g�<���O��=yl�jfsi���:�����C�/�qm��Z���w����M� �ufc�۽Xh%��%n�T$�Vjm<.��6��CV�#3p�D�J���|֕nVRs=E����on�g��`��M�}%Z���( .Mx��6���H/^{I]����uB��%]���$]ӀX�-��e�L�Oy3�Tse�-�o�|��v�+�J����zb���NjN�F��e@��%&����7��s��.FTD|Z�75���7�q1�c��ڮ�eM=���r59�6��C5'��#���s�i��u�u<���Yj :����~.��x~���	3	�Asw���<��g��e�x���ӕ�~=����Ֆ�fq��Z��1`h����:A�j��_<I��4��E_A��7�nF�(�<��S��8��)�w�,�E�jx�a�m6�t��|�����t��af�ꬖЇ�zzb���aܕq �H�v#̠(�.]v�n�~~��J�Z`Gs��L�N����gd�1f�~��V�ݘ�^�Q(� �mJ�3�.t�Y�Ĭ�e	�|^�s�xtoU��8���1Թ���g�8�1� w��D���*Tt�kpns��E�a�x0rnL�"�!s������ �>/�ܪ9�+��+���8ar�"�K�'���X�.Q��x	�|1�&��/+a7J
L,Y���c5���l�_j�>B]=�>;���qy��
C��=e;O΋e u��o,B�yI��Y:��EZ�?ʔ����2�����7v�|���z�Y$j0˽M���qr�˯Y��o�FT�5�&�	rFf���(��40i�	颲'���?�� ݽ���ݧ�,XZu����Čl���	���i}+2糺0;]7�t�
Lz1�T^:�&z�
b�јǿ���Z-tHVr�p��ڤ�����>���ѝ�'�X�mt�`��"����:�IR(��iGox�lߔ�~&|]�[>�8���y�1N�S�5��ߴr�������JFGU�����9�?D��k��Zun߳��ajj8�$X�c1i����˥����oi�Cw_��j�Z��Yc'�/ \�~(=?
���1 �rojQ�Sግ�?��7,��o��׼c�0(�1"������s� ʇ�T�������u�g_6H~u�2ݬ�W�P�y��2A	\�q�_Yiy�'c1ԡ��)�������t�$A��[C*�
kyll�g9P�sJ4q�6aOڶJJ�^�J���eفz��踚��!�3���hb�[�����\QE�ǋr����x��9x�Q�Y���W�2�|���}N��Q�v���#t�� �g� Q�޵H��V�g(d��[4gb�VG?�"������<g�%���=^�nňhϧS{�KtU4^��V_�͇��
u�[ 	;s��ut0Y����;cŗ*8����r�咢&�X3���c,�zё�@���G�GDIn;��TI�{<�wxd߳�_�okQ�0E��@*�M>�4����v����Ԩ�L�И�MOg��E3���xp�� �o�>�_Q��� RkuF�96�Zg�A2�ZL�����۸�UͪE�{��C:��6���9K�፾��:΅��ӑ�]<
b�S�ڃ/+�d��:ӗ�a.o#�O#G���5��S]�X=�/�����s�����M�����������<l�Ē�eb'�e6*_-���h�|62�E^뽫rn⇟*��Ϗ��]W��X�Q�9�/��j�v����^�"�6���3ޏ
qUx:�=�f$�H��3T8�:�b1
���mN�ξ��N)T�����J5��Ý'��Dt�����~���6�N��&���8u�gF�ܓ#�,�/�v��ey����;���)[9A���s<ʱ'��`���K́���7������qv��F!�#��a�9Rj��L�nH2�q?�ɔ��uR���᧔V^n3:�{$kT�p�^�K��Vx[x�٘�������8~R|(����-?ET�(V���Z�y�xF )BHl<E�����#7�6� $֤dL�s�+	��Ui�+�O���/���B�.KS̗���Ì`�M=Cō�aO��: ���M�˰8䊍7�����s�Fa�>�Ta(�Ð�<�Yz��=3�W�y��)��F�Y�~�C�=�jz����\_����d�>}W��Qn�6�$��6��+��T8g=\d�Ĭ,�T�(��@`.�0B����lWh"�[��ͥr��9+fLZ����U�n/�
�W���͎�ō��:R�U��	IB�Gu���f�|f\I�H�uU�(�嶈��gT��-jX�ɰ?w�/%d�1W���NȢi���*!:@nYh��-�G��aH�P�|�@�4�[ͧ�b�X�TP9�=�����>L�k��ډuaH-;�*N�Ly����6�5X�snZ$�	�j�<��u�������J� �:@�fZ�������N��Qs��q��%����n�9��h����Ե��U�(�X�8,�@+�6�}/maJ�l�.ռt��S�&�A���z�i���D�E!ƈ1UM��ܟ�M�FI��g�3ַӝ��]��n����y����x�u=	ɛA��%���"��I�sdUY��ܸ�[!�Y��R����>��Gt�
 ��ർ��#�o�t�-�Fk�	� ���,�s�lW�&v1@X�k\�z�Ӡn�֌F2F&z��<ǉF�@�ζ�~����Gp�p��=�ȗx\�Q\���F�l���S�OM�T��
���=x{������������}��G�0I��n͞�Gd=����/{][(��5��-�����02��BU(Q�����SRN��}�l�srL�Ï���L�����AK ug��D�&�-�m⺟�4y43���Hn51�P���[����.��N��J�*����\��]G\
��:�	����*
n��ݗ?g�G���%�pB]a�u���.�U+�v�-#���0nz��[gKN[�j��u�%�$���=@#��vF�荖cNMsI���"9 $ؠ ���׼��RG?p0�*������6[S'�\��U�ȤsK�K�6������ŶMzü~���"^o������s��b�9����:YCa)�]���H�P�0��9!!�M���� �q�O�1?e�%i�3�_��/ڊ�!KJ.�$��YbvX�p;d�3a�xAw8���@�&ꊅ��j9��:��ˮ؛�͒2|+@�]��Fb�x��E��2ݶ��WKr�@v�;������M�N�e����_���0�D��zk���ف�3�)�3m�ڬ�>!^Vy:2z���ͣ��t4���-w��\�/�Y?���a�"D$�;���	3���ƈƅ}5��~e�%ُ��̴�V�%Qzh<j��hK%`l��wH7��|�hO�neYϺ�M; *{�}{��Wͤ���&Y��V�/��`C� ���?z�g����#���N��ɛ��l�l땍�A��>�\�o��P�"F �i���=lC��O��āg���8��?w�8_9��SJ�D����z�@|��Ma�ot��Z�{6��ׅ���$n ��]�;��A%<Љ�_�Eh��w9��G��t�h.�����
�	�Po��5vh��#rO�Մ�$-j�04wC�e9��|��PQ���9��2pc;r�������R�.�>eӷ;����鲦٩Bt:�+ޖ�p��nʫ2�P�� �a+��~�'��i	�Gȟ9�`.�QG {��P�q�i�7"�opbU��ha�Ï��N���+oC�r�E���bkۻȐ��{-�V�)G��p�x������+i�����~��>�jg�/�-]�De����}��2l/�t��(Y���<u!��[$�^�(❽#a4ok���z��cFːTd�\��a3���Ӡw��q%��>?�a�����{�2��V��
t=�3���P���IZ��&�����5J-b�E�C��J�Gfje�_��0�9������^��m���2�N-6:��`9	$a6�4�}�f���0���{�hf�]��XC�2�`�c=}��[�����[GN��z?[E���N	+�[H�E�����T�1�@�UHN��GL皴 I	�}���ta2z��{��M
�tS�����1�7����r���ݾõQ2��ͦ��A�~v*Au�Ư��+w��3;��s4"���8!%l�f��lY�VBd��K��$`���ĈMk ����>�}[�۴���G�~6�	]ExS�ν��]*�����4hYc>�g�6��x�@ �p�!�ٽy�g�F{ i �Ho�~$�&��	dTQ�γ�'Rz�<����oRSRs��q\
E*(���t��P1#Ǒ�}��k�g��d)r�oL�aYZYq���U��;f��ce�NRq_1�G����;�Ske�Έ��ĩ�Ԯ"�=34F�Ln��CM����=@��7�=%l���/����X�uSғG~J��Xi�"�e�Vjh�:&�-8_�b��_��Ar�XqO�_LV�i�Kv�ք.�;�m3��N��
ǿ��R��>�����9�(��e��r�Ӣ��D�aLCs���/�uo �0��\>�W1��-Y��FzfE׭_�G��`�'}�p��G��4��*��B/l���R���o�u8/Ej��1!���ѩ@G>�S3�u�!�wj��*F�3+qL�9����&���z�	���eJB����:q� �i{��;��"���bp�<NИ-m�w��)l,�_�(���J_,��[�'��H�Ó��DO�-A�k%�5����	r��j\�khz�f�{Ɩ+��,���5y�A�wKU�W"�`+XJe"UP�:.b��i�mn���%��m�k���@���q�fYt���j�����]V���&�'�m�؅8�r꤭vEC�n���WD�/Aߋ����K\��ʲ���xGI�d
�X�� Qo;�&A>�k>zHD�dT�`�K���v���zLY����\�К�+�?8���χ��g&�V~��GV�AE�i���p ���V�k_�2����u�)&�W�(��"z���U�
�����kZxo0�H�3���k�tR���h����.vpI����nA������G�����慕s��&�򣸏L�-��u{�H�)n��v��ɂ��C4�d+��n���#5�Կ',G���qv<�~�ۂڊ?��J)].��a�B�PA�q/�DU��p�a�PYhb9 ����#��!f�-�s�|�LT��/����K���+,�����e [S`�܍�����%�wKs3B��#�j�E$�<���j��w��C�tk<I�N���h��O�g��[�`�ZO~?\�d�u���52�Zκ�5W�E��I��;� �K+����Ų��_���"�A�C��e�i1�g�-�W�h��*g�}��{^�C���m*����
V���(�RbS?�ǿ(v�6��5���4�h��9��k�>�)^�h.���j��YO"���p��+���"�-�re����������¼����H@$�m�@�S��c�2�(��ݹ�_HFk�O|9rY�Ռ���>��sa�?m��E�*�ji���k�E�U>nz��j/ڬ���Է3�9�[p�XW�����#$�f/A=��x�2��y�˕7s��gTε  �H1�/��4>7�z��%�V�Q��¿�ߤT�z@�(eތmt�u����d��t���dJ�AB�1���{[��������2�O���o>��s���=L\l���3�=Բ���	�Ɇ��ZY��_�">K;h]�o�G�R������F^I��?ǒDrR�����R�L��9�U�	���럾	�d�J i\���k�"����0U<���!�Y�L0F���B�R��|I$��bH�IӶ��25�'�A��ۮ��\g'�X�A������9�`6��T)��N��Y��ȩc�ꈪʣ��� 9�S��� 1I��^7�躲�(|��^%�B	DM���$=������v��4�r���I�0��W�x���Sub0���O��j퇄�@�ɻ��~G+j>�n�6��$ғ���"N�tb��R^i��H={�Y�G�9ό0�H"�#�:����*���������O�D�fע��B��:�#&z�ܳn+o����g�sx��h(5�n��������5��h��c{�B�ك��DļH!5�Q&��/@�>,b̀Rӹ������E��k���,���ܮM��yϝ23ױy�!r�+L�=*��	wr5%Na��m{���X�J!��ݷ�7�@�j8F\ƞn���	3:��(���؈����N�	D�s<E[9���:���/7�P�����y� ��[�{�렙߀��ިd�n_U�36%�P5�T�ʐS���'���)@p53�;�����$�G��}1S�]�D��G�K}o v����_�gH��84S�5�o
���|3��1���Ae<0���k��$�cG��b�#�j�҈V�bUĊ����"���;��I����6�f�d<i�N��P��Y���H���_�V�5�1�0H��{=K����\O��.��_�skLO��9�Cp�=�蟝1��$��4�gof������D�/�����d��-%2%�"�]��9�@H�H|�2#�W!�־�b8y��G?��/�,{n����F}���~�x	U��*�?B�+	�`ĸn��N\4�Q���/��T�t�%b!W���H\��l�����A�zƚ� �����UW�i:T�Ѳ^������7T�͞���aG�(!����)�$2v��TY+����3���},��-8OY6p��Y]oO�%E�bm�"���]��F�w�8 #N�����E[��6dT���5���;AV��a��Om*CT���~C�'m��Z�>(Q{ˁ}ͥ�]�6Q�����!m��֋�x_��%Ô���8�q��6���P�e�N�#i�`#��y������/��J��-X�!q���Y8Tl�Vb�%u�]�B�LKU����~KLu�I�����\�ۨ�Ov��LRI2"�9wL�ձa0� �{��V}���q"On���}u<��l���X[?�¯N:�8��y:��?2�%��=�;�j��3��{�M��iȄDM��X4��&�o���cb���?�f�6�Yj*�q��/���O��ȶ��k>�A�Yg�Z�&�WGP��us��Ջ˄?�Ew�A���픣��#�ш�����*�u�&�>�v�����EiV�<�<2��e������gbP���3��U�2�_ߥkiL��|}��b&��xC�L�ɧj����"�G'_�i�&�"��������J6j߁��	 �����?�ЙO��6��ԟL$9��r6P]1��}8��?���W,�td���%�`Y}�#�h��[�{�3�s�����Ă�6YD�aa���/U'=7�"_��2_-g�����8�v| �2f�b���+�	oBޏD9d�ܳ��<�V��M�7Wů�3���Z�]����[��a�X�D�N��<oB�Fv�!8����^ݙ����-����u��ʎ<�	S�N��#[���v�6@��'uw�5?����Bg}��g�xNg�X��jv���k�s?{v?��$~c9�D��[�e@�oH��ډy����E����1���y�C�8���ކr�&m�*
̎^�z�J�]�&o�Ր1|���*�H+e2B� ��꥞6�s�s.�^�N�@n����G���J����Ȭ5J\ e��QX��}�6���wsУ�|��LX_��Y�W�AZO�|:���e��Ɍ�̀�u)`\w�����/(�p���>0���Y�� �a~BCV��Q*�y�Z\G �T{�D�n��0� l���7�ڃ8�n?N���
�ڄ$�G�����1f��1�����Ӹy��F�y���-Q���d�w�_sȼqM�|�>�� ��Kpc�^V�y�U�AX�F�i������Hr�l��N>
�������ʭ��D*��K��%1G���k�0��Q��^�g�%�E?E��;��zi����2�$��Yt����/e�곳ee�Hݧ��F�и��v���ۚ���*�:�0T˫�qd���g�s�D I�]��v~�2�<3lc+�7��r����a���[5��8I��35c�2t���^M�|{��ӖA������4w^����ݘ�՗�=�Ә���4�g�'�v�'�2���d ��|��S�U�r�c��mr��f�*������^C��c�)��ʋ=D�iN�g�fs�m�� Q����p{�[�.<݅%D��.����ɠ��p� ����g�;�6T�����(�EE�Ц���jqpC,����rk�|�;5�F��+�Fb�P{����ԟ��y��^�9݈o�vS���
�X����F)"&I}!;�xngX�J�ɜ� �d2��)��G:h�A|��Ж��"k,�M�9T�ѷw���ҷC����U��� ���C��
���k��Q�|��M�z\�C6\!��o+�ؚ�?`��s�aE�+��f8�i��x��i�j��J��͙�.�f%�d��	}�v��Ȥ��c]&5��G6vrÙ�X�a����!KL;ZSYM6�n���	�{�Pf*.��i��2�G�[W4�]{v���b�&��;ö����:\Qy{gY/�k],ѥ���v\�#�d�
v�6�Vn���`/i�Js���.�&g4ع�����:��G�S:���z����p�^̧�G��ܢ�(&}��0O��z�S�y��d7�.Y/�r�u�ZH�T)�1���]I�?�^~�m�\fN&��Mn��5(���O���m>�Z+AG)��G��4��E�&p�'���̃v=�I��Qz�O�;X��e}/5���n��&��[��L۰�~<����^P-(��	y�t�?��ԯ\/����9%�iR��lӝ�xX�9ˤa�|0�eم(RJh�
�k��A�Q�>�ol��u���yx�R���?��c�����7�l7BM(T0� �+M�vV�ovؐ�4�Qݙ ��k;Ȝ�2����.�)�)��7�������5%e�t,�;�~G�ϒ�B���j�M��5��RQt*9���8��~?�H����?��"��1�#�|�s��C��<�-�I�\x�k8�0�L�C%cOڳ�^?Sa����k�������$r��T^�U��'�i!�:ڷ$�ƙ���GY,!O����1	'#t����I��u�3Tx�~}��Q�OiR����&���𥼓9_J"�M�(�?tY�CR�������#��c�B�#!=�d][��7V�2���RQ�/|af>K��r2�ۯa�`�<ƿ��p*��.m�u�`5�������'wOB�����>ۍ�ۏN}Z�lEN����g�����~��z�k�P:̉�>�Kb�|�|I�9��O�,����D�fj���iD\���ٻ� �<}���bk}����J���6>C�v��ÃP!Pb��T�j7o�;�H{Ƨ�J��$���P`������:R���:��n����' �[8B9G�'������u��[��u�������}K�h6f�D�������"�qY�'>W����dl��˂RP��=���A�V߯hZ�*=4n'�]�Y�<����$x{�q;'"7�)��^�$���a�S���I�3R?1Hݝ)�H�
!���I	����g�ڗSXE}��ߧ��(�����opX�Jt���ʏ�S+��έJ\���k'�IX�s⌿��м�k����m,BM��Ұ�YS�2$��ô���B��,��ӔG�7RI��$�Y�1LH����G��̸8{gP�6US��sǣ�`� �546�m��z@Ԩ$�3��A�]ڠ���d�Ŕ6��T栢	6o��S�j�x��֎����^�3��Fb���MvG�Q�X������,G|����^s[��
����ܙ��B�$�����u�\�S/LE�d'���I�.Z^!�r-͛�����e��)����c�~q�|�H/N���5O�G�\,l|,���̷�z�F�����I4J��#��1C�9�)����]?���L7�.l�C_��'~�(�p���D������<�R} ���v�*BK}�Q��2Ud�iu�e�͵T����sͿa�߲3�o���!�/���p��(�rBWQU .#��D����p��^��2 W5���(�}T v�n�6]�M��h��Z���M+������.<�N_Yɵ7�,��X,�vq@.�m�p*��3���m-�MrA�����/��[3�5��T���m2�9�jX8nҬ䴗��.�\���W�� EPA��o��9к]�����)o�T��J��9����R_6�I�S��q�V��w0�t~8qHT�<�J�5��_y1�D��<@�Ye��W�D��I˽���k�dA�-��c�f��9�GG��Fg�ߙ��B2S]�;I5�d��+�]���rǻ�w��(����Q��/����d	q 9�+'�´'�p�-�o�0�����w��"�#ks}���/�5}�][���8;|�~�%��o�4�o=M�R�j	�FjK@'��v��#�u��N�*�F�O)2�:ǡS�wU+���aN���Mg�*$Г�s� )�������N���q����)�v�-����f�;S�!��Z�W��v)�ـX�>ҙgw��Gt�ǩ��V��%>����LOD' �nꀐ#��@��K78��U�Dɉ݀���A�`,}��dc��?(�z������Q�@�]x�P�)�T$�%��z��V;�x �i�\����k�IA&��չ;�+��
7c[�֧4jBK�����[$Bh�!R�	��G�%��+����r�ݸca�	�!J{* ��*�n5O��q��->)Qv3g�TS5�y�;pGL.�A��1�63�ŗ6<�-}�lk.�Ћ �[����.3�(��X��4n��7�PL���o�*����nK���Mg��a]0��8�_i�<��{��=�vM�t�.�'M��"�Vu�����2ֵP����&�b����t�E��1
Q��_N���^�_��Do��jG��ε�|���"gC�\ʇd��A�&�R�� �����:Q6�]�~�E�����]1&�Ƣ���;8@1�^<����vc X�	[Y������0�w������=��X zV`L���N�74��,TO{ąj�]y"����y���<TћȤ������Z���x�		���t{i��&6$�&�^���]堦�&;��h��L�FE����i���R�=6��-������ ��^ �2��N��2d�^��Ҩԣ�k�\ˈuꟚ�}IV�`dX�����v�@/��ù�cD����e'�{�yX:=�h(�Ŗ�f`#�/N��MZѝ�,�����B�GlQ`*��-��>b�dR�������$j��T�)�,2A�[��L��:�{����vZ<i�iZÕ<���u�ÕDOr�7�#�'ԟv�i�`��᥋�/��ofa���� ����#K�H㛡�-�W���V�C=�:Ͷ��mk�bg����@Yih��n����^~�ߛ�d� �W�U�w�\;���d>q0ɾb��x_�ߛhٴq̚x�؆������|�M�nK��2�?�ٹҠ�=:S_����P?�P&�D�z祽5J>Ɩ;k�G�D^�h���$q�hݠUk�Y�N�l%ɳ��F��h8��$��d1ZX\`�r�d���D\F*�1����Ehc���'.9&;�U}�	.X?�??�oګR�f����)�ˆ{�%�`�q�̂����紛�Pҧ �O�a	,g�GR�����I>�p��k5�7
�z����`�v�o]�;U�E^r GxB6QQ����M��p �L��!vU]�o>�HE��];qo�F�3r�ctpV��U|@R�ml-�iq�F+'%��%�M&C==��oN7￀u�Z�PԄ�Gm�4�N"���/��:���ÇJ�%� �~��!ۮ�!�Mྻ4~y�9q���.0���l��j� �+]΁�"B�)�u�*��Og=
~-���$�u��퀎��m'�w�˞/�.v��c�8F兞�|t� G��r���Uh}-k|����%k�*nJ+"�y�M�S�6��~sڧkF�o��Q ��[�eB��$E�P��\�O0���('i �ʊ�?���n���F�;��T� �$�Xߐc�5�
\�U�sr���?�T򞎫�E��Ms���o͊+���4�̡�{�Hh�bP�,�*�#�"vGC.� �̭zX,�^��O�>|Й�V�p��T�z���bYE�G�e�WUoս��M���2�ɥ�!P�c���{�O�1w	���Pv2+�T(��4���l��'Ht���"�����DN��1���P�"Յzܸ�C[i��H��=�<�h?�!F�s+F�#E���d���T�z��ƶpƯ�$V�ݠ�`\���;�'��q��}�'���F:������K5���G�Õ�zW���Ǥh(q]��b���y� S��M٫�/��ɟ5A�R>���k�Q�����%{mאSL��Z���Um��ؠ���Gy�*��0�����}s�A��H5z�?\Ɍ�k<�r�P�'ǽ,Q�����kS�<��Q�2��Y�S��cmҁ��JQ�:���ӥ$%ƒK/�I��A��<=0���%� mP��Ii��|R��ס*t]p��`���m���2�Lس�=��c� �.ԶH�bk)�]�x'ﺣ#K$��u�y�>�������j@KJ��n�W�w'�-��'3{�ؚ��&=R��A�%�J*Z~��@��oz6�^|5N?$���������Z�N��.��ܢK�B|Ģ�J�9�1�������+^!���<��]u�^f݄�����FUe��ԋFm�
� �w�y�ʘ�S(����y]N��4����:��'��~�j�`�����I�/Y�Hjُ�g�Q�%'�w_�)�?a<|��;��&v��X��!�W�8%+���3�����$�vpkaO�)Q���Y���R`�Ovx�~�(��v�q���}Ӄ�8�O$�8�K<>II$w��v�=�eR�R����jF���
X0j�����%�71����c$2�4�BFl� L��W`X�h�A�����e�n���YI����˺��l�E��c��QK�pH�0��,��^�����ڬ��J��TiU�n9�H�8������cnpDZ���B�>� �G"(��9� �p�0�N�����y���m���J^i�Y�����He�"r�����V��9C��Ԙ:�T�9�@� "كٕW���C�x_��No�/�J�D�w/��z�0���|��#O�yվI|ɋ1o�Bx �Sd~��e7@Ϙ��!�C��//g\h��7s5c\�����c�2��_��	<o�	�k��5L��5����˿�&7�a�07�I�B�۴';�gz��KQ�J�YI��%p��U���[*����@6��f$�xyzǂ����pW��=(�N�PYW��MR�T�z�q��	h?��V�E�!Y�?���������f���2fe7��|dv �n�5bpBh��f���3k�#�IC��ʻ�ݐ��\ݠ	%ԍ��G��s��a�D�jmaE2M�7��h�s\%{Bv���.��!Q�Vs�
�D-��a���9�ně<'�S��;�[7	�d��n� a�7I�k2�O�� Y��p�7\�����o<R�.An�K��̄�X�[��Aj"dr�N�=���n�$S�e;�
0ݏOCys{�{)@]�J������x�
z���+$��.b,�'/�t@��RG��PU�Aܹ8��.��Ԯ�{q�#�E��B��j�<*Z(���tր��b�i�u��H��Ot�t`k��SQ�o�3�l6؂�nB�����s��(J[n�h�w"jgi�{<iG��v2��>dW��oy�\�W}1���BU��w��a�H<D~Ӏe� u��K�X_�(q�OI�<��-oޚ~L��[�4���_�y���e0���@?͆��p$�<l��P�F��L���R:kV�(?�HaE�q{V�չ��9�L���FD�a/ޅ�)ľ�!��zY�D|��n�͟�jSg	���b�l������j�0	ۮx�*�]�b>��ȁ�s� %;��_�Ji�t/;d��xٶ�,��φbudpM���}�����w�*�@����gce��(�A:b�*spo_*� )
��)AI�K��vl@��f܇�"��5�媇;�6}7��E��W����f��l�3��f�F�.o�ތ�d}|""����) ���'ɡJ�L9���fv�@6���}Sa�_O%�R8���a��_�bQ�h�@�<����g6�G��[8����f��2I�I)�Q7a��ΆS��q�JS��]S��h����hi��q��I�~4�����O?�
��7F�����o/c��5q��E����h�Rc��FH�q�^���]���%�~қ�c�_���}������87��őݯ�L EI�ӥ󣉙X3��t ^��*�Z��A&�0�����܊g��%(��ɔ��׃����z]�Z�g���C[[��8��w.�4�	:+\,�AZR<k`y=���K�B���v�k�h�|!-fq?���{�~d�2�慿xu�7�ƈ� �m���E~?�/mj��	��FF����Dr���6�D�>5A�߯yx3)C�EG�z���'໡�:4���,�3��S[{j��$~���{b|e=vR�S-�/�D_ 7u}�A�����:jJ�N1mA�F\z�L5��-A�:�d
%���_�sܐ��-�8q���*A�6���I��Qd$������\_L���땫;���~�YklP�h�C)l�͸r�DY���󐷵�.�g��M^�ֵ�~�Ż��.�Ԇ��W�R6,�窘��6#>%�`�����\�W�L@?����\x�)ץ��y}>JE`�eZ
�-�y�H۱�f&��/Bu�%���e���?f���|��&Ȗ���lt�{��|�8��aө�
n�chM�P4s��h�-���5O��#&; :�.{����m\� ��ց�+ �Y��G�N�3�Z��ߕ	����o�f�nF@�o��Zŭ�O>��ek�����ߺyi���#�v��`Y0�w��ȑ���c���xL��(�Є�8]��&BR=�뛍uD)�t��@���;}��f͉�o�����ڍz��Œ��p��0�F�j4�B�����Dˋ�u��k�μP���kI���Nk������ s0��]C��A]����JǝR�]����+�M�M¡i��v͒����i�R �k��l�W��I�Z��m.K��g��q3IF�-J���5���ͭ:��J�Xaڨ�[�GN���{y�����U+�woV��*�)׈���W	��5kﶬ?g�_~� �,�v�@k�밻?��"�����쫮�,����6�٥���z6�
�i���w�/�c{���Q^ ��W(��i1�#�T�B�$L~h��2n�r��a�vV��D9I���x5�ҺǶ%
Ry�puop�g��R��Izt�dzR��齊k�4슠�/��6�x���"�3Ƞ��Ic���|&��}�(�4}��qz4�
_Fa�D�nc��	W&��Ȫ�ݾh;EVpg�6&w�:�gOa	p>)���-}c�d���`kW��L�D�j9�kfx˯����N��l�f�Nذ��`����9������q|#��Jސ(��	�?��K��>O�c���AH�r�|E��i��&���5�1>a����7<�/ӄ�ػ'%��D�J�H���$��;b]���2|ON*i��5���<���(K!�#;�	���﷏~�/�)[�{�2�l��',T���9�r����e4�1��mX�r� Ω\���K9\ug����� ��*
NuӐj��fR��@F)�`9=ܜ,��n�A&^��gqz�4����#���ؓ�6&�۸����h �wѬ�v��Cٝe�t2�E-���#�x~�脹L�U>��Z�Z��# }\�j�A�ng0P�;,b�Q�3��K�#��܊�M�/̿�S1t��� �I������.oZ2����߬W�X������-~+���+�ť�y�1��P�\y/&%E�[�9}�v���p��F�>�ٺ���NF��y����: ��"�~Rt"�Ikǽ�P���<��?����j�v���D�!?
�Aٯ���A��
H)�1!����\���h�Fԋ��w[�w9���}�son$�z֗W�m1�Pȱ�����]�؇������w9����崧�`kr�yf2��B��N�:�k�LNgsY305>{е��-�u
�Y�$R�E�$5F���Q��"C�w�����O*��e,��RZ=	φ!	�ˑ4a�׾�
���`����wh����@�@@�΋;Y��-�f������<�ڵ������ܗ9�z;13�p;S��2ރ�7�i��E>��C����NqL�s�®w��&h��A�4ί!$�]��$.q؄_��>8�ͺ8<�z�u��E��Y�*��J�4H��h�`�ߚG �m�@=ϜeaF��)�9�7B_2'��T���=ũ%��~"$X�tL�P�];�{{ܙ�9�݌ۙ��� ��|"&M��)	��TQ���o�������.�졂�����-Ο�`�T����0b�B�*�̣�~_Jc��3���a���yP#����l�,@P}�r�f�26ep�I�3�;��y*k���UbC)�:ĠB�'�?�-���L�+�i�Wɍ�;eTʚ Y�-]vl���^�NT$�&��9ྩ�FO����5f��yo��.F ������:'�s��Fu�"mc�E���t��|��
9�:�H=ݪՎ�JP�t�&�R���"�s+��"�d�I����g�S��d���g�x�۷��%��伆���B~��!�jxV<��.I�򴁙�vj+�ٲ1Y� �P�x��3��	������	��Je���X�*�������h�3x9���z�r��l
a*9	{~��ٺ�#���z W��8���s�rv�6;�kG����� j=O�f �����H�"��̈[�.G���'���o|B
�`׾Y}�W��{�IPy?1�@���.�v��b8ԋ���w��1��s��ji@ �쯖����3w]�!r$����Rc��R����h��Y���+mՂh�b_2�3Mt��ܳ<�'Y>��vR��E��4D�M��gGR��<�J=ξ1�jo�����e��`��ݪ��m}�����
&�uKX��I���V���\j�\����;%����1���j@F9�,�Y*��V�Y�l�0ba�����ͯ�¹
�k�mI�Wi}7]���1a����e�l���x�����<�s�R�4�}��o�r��6�j5?�jZ��������<���b�� �G��娲8&N���i%�>/��%t��^��~��B̪�e:8��'����p�R�W��~V�ka��\i9��r��s�	t�I��{��}����Ť����� @����](j�c�P����������V�7�H8��b�����<f��+���M�E����yZ�E�l{�� ˑ�_-�-���jV��x��a��Kx�)7�ƫv0%~�%�=7l���/䚋�/���\'j�s4*�,cq��>��"��j�����&c�3�*�~NJ�֝ֆV]���EA�$���2Z�iͅ|��v@�:�f;�A�<��"�x>]���/���BsB��LsE��Wr�(�<���\��QE�E`7�8Z��ҹ���W��)�n̥F���4>Z�_�2�z, �7�Δ�!����U�(�~g�@��[�)
�L��������q|TN1�s���"gS%�=M�0I���'�iީ���6%F�p���J
�ͽ���tm�w<��K�'��^_	����؊���ܟ�О�$�E�S�'���ߧv
x�5F��@6o�Ekc�]�&<>j\���F6~,��-�?7�6�C�3�bxf8������w�!�j�s�X��!>���ܶ8KS�7�j4�7]Ӿ��]=z5Әw�L?���`��R���f.;��i{v:6�TH���
��j�a�>�t;2;��El��&u�J5�8�9��SJ��{�e�r�(;;`���F2��-�����
�A�OEW�+��kǀ\�ϫnF���N<���f���5��f�p�.�C���D�վ�C��N�Q�<�_\눸xէ�k~KT����;�{C�>�u8B�)���aP1�9����{{��u��-�<�� .kMЭs�N���x�'�˞���C�x�u��baj��� �Q5n�\hUn�^�e�����$
T�L�sj��s���H���)\��A[��|��[@��[�0�qЮ$o(�r�����/[��R�pK^�;���jS�` 7s7[� �I�Bʵ�4�Y�B�"a��}���-=º�~��l�}�/&\=�gL��?|��-4@�W���5=k����L)t�g8�b��g��?+p��Qy���g�>x>�9i���$VmaJ��/v�T�l.���i[�PS�4��d����W3�йga��>�ܹ<����P�q�Z�9C�G5�l.�V.(mw�]�ۭ/ߥ�V��O|����,��~��!��U�H��Ӻو�J��<�F��W��H��I$��e�A!�Z�H���-�%� �r�W1e�W�*�$αkL�|�&O��c`+D��Q�s�k��%a�� w���V6��r��l���Eٟ��27�p���=�#�'ȾM��f�����L�~�	�m�7 �/lIls���/@J5'ç��p�%ی��l2`A���`�ct=x]<�R�GK
��xA���:!r�=i��ؑ%"
EmZ;��~�,*��Zͱ��8���f<5�!���A�ha��+>���ET
*��,��%` < L	��:��wbd�b����Ќ)�6E}` ���)g� q�k����f��"慜ʶ�T��A���b0 ��B63��ֳ;�]�� �2��_3 ��M��~J�����^EW�ϭ=x}����B�Q��/8��7!i���M�	0
4�e�8Z�[������C���Й��6yW4�*�Ó��@�Y�0�J��},�&��|Ŝ�9M��ǧ�RN��p�l�}oBOUr2'��ܽ�x�h;l%X�~yQ���s�v,��|��ZĂ��rj��U���x|���gQ,(��n"��F�����z�uXF��ף��D�3�;�Y<��o����k
�m;�pr.��� 9і���#�ȇ
�>{1S?�$�.AZ�ŖgW��H`uExH����3q(��|N/�n��wX}����)9��8�vE~{B<���R�׆�7�ͪMY�ݗ��.¥�p�_VX��kiq����=��r�ff�,IN��-D�u�������%+"ybi��YZ��Z[������i�kfx�44^mËD���%�^���{ɲ,,'�u+yv���:@����S��a-+��^$&�nݘ�A�Zv�H�1�5�M)�9](���YN�I%�L�d�
J�7wi�_�,Ho�|h��K��z�֕ �w	y7e�u*Z��2�g͊�p�4"��گ�I���ۨD���^=�8�������,�a�WkN��j"فb�5̈�ձ�D�ޙ΅��H��'A���O�(Z⼾�U�~"$�4-����w�;i�2�~_���SbXt�׺�e��1�*��Gt��1k~���l@������}����$xq=������Q3��Ü��>����3�)�-����|�$ӈ�S����fm��^�W�VQO�z\��1I̖�m�!v�R�L-`�IXGn�g�ט��, X�W]������AcfC�3�j��[i)��,>�I��5�s$�L���J��"˻c�:���x�- ^R�$�U���t�Hp�Q�y3S�
�A6&A�#70�t].H��ߙO%P"r�KB�+8�|.M���AF�"�m�SC�Cڱ;�v՗p��( �\�h��'\oP0����`���׉�rAQ�ƽ^?R0KK���C���������#�6�gh�n37�XS����|G�CȞ,4��E�����^K�x��R��<Fz �#=��3�~c. M��W���@��lp��N�"���`����eX�+l�_$��ߑ�O�2E�Z�0��[�A�~`1/��R,X��0�V����g2W5���Su��1�^���N���.^v/�.�UR)��RfHtjChθ��J�-xH�Ta�$t���������iNg6l�pj1�X0�i�r5B�.M�m��mWQv����h6'�d���4��q�Q1�Nɾ��6&�=��a37Xһ�ך ��5����T��X��F|O���p�;��k���(^:��4��5G�H�H����d*��i�I`3��WV��-�Ƣ�*��_4�?���Z�]e�}���|�n=��П,y�������ޖ��Wz��ҙ�G+>��!UU��QȦ%K"b&z4�Z9y�� ։�oD�﵉I����8P�f{oM��;=f;�)Ҝgh�2�uj�؃�q,���ɝY���I��O�4a��>��쓥�8�D���H��X9���d_Fj�F�t�X����W��<��^�b+��{�[�;k�|XJ�eO��!�|���,�����m��V�s�S~�`��cs�ůk�͝�GcO�Ak�-�1����ͦ<Jp-Mk����-�	��2���t]��!������P
*��I�3Mg�qx蠸M�}�l��Cc���c -4\.��Q[��Y������j�2q�YX��5O��8؝�I��/1�y~���_G\v���&SO�s�GiY�o�pjwv�KM�nL\�K-e}��=OǪ��|��6��8X�*�����K�-*�חi�{�r_sD���>�����ADFT�H���g��R*~!K�O5�T8��En�v*2�+���\����ˎ��d���J`ݎ yu`��YNg���y[c�L��%���g�m�@Y4�	/|׉iG|�
Y�]/��7��K��w.����'��ү�>��}f����/�U��	���`���v��)<�	�~�^`)8�YMr'���y�Q�5/*���Q,�DH�x�MG�-3d����.,���taVL�3��	[��>bzֺ���V��c�ƵӰ��1���{�RIs� �Z����r r<�1���х�Ţ^@4/�5V�[���
ƻ,V�$>�6�;H�
8�i3�зSd�L��d�˙�$�䮰kv{#�d�*6����@���b[�inc%�T��	L��SG���&ט���h]����<=c��s����^�x�ѧ=rP�2�D8�J=�'F���}Y�蒴#�I��$.xָ�_�|�E��sX��yd��Y�;0ՉsF#q������஄�z�a�kB�֥�B����_�)�f�~txN^B� 6�Z 9���N���L8M�Α9��F��u:� ��E�r��)�+q�u��1��	'�cP���*��J�8Ԃ�WE2�nc�*Z�Pm 8O�����b6���h��~�	�*Wn�<� Mu��]W�8��ƺ����SҜ�^i�f��ZP��D�*�'x�.�F�!�l�
�]%ʲ��=��ĺA��^6�q�A������o3����@�W��L�wo���v\bH&T�Z`��(z�>�]�R��G�*�i��X��+?���_l�E�ݚG�ݞ���^���$\I�(����纅�#����A!ۜNY f�$K{�B�~��_(�>C�"Ѫ�7����*!{S�#/�BJ�G[�f�뻳ZT�N�r���xrR6�he��)X��@�.Z8
�"p~�ˋ��Xa��t�;�s��Tq3CsY[���.t{�Su	����o�K*�%�V��o]�ܜ��,a��k�~����n4���dI��?�5���Rh��~'������W�\q��nV�ɝЎL��b\��W����_��eǝ��Q�n��z~�ތ�}��%���F7W��w�-bZ؆�"�Q�y�3�7�o������Ǻ��<>R�`))�C}���~�#�m�}�v_n�(�'�i*���93���}5���X��2*�.����HY���¹�G��'�%yGoV´J���Fa}:I���b���y�+n�i��(c�6z|N�U.��^}��L)�+ ?���K��^	��ܥs{@�hz=*��F��P�޵�m��Lj��n��̆�}i��)F����p��t��Xu&h��G��̓�V3{���'�r9��8�`$�������=?����D�GV�6��vAE��I�4�Y��E|q���c��b�+!{�DӸ�8�
V�o�a�P)؉Mw
֬���G�C�x�dD��qR�b�!�%�t��^�_�P�C.ȋ�Ϣv��T�)�l��k�O�Sd�2g�Hx��rI�cCb���=Ӎo�k_|��q��,&���Ȓ����D�j�]�?��j�����C�X�p=ϣ%�K~O�m��nB�?��h���.&u�%�u#�p��6��K�jM�K��J���u�t߬.�ܘ�H+��٘~-m-�;O�?R^l?n�,���/F��(Y��/iֹ�C|�EЭ�L����]��"��xV�#=4� 0�rD�휗�a�b�����z&9�*C�9�|��VC�l*����8��r.�t�S6D��Hwo�w�3���2N� �~��V���)�����#O4�_�B��f
�oѦAwkWW���}2�#���b�Z�<$ۼ拻�P3v��e6�Q=�]g�Ks��f&:T�H����J_�P
9]��I1F�U&[F/����W�m�������aQ�'�t���To>E��yѰW'%�¦U���F��u¥������ݼQ���[�����M���[�.rzN9�����ü�-ϡs�F�N�<��gs,�Arχs��e"��b%�1��ڙ~Of:����#��(�=��%��N�F��*���d����.Qp-Ø�$�WֽD���DPu��,u2�7��eJ�H����A�Q�rp�!��a��.�!8�k@0Ǘ�~e�n��|����5�����������cV��d��
�5"Z�R�;������J.fJ��"1kY%h�5'o0�Χ��M���B�Ã
Lq� C�t%��9fd4@���rc��:J-���-2��"[]�4�J��8��³	�}R��K�U�~��
���%�T�v˞-l9��D�Ĺ ��ŢN�kR!Y��#�RIe"�3�c���i`�݋�	R-Bk)ɳw��c'AF�)Q����c�_���=��7Ԇ��W �^8Z"1��m6�^�z�Ӹ.�&���D�n�]�:��&.e^�'�QsIV'�]��>/�?������e��PL�}A=�ۄ��nH��<����I���i�yU/m��?^
����q�?��kӖ��q����.���Uf��NЌ7R�10����j}~WK,M��pYOڵ�����ٯr�%2h%��S-�TBҍ݁P��0$I���T��4�N��
|z}�����E�)��(Yg��uy���Oڹ�%=�㋓$J����wbs�����I�$��Vo	��?�r�ұ�}�o��yDQ�J�u'kp~�!2���S����g�	����C\E�z�+�M�_Ek��x���j��67E$�+QY��lBdFE�K`]�����~�`���|ܤ]K������uy�D�!�Z�UKA����?�4�tG})�̣p��3s$7D��bI�x��J�U��~�+�?�
 �uwC�
��d���(�Ϣ���[��'������%eƲ�d�3"K�^�WT[��ч���z���ol��D�tp�NJ���v�uUg�AJ�ȑ�@�����PTDc2qp�[:(�S"f�@]ɿ�sRGD�q��Ś��Z����W�9%R�w�ǎ�<}�Z�j���^)q�H����<�3~�FVwy����KDf,
C ��~U6�ȂDFS\W�`�,�̦�PG�w������UR�%Q�q]'7�-�Y���c;]L��,\�Ґ�FY��r���T����zZK�L��&e�k��S�y��:>���͈�ȿ+������O�.`F5m\�$�x-r5����Xh�|4A�f��Lz�,m]�|A��������������:��18�������T��@v����ժX���ҜMRD'w!�K�rQ>�3�������t���~=�����sVe�6�O����RRN�]Ȁ)���v����7Cٛ��+�+��=��'c)'�5n��S!���t�J<gXk�ǴNs#�&ҝR��]�����5'qP9��Gi񌠌k�d���s�L������4ja�Ì1�uP4���-�l�Y��T��"�d�.'��RZqX�α"(:Dk	Ͳ,@�%^�Q���7�cӶ�� -�O�\��r;�?��r��R�R����x�	�Z(�+�Ǿ�b+�eU�8��y1�]�= �`!|��v���C{�3��:�6	
$f���t�>֟f�`����Hg;������]�����9L�mh���g_H��G�����K�^��@����F�_���7[vm��H{5SZ&��%ke��Լ�O�G]F��GD_���#{G�p2u늫��US��w���⁘{˼8z�w��}�rwi!�xJl���"�Z�m`;�.pʯ��Ɉ���=&�[��*,v����:TId6�M��D
��_~�T젚�嚣>����u�{�P�im�$	όǺ������K2���	&<u>� ��X���	��c=PL85���PlyШ��I޵��p|5KV�rq8�+����E�X��
��T���w:�;\��j�(\w��}�`�\�=!i�0͸Kf�}3)޼�ʁ.�5�d?��&�GRD�#����ʑ�p���4���t�aTJ���v�����Up-2$��n[E`�	������C%��y��ϳLX�a�9�AT:B���%B��L]y�<�_�{<GM�Լ�Ic�����]%�:@fr��^�"���*HJ�Xr?���RV�+����#�Ac^�Z�e��<eS�I,,m��k����C����DWF/�����OcP�4r��������nc��2,�}l#�2�� Q�@?��ś��@%"0 �� ���q`�Ji��a	���*���3LZDb��b�'IPq�-S��n��	R�*f&�&w$S�ő.����u1�^Jm"��w��=��	��|�ؼ����G6>O�}0�반�MTa������j8��]U,j(j5�����Ȕ�Ӗ����d����?�ML�l��x����(�M�$�x��M��#2�D�'��!n�����
133�����w?s�u�`��J�+z��ջ���؏�y���U�x��V����ٖ�q[\��������5y:xy9`ց�2�8HՐ��d�/dj@.�����*i��!K�7q�_��͂���q���m!��\�Ðo>lSvl��V�Ýc�f[��3��aSc��|* ��T�)w_a���)��&S�Z�a���r���������^����c�� ��ϑe���m(ֲo�(M�b�/M?���e!eH��
`�v��h`J�o==�����c��Oq_�"�����b�y5}VӃIۦ4�F�CN���,��3�peǙ��#fr��x���(��vLo��F��4����-�Swq�iд���9�R�v�R�k��]�yC����k����@Y�P��s�+�G)�!����f8��(�Kru^�zH}O9ц�b��P�}ӬO�1�I��V�[�����H�c ��?��gU�y�g֗�H8�{@����x^ib�.|\2Uc�[V�8�#�U��Ҍ�N��,�|�Ќ]87���*9Jmz�J���u[S���ք�s}r����o�V�1?{���C-ŀ��c���Ń�*��,��q�6���1�!6��VS��D##�
�T��/r-ցh���3 �I4���\@�je5_"c>�9�eyj��8��������`���:�da��0hcQo��P�Zq�d���4{���pxW�����hK�GyK|�iE3qLJB6̰�i���ɳ�$X�q�k������W*-tn�p���^�
1�:#ڵ8gpqPjԇ ��>����b�%�/Q�Pe�ㇿ�?��Y�&�C*Ɗ�ן��:��b�h�ߦ�����pRo����O��s�ݱxň�j~���cd-)�~�L%g����'����!�lM���3ā�� �{�~��F�c��HM�'6z;�C�eK*u��^4�8��>�����j\����;+Hen�Y'-r]��|��bJ��5��&�E)���P��M�N�������wG"�uL����C���ŗ�/Hj�~#��i���9C�?�w&�D�2���V����׭'�\t,<��E3��h�tn��e(`ܹQJ}k�<�5������+���ln0&�]�kZ7�UX�J�%��0�#����!���;c���e�F3Ċ�o��=
�[��9�I�0�����=��KG	2/��ٴ+�� ���Y�ȱ�+��v��P��j�쟨�3M�`	QW��{�l{rr:��'�Ѷ9j�$���\��T&�h�S��R�ʣY�r���;��e�cGm�)�//F��8|�G�u��h�ҁ�	�\�z����9fdT$�@�����G2���%����$0Hjp��dk�|����0r�?�#M�_p�m6B�)�A��yC�Y�YO��MM@lu}�);Ӥ{���<}�K�@��Ac�I���u�ҩ-�6�7���[��q7�ŏ�r�5~Ϩ8Um�Y���a�z�/�5���)���M�#�rwH��5���._wʼ�.`�Ъ0Njo7�`��|�=���(��q��J0�ʈ��>�wnQ�&�����|���k���e�#99�9���~�E���q{h�~&��sgw�9����(������������,ȅ��Ȭp�J��$l�گ�7Q�A��
C��Z�QK�^�nR���e���$�<�?b�����p���{�][�5I��(���(��q�6�R �;�_��:$\N�:�]�G�(Q�E	z~R�忘�����E]��ڋg��U+�~�x;�-:�������Ä��EY������1X�� ��^M��ş�K%��ha�d2f����Ģ�`쏖��O�O7]�N��Yg/n��z.�K<䅇��ŶK��T���䲩$��-���9��Ĩ�/����	O��ۼn��B\��O����hMT�����Gw�su��*ᯚ8lqd%�E�+�n4�ebq#�x�Ћ��\�a!��~H����m�C����"6S�BK�ƧH�V?	\�d��cTHPV�+aFܧ���E}<kE���<-&$�"M=~K%����!����������(`���ƾ�d���X�C�{=:s�Ľ�Ԛ&e.E2�I<B�o��*�<��p_I��]p�s��������)�V��g٠�:�qW[�q�㉗�2�o����l �"�SR���]��V:�s��G,��Y��<�;������j��,�߄��φ8��5��������|v�z��k^*�ܰIT�����,F=��^�>=h�*xZK�~C<c���~�Yz|��T��"�&
��xS��"����m�x-T0$n:/������P�!7�Ax��g1�!�@ l-�6���-���_]>n����+C�p,���$�<Y�U��Mo���S�%�W�_)�_�����97����kX[���[���(� Y�_��f������@�G�B�?��s�9�P����r����:����걿X$��V^���kӑ��$��)}hy.d?�-���e)ŷ,&����U��#|�d�ѱG\��������L�a6oa�w�5��1�{Y��B.�}�]���q������g�������l8H������x0�{
�a�ԗ�����|>wJ�4���ǫ��V�W��w���_U�6�a�(/!D:G厹�BHG�oBI��%7E6;=�D�(?�%
g�w�³F;2E(D�|tձ&k�x�q�1~����4Լ�w�w����;�n?T��\)�Տn����!W0�>/���r�jqU9mA`J���;V1)}��*��AƘa��S@�A�B��JB?"@;v�@xZ��ͧ��,��e�*"I�_�-�9����T�K5�D���;Tm�Y_lƀ��nO���q���8��<��[3��3�)��;�%qW�� �V��$��$m�� 욈���KE�k�O�� p���1�s�۽���t�/rݻ$&��.;��;�$?��Z<�~������N��_��o����&VtS�*���r���m%,Ncmeih��`�����sˍi� ���է���.P��}%���v?ek����9;2�B�fe��{��N�Yg��>6�)q�0�"'�`b�s�A�G�ݨ���j�P�w��ռv��\�|�խx�J�=p��upp�r'���$j���J��9Ex{��c ���`)y$�C�/���Ot����Э�B���K���y�)�")�G�?x��Y(�c" ����&�����g�b�
[>�iV;�nQ�͐�v�-��>��(����Z`8��yK���N\�V`��d�qħ�J���$d| �UWƸ>��v� Z	����=(J��.�Xt�Ԕ�C���^�x�|���T��(��������9�݈�q;PjN�[���O��f�ʂ���mK�{�"��I��֘b�j��T��D���)��n��g�#inx�5d��K�GثB���#�GC���`'�8E6 �֙<uM�Ä�k��`���&�8m�²�s��po3e���uyj��_;ͧ�.~�`˪�Zߚf�)\֣B&��;�c7�u88�y��󔑯L����>H�'�>u� �8����0OM���h{�'<��bχ�0Q&���s��Q�i�"��ȸ���c�9rRb��N��E��Ntʌ��7�����S��sH��O�"�7��+!&i���{��/�dD�3�t��,3^�P>�,�8��F-5�൹�Z�: N�Dѧ��k�my��G,��1y-�5V� \�!GB��O(�L���EpBWY�h�;S* @�S�;���o�g~2���w
�OUi�:�X�>�:a�r{M��Y����,::6�XW�o���o�C�^j�]�b�HN�=�VكQ4�&#9�5u����v�L:�LT�d�r>Iy�;Ƕ�� �u~p?�5��2)Z��B�7�(jEq��)w���y���7&&��:.d����iz�o�VDr~P�μ��%J�����6{���/����߹����7-CF�Q��ℑ%^�8�]͑g������ ������M�[Ǘ<|B�}!q�Ĳ�����ԗd�Ϫw��巅�<q�$$�/�<A�8�"�+�W������C�T�|E7�\�Lo�`�yQ���EjL���źb�׶�	��PCf���R��n��2�d���A��hy�̀p�F�{5�$�-�Y:� {�t�| 1����B����)c�H�-V���#o����/	��i�#����[)�Kk���t�d
à��Ȃ"ק���µ>���ڽz4�_�`

v �!�EUm��)����R?.�ނ^�pO ��_�:+镗�1��a>u2�>��*��_���|~pÃ��9v��7�:�^��w&��d*�-��&̈�D8��{�I>�yp~���캮��X����z���똃�D�f���VP��:� �J}yM���2<:��,�q�sz�TP|bi��<yQ4��Ԏ���к�:*[�f� _<ߛH�t8���PpGΗ���[�	��ͱ2���O[��"��׸c��o�Z�0�TUXKV�Fi����l@���g������]��H�I�g~`��Y}V�@Ӳ�BH��dA��� ���Z�4��I7K%q�iQ'-�F�daT�(��[jl	7�x���P;���,��nVC�J�Z�bv���ԛ���������n9�~�e��G!_�%�J��e��U �K�K��1�k�%s��õ�A�QH�Q��zE�ϲ֧ ��sa��O�-��0&��[6�"7�('
�삟@&��Zُ.��	������6dХY|��ſt����>�{�]D����WN+N��j��&V	[�h���I9��l��$���~P�H��VN�"��e���}�A��͊נeh�������5�ֹ-��^�p@@"���2�j8V9c�����Dz��3���T���H(�إǧd�5�	�;)��\U�@n��R��f�'>~�F}(�h�@��v/�T]P�4�ޣ�?^��<���U5&�a��.�� �H�<�}#�ʟ���iɊ��������&w0�z׆5:ɳ��.�t��|��9t<�!%����`���U=M�����'�3p��R��拈�d�S���1�,!g;�ᩩ�͚�Ƣ�� x�wLy`�Ƒkʯ̕?4�T��b����
������ݑL���MW�� u���u+�?;��-���r?�����z\�͋���M(uCm���YN��ԫ�'���糈>^�qʵ/,���lo��;�_	�; ]Q���/PT-��;Mv�)\yzRهl}a�A��z�յ��	'��e�p63���nXo�?�[��W�v�v����B��t�����-H�<w#0��7�V$�g�,__')l���Lx�cw�XA�h�{6!ޒ���,SSB������}��Bԗ�r��6�	Y��(�X��說�$�S�7=k1��3rLՐ����a�@�a}X�Ȁk�A�éS�ϴ�M���E��H��3qK� =`��%���9�~�{ ��U[�V������?d���s�aԓ�v.z?���}�b +}��Ívb$��U��x��0�8$�H��NMDd�ޒ��I�m���"vsn묞�a;�(�W{f��	J�Bրc�H}�,�j�c�i�m��WT!L��ρ�d�i�r��%|B\���Yr>��K.�0�i��IT�DnZlD#�%�b0��s�<�!I�JW� x�w~Bd�nS�ɻ�G˸���!��}W��N�|0�t�O�+�m�M-'��-�͵'f�.>=��[JS�)c�܂f�R�P�o.	=��� C�:m��"�|�T*��Al���6t�v]��e��Fk.���U5��ȟ�0�je�22��w�4��aG�S8�k�x�����m�N+����1/������+�ͼӾ$�s�=�� �WD4(1�H�l�����YtG��$k�Q����g��'�\�!`� �f+��2J-��<Q��}��t�HB�~5	5�*8��K5P��d6�oS�é��By9/^��3)���C,��Y���,�t���&�!�WBV Ⱥ&���C5D����i���W������`(�4�bVqa��E��G��/�ӽv��|&h�bT#O�$�0^a�Y"W�4oe\��ي����u���<'������v��H7�hu\2�H��Ц��g����Ct~A���$;�'��
zۋ�@33��Y�c�,;��:��T&��7UTGVd?� f�V4���͐�BloD��-�� t��Jz==^;�P�X/iL�-x�����k�8`S���| ��Re��"����,���_�����BTq�t��2PQ�D+Ue�TK������G�I��䪕� �$�ZMiܦ�.'Y*:�y�M�J��Y5/^2�Q��䉓Io1���;����+��K1�P��݇�q��~גk�_څ���
�%]D����V������H�����'q�U z��E�ZjF��\5=LuN`��MqP�EK~�-�+���+�m���M�0�����d�rb{�%Mr��>Ƹu�z9�|�|�F�L�e)�Ɛ���S��c�Oi>�c}�jw#t�0D�X��d��oW4RC��c]9�Ј 87^��=��0?09�������Η<$*�Ώn&��c���"F��X��6��a��'�&��9�Y/�m������n��Q�&^��j �pqoe��}��бcŵFO��1gW���A��T�	S�Ȇ�`�u�Q���o���䓘�CcY
���|�Q��ḸNWZ�&�+��������:�:����p��+�Av��J�et��_�wMa���-���@����w��~�&����!��)�ӛ�'o*�=Zv6��R�� ��9zl�����"N�L�¾�d;lWF�Ҿ��:3�P��'@I5�x�ZJd���~��粢X����Br��ڟҥ�>�Ƚi�L��SDóL"rs�%Y��q���W�L\��+��_� )��|0`�Wס�? ��:NLͥe��� ¶#G5ɴ�~�"�0Ryá
!��/+Ӝ�]�X*������	�Q2��Y��[��C�V���YD��/��xsX��ve5�k��Z���5���UIvBs<�Do���<))��+=T�7�t�?�<����;��eS�?v�x�}Ę
��i�[�3�RI��A������8Is�3�>+9��C�>q���rΊ���D�X�����rw�>F ��w�\9��5���阈���5dib�xW�<M������t�L���Y���~�vY��Kr2��˃H�P��]�?ժi�@m��
�ӵ�E���%	���m���a��Xg�*]��I�恛��`�u+{��Ap3�a����&Iz���Qgc�fgH)/�S9��,���!IYZ��*�٦�\����[ٛ8iA��c�����1?�'�W�[k��1��5��͝>�Ea	M��c���T���9��
�6e�L�������Y,�By̅�f�T�dY���j E�L�o	�)+c��������߀�Dz~<�B!ݓ���!��)�E�`���x��̻���6jO�F��@+^�"4�PCݗ��>�GC)���ʭwT،Ӡ��J�7+��C�5��zL�ԓ��`���]��ߠn���<������4��#22�kĿ��
/r�K���F&���ǃb�c���T �+�K�j��,��Y���t`g$��]�^b$%�F��J���Q�}y%�]���0Δ�p.��4��;p��d �8CbJ������?�0��� 4�������.��{.�;�?�����U�3�h��띰O�6ʵU���E� @	��D͔Bʜ�]�T�w� K��][e��2]�~�n�>�B^-�G֝Vς�8���bN��"I�(O���q�憬,�iU���䩭�K�߁fߎm�M�VŨxGc0n�d��-gM�f�{�>������H��"+���XT\���̕�*���Taf� �vN�bhQ�8��Oy������I'z�M��mpx�y�Qyj�ϥA�zJD�#cn�����П�]�����3�[yu�o��>%kS\=s�?�ߕ�#��?o�3�J~.>����2(��{��6m�
��~�D�t��N ���7�i{�`����i�o֖q#\�i��m¤��T%f����h���xy}��DA�$���
謖�b��6Fw9��j�?��|�E���rN��77.M�Ws�'��z�>m?��)�|���
�/��K{-������K�Ԓ��X�4��ڟ%h�i��dJK�k�p͐%T#ԁ7�o�a�I"��O�6V�\tAw�Sd~ޚ�WN
ސ��rӸ�h� �F q`eY��/�H�����������D�
�H�y���~���:<���Ի��t�)�_���ɟZt%��o��TO8_tdIuQ(k��d���R�+}��]�{l��xoJu���
���X��7?�\%="[�;O�*=p~HjC� ݊�}��N�mA`�;�������?e�M����&n�v�N%0d���)+s�o��Ӣ�?j�'�xv�I �ǳ��I�[�*��X��=Xi��Ck�3I�'��7FֺR�B�D����n��X�A�)�p�:���nDY���"�)]1����?kFՄ����X��8Y��'h����+ :'bE���f����
 �s��L!���
X��|{}haY�#��|����������k��ށ�W�/�V29J�];
��ғY�x6S��Bg���"����r����z�ٖJ۩�94�H�6qQf�^Y�ڝ�$2����X{|V�����5����ui/j�İ �;�t��kp�%R?$j�@X�h��t�4���fr��]��|�('�%0�3��f��<<p��h[��sQ��	uWA�*,���\4���q��&X�(,fNXh���HdBf�i6,��k\q�t^7��'b#���H�"�^Zq�(�ӗ�!պCH�<$?w@��ʻ�St3+UmU>o��v_Fټ�|�n5�?ެ]�/c0	PO�/��fIw!m	�EF�k}��RU˅�3��,=m|ss����؈���)��
�'mP��0���Iptx%��pv�D�u,�f�+:���]�P���7E �
h��\G�����`6�}�ArL�����\9�E������Y��Ѱ&Y�f��5���lʻ�>�ʠ^3)��w��I��;5�
�䇴�\��Y5�����P0[�S"����W���<Q���B�Mne�!z��ΐΤW����r��%�I+�iDY�&%�BIǤG'�i�z�ػ:v�*�iM�����|�K���B�8�̂�NS"��UDz���[<X�{�p�G|-�8��Ck��@)P�D4��NY��ȸ�I�h��X��c��p��q��6�B�n[U�L�UU�'z�D�f4��g���t����<>�@����3\���b�6;��>�K�_��)��h���di)+��O�|���a������.��>Hc=��B谱�5�-O����^��&%pv(�v+�tl���Q��U��N]�Kd>ŢV2܁�)��Do�X.��+���ys�������O�d�>�\����f~19)����.��WW���Аq��jw�#���Eꠃ��l����3�~ߴ�*���
j����Ui@G-��RO�XӲ�d�`z9'���'=�֪���W���w��kw��"Hw�.�݀�܀"D���!�*�$�Q�u��[1����d�%�������Ŏq�F�k���>q��,��g)�})�Ԅ��j�2=�4a=z2o+����',�M�U����Z�Z(��GL�_t��6�:M������ӛ�S�D��,w�#���	�D�7MG�22��GHl�~&��S��*��͂�nNw���-,b�	
�F�Ŧ��9V���P[���7�����I��ħV�6-���jQf0C���~t��z�,(�EQ�Z�x� ��Y��D�yJ�\��I�9���b��(Zb����,��B�H�F�ew����E�'渖�φ\�V%�Ŕ��0�+HR�#�!�O���: �ݑ�rn��Yv��/poqR�l9䔯�R^��u`������3���l�/ݘ^�,J�J� ����1��f4��(�1��Dk�Օ�3�|�(��S-p�.>P�0�e�g�>_ �e#��c"Q�2�+)��R3P��,��c�!��z#�ֽӬ\�
z0�����Q8B��0����u�?�3��
R�8���f0itP�Rx�h 2I��t,��n�oL�VԺ�+Z��R9��ً�.��SP��R�Ѵ�H���� LO�U�l���GTS�}�4�:Sx'���g1?f�� �ӿv�p���X����,������A��un#4PW+��J;=�E*T|��������{�8@��;�O��������x�<o7�f���.=f���l��p:�ؠ�q��I^St�*�I�����	u�d��W�<<��i��u��?�lPzf�gǊq��n6F�$:��x)"K�l(�xxb8�2�A6$8R3a���Pq�S U�|	�6��"&��)��5���3����u�]�p����x�0!�u�ab�T ���-����	E�h���qG[TͿ4ǰj"1���55Œ2B�^�-RB�Q)��G��gֲ'(����#Hj�^�;0���������8]-�-M>�q[�bB9��5=wa%�q����e��zq��[Ip##�]�;_]�,�_��';珴����b8͊ˌ'���T�dW��4?(2u�}����2XX�δ2�y��PNR/� S�k��e����ep��Y3ȃ;C�F0-tZ�s�vW�,�H�Xd�'�AS�
�=��3w���jKePɕ|�Q|옸EO;�M+a���0P���1��� �-� ��](�o|��BM�璘v�����NL�Ýb�F'�o�h%�r׶���$ErK�3��dy�w�Ғ�������UE�9w�䅯��iʺ~t��#b�w�'FJ��
a�`KWѷ�E،&r�_�,?:t���ě}N#r����J~R����V��Yr�̙R��-$MV�י�T��K���t6O�ϯq!\��j�!���]�6R،�.��YH��ڵ��@��YPi�Q��A�A�7/dA+���������;�7K���` bЪR�� $؞�|��"�?j_^!u2��IEj!!t�(DqhE���^1��Z�;�jGֱ���}�i�Q��/	���e)%�5��2�諽�"��ˎN{ �ד�kw�-��p�#g����c�n��ѝ���1�Ӂw\�?����?z���vz�gZ�t�^��]�g{��X6��T�0�P��LV�-���n�=�R��q�<�ʿ�����n�e�]��U�m(C�J��Ls�c�ڻ,|G.���8^� 3�ݯ�S��ÆO��e��H��e��P�1�|�?��c�kZk�J�49�I�
m��x:΁G�m�u�|$w�D9�	.ZɒY/u�ӈq�$R?��}�?:��=����c��!T�k[�1��Z_�f�^��T�p����w��1�����P��_4<<"?7��dY��z|�B�壬g�J��K�ɘ���$/����2�<s�c*�����m*��b$�,q��>�5x���:�P��Q�L�$�:����J��ɞ�(��?z��<ÆH`��q\�c����G%�GpP���1�L��r�`D@��1���}k�x}�̺��\k:��׋�`�w�$�K�;5.�O��ؑ�8�>Ǆ�"�2��G)��T�u�����z��@|��U�4+�j�z s`m<%U$�V���B�+Z�����o���E��I���*˫�禪x���X�M�ZK����_�QO�頻���,O�sQ���_����d�
p��~'��uC�x[��I��lt�Qף��ҽ�ϝdڷ���g�ג� bj��L��>����0|��>�����"˅}�f'J��'͈��^��p�����l�m��2..Q���OϬ0�k
�{h�t���N�^Tw�L� ���c�~��El��#�)��#7[z��@͔6����0|���]f�j��+ӈ�A}Z>��[A�xf���8��h��j���h��8Z�<@���T�]�	����b��N�E�l�5a �f����MC��r$IW~J\q�.�6���U�9&�����O[5a�>��i��,�[V��;Òn�}j7��3��>prM{��.��J�kCO>���R��1�6i��Q�HHn3p�[�Vv̫_�����IO͵�Ҝߓ�7��p�/X��*W3T*X��H��"�}rĞ��W��14=ocE�5�����_5)��Yu�%�K�Q��ҕ]��TG^u싶ī�<���>�c�./�KMinVN�?��L��t�[�z_9x��N�oc#�o�:�srm~g��v���d���
G�8͚�s,/�Q`^�޴���͟Wr��- 9�3I�Ư[��	d��O�ٸ>,D��?��d�T~�V[\5�c�',�&��]0�{Pww(���� �T�[��{�'}
���{�i�_3�%��a�/����X19�rzR��̫��#��	�g�N� q�F�THAX�@"�tm5$r�,��O�Y���Ⱥ>�����vUO�=�N�o!�R2R�Y�3,�K���Vl�	Y�"
�����>�D$�?8���i*�,�敝^ց��s��A���-��M_�ܠ#S�.�e�kE���GY�����c��m��(D(����<|��C�U�Տ]����tQ���n�tԹ�hV��%�
;��*d������Z���ieM�Ue���>�؆�Դ�-A�����El��O��D3p/!ys�N�y�9 Tl�"�o��o�dkoC�S��p�3��$�`3@���.;�>�Q��H�^N�ӎ�a`��I8q1��$��̬�k�j3��~��-y�[�������n�
�Xn��ۗ�,;���ϱF�=j�n�x�l|޽�P@�p��x
|���J�QA�����b;� UC�������f���ѫ���J(���V�&�]'[}������e ʺ�jOf�{o�wCC��)e��7�v4r\������f�u��hۏE�D�9�;3 5��W����!���/d�QPK�5�̣]:�~��+A�hV���іLXih�!@�P�t�"pp��������G��q"�3d��f�a$\�kMO��`[U��2��0�e�ʛj8�3=S	�u�i��&� ���m���d�H帑���Y�@��r���.�>>���*���� 9΋����A���*�����x�v)<h�·�S�z��~'�&QZ�(Ry������6'�2ym��] ~�$�KQ�v'd�:��fM��X���6`1���B��)Y�\��l ��
$�(�	������A��Q2X����hv� g^^�e� �L�H�1��'����� ��6�Z��m�u��fq���X�o����W�(����D���'���~�ga��J��v��)� f�Hehx��28����	��dEK��f����
�D��+�h"w����&k�y���7d81=&�KZ��h4�8m�!F��_+��=6��"+p�u�u�Rq5�	�Qbm �"�IU��D����sE� �3��%S��ŖJԦ��L������*z,�Њ�8��U���X�+Z�ܛuH[\��&�{�F�J�sOzb��",�'aN�D��/��Yj��x��y�|��s��E���Iu#�3˞$�4�&5��	�h�@��卢�{���2K��,��cv���םt)N{ͺt��N������,v��F�k�E�b��N�+�S.M1���ޜdH��O�i��R������$�U�,�y��[FW�s���^b�m^��۪s����
̎��)�R�c`�� �@���