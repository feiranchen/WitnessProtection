��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX���@@1�⁄�R��{���-���T�ӟ%��X�=�NS��h�X+�D�[eL8.���jU�H�=B�R��f!�k���9� ^s�V�fcb��k�k��@��"+3����C�AA�o����DK'���ĉ8��Î�cR�ro�?�e����1�U�F�}
��"��G8�
�Y,���5��k��d�sC�p�Y����T�|�X�����P㹑c�N$OZw���A�P�0�5���	٘�.��v<����+����K�r(a~e��9�ReCvJ�����}��~Ҡ}*H[�RFTݎ���g�m��q�4pq�ԪA-5t����hP��((bU��)�maO�|"�$�ƇY�"d�eH����^��ӕ�
O#�wE8b�Ԋ�����;�L8��,��X<Vg�p���|5-��X���9�ՈGa`/}��ˑw���+Sw�?��9"Pj�'9Vzj)�B���%
t5:T��V��cKm�|%�h]�x�u�&��9�>��g�p)�uJ�tڣi�g�=`m4���*CT=��b���M�ț$�[����Ϫ����?�i���)�j��Y������	&��� ���=���~
(�B;wa��vL�)��hq�lrg������[f���Љ!��[~��&�9z��`�Vt�G�8��$kjC7)&��f٭Jٲ�B��o�=����e�;TX�}��[3�c^�s�'�v�Ӆ�7��T�(��_7�?���0iڃs�F��j#�&u~�����;*��`�E�#szE��g�M�wޭ�ɂ���f]Ȗ��!�|.Ƒ��p��
̷6.'`��a�^G^�=:z��|���/�2��OJ�p���a������N�m��>4��d�1r��Z��5��D'���~ڧpX������H�o��I��4��r�����������S�S]lP��Q�CL��ڴ��8�߻�Y(�&5� ��h�`�3��<��G퇶a��� ��n�y1�����,|��y�]l�ߓ-A�VF�[���b�"���R��+�7 �v��='@Øیj�-6�`��h˯�fϖ��cLP���Pښ�8���"�#�c�U�W�0af��ى��ڕP���=�Z��h�:�L�d�{54ܭ�=���@��2Q�1�.9Q��y��YV�a=��(S��!�����D����.t�����	��٫�(����U�@���3�L�8�f1#��$�JGo�ˆ��<|w�]k��r�,��>O<��8�@�����1j]��ڷUyY?&r���{�b5�\�3'�|<�Q8@fKb��Sucˤ���&_V��#�^��8̩���?S�s@��y=3�P:�v�P�pǪ(�qv�{(��)`ua"�[�
@S�<.kI�jv�����$�ϛ�%uۢ�s�',cց��bg��=�6	9)�Y^�L�Y�Q;�l1��X��@̦浨.ZY!s�L���ց+��C�i��9�J�	:~I�KCݞ �*����Y6`�2ec�r'2 ˡ-�+XJ���Փɾx�J��>�a���ƴB�Z	���*�ђxkO�n*�0�`�7/@߲Y��[�|���c�ҭts�]+��nv���x�Ĥ��v�b�����-;G��i�ƩBp���7dT�i�8���Z7�Cj;��;�Ȣ4hW�<� b�S%��ӡGU�;� AED�ȿ�I%3���Ӗ���E��b���Ū��C�2��E��?e{�}�zx�:�wW�R�F�*�&��A^���c�]��a�r��.�(�m��'j��ȇ���
j!ʋ
K�j��a
��{�9����1��;+^;"��QV��ҍ<�f�/�E҆�����saW�]Lt.�pݟ���(knߺF�!{/�Z��e*	WFɔ����T�H�~Q��#O�^��U��	#��_��H
\Lp&i����ӷ�|>�}�R�s�آ����"YvشU�a�pO�W��2�B�f7>���M2�`$��%����@�u|D�J�Bz�2�v MZWZ��x�ɻK��5�bWg}��(�x�ʁ��	�J �t�2�.o�f�`a�b�'��"%]eބX �fe��� �젷[���2f��gʖɐD�������	sY��n�*҂������KD9��xUc��c�P��2�pS~Pѐ��kv�gՓ��~##q]#H���.S~��dn� ��m�
+G�@�h�d^�WC�#�g���[b�Ze�\����1�ү�a�y��#`�ۙ�]��9෋3�|ǈ�����L�2���3k��qcBA��/L!�
r(^�w��b
AO\���RQ�7F�V�#75R����6�q✍��f�keI��3~
F�"��W��n�!|кƾ���S��
�JCB��jl�Tܳ"D��-:1ޑZ���Ш��Xz�l��;<Rh�Jbz��5C%��o�s"���f�{�kR�9�A܄��ػI"Kn�+jٕ%�R4h��v��UYv%T���!�*�J�0#�g_�@�����F"�ir/��#�A�P��l�TV.����'Ŀ���4��M�y�n&�o9�	�螴��/���W��D[���ԧ����� ��,·(�N��9��Ѯ���/���΃v,��k�m���:bZ��{�SE�%twx�֚�\��Tt{L �\�� cӚ��D��ܖ�:2�Ä=��:��y�������T+j��q�����v��.� �*�!�Yw���͔~er���
"�p�0/d�fqAJf�^�T�%p��ɱ����8�U�-)r��GO�x�MY�����7Mue�������0@����60Mz�������n��t�X(]B=�ט-%��`m1���np��\�Qb�����FqQ?��fұ."����l&q�|h��H"84yM�Dfˋ�u��
��.�F	\����i�O���/A)0����߀pt�f� �S,l>m����N���Rc�K�\�-X-��b�v�J*��1�	�`��-	�]i��}��%��V�,l/�Mʊ��$�6�"t�8�AJh8������h��O�1����b�#������դ)d���R/Ab��>��N%l�����p�ʖ
�V�1�����s}6g���0� 