��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��@\�r晓͋�ڎ���ݦ�1���Q|��	`u�yt�W��!J�����7vf���(���>��>Ц��E�84�i+,�PR'9X��-��@�g�'J�h9J]� m����J��������Wӿ*�����
0)�/qI�� �o9��3��k�8�I�pΚ��&�[���#�G=@t-��P/@��=�P3��r���\�d=
Z�{�n}�|c�����P} ����H&�x��=���K����?�xyNΥ]�˛ְ�3�yQ�ją�:����B�[x�,�P6|)�j	�*��Qr������k�65�����������Z�>z�������e�q6��t����q��������m�r]�ϙ�k��A]�<�/���#9�'#���.��;}/M�ψK�^|������Mjk5�����y-g��R���GDi�bg�����X/x�iG����|7������
�'-Q۷�����QӠ�ɇ��<�.�@3c�F��C����>X���������U�����1��������Q��{¼:\H��$F���q&V*����`e�f;��6-Lֳ��P���`3���������g*̎�w�ٟ�Q�У-�j]=?9e�5
u58FWw[������ėJ�sZXNH |���wHe@��6"c=l��/1b�oP��0�Ie�	V�+$�S
�}fr����R��^��.���wx����{����\�,%+���/`��V2(������6m���'z�<V>��R-��^�O�$�ח#��m���P�6{I�/a�k���
*6�L:��1�#uG�,? �ZqH��!����aj�t���|'9����r�nh�
�b�0��y`�9��+�*�:R� �[V"i�?**��tM#ro��$��3Y�a������au.>�b�=��ϻ�����'x��r�߆����GӨ++s��3G�E7؟z�2��ox%"��3��x��7k�-K�Q`b����䨴��������=0�W]͇��Cy��N`T�pSI<���E��؎9�=��ֻO���R6R0�Cx&��
V�Z�oZ904Y��:�:
�$D�~ްp�=r�S@z�~6R����g8	��0=��ܕ�;a
{D!�݆;�����&�{ġp@N��8�U�J��I5���D��?�ِt�)��z�C�tx��S��;$�LJIni4�P�pL�Y4�#)���D~���)��`s������&A8����9@k�&@�i��#�y����@N��d�g�6�e�'��TR6ԑA��,��H��0`�۬��<���%�:`"��MȢ�+�*�Қ�n�~?��wLl���$�@�b���Z=w��agFW�G?��o`4��wڲ�kȀ�$͞փ���%��]�����\s��[�����:�Kb��@�t�Y�7���w(X�]Mc��B���_z�֚f��Ѽ��*��U��
�C��B���?��&�#�6A�J9`DaQ�+.A�l�Ӏ��§6x%P��^�f��ۘ!���[����ׂ2T��/�U�x��2D�[L�N~[��4��{�k]W������#�#���L|ۻ�P%2S�؉�'�y�1
�mx+�hn����-��YW�).L�;�T&����i��ȣ�-"�@��J�	�^MxȰM���}ąe`����+��s��>9�:�vR`[iCy��ga��ҁ%֛�{Ա�-Z�8�@#jҠ�r�$�Ɯ��2E����Qw����kfIMSŪԐe��"`�{&E�\�af؈;?�8l�����G��V7��Z��pwD�o^v[����7�do�p�֢��T�-��܎��z�AW1A�v������提w��i��6x}mX�����M����L��kj�J��#��?P_JR[q�z��
#W�&'z�B͝,,���]�1�C�/��Qˌ�`�)x�&���;�,�&Ld ���J�Эlܒ(	>��F�~�ꉫ(Ea�,�J��̕��S�ҿ�lbh�ȺK�p����b�=ZX!����x��x�F"��i��%
�k�k��FC�R�@[����]s�%���n���
��/�ݮ���@N-��k�Ҋ�$u?�b��Q�Z��s-1SS��-���d�/�f��-s�8���V[ie�F�/<��O�v�ˠ����f�/��3�R��*�)�`ߎT�d *P0+��t�߃ֈ�h�U���,����ʅ8b?3���['a�v@^*�'n��[���9���[��:����\1"p@�z�dw��}�q2�7VW"�������e9���d�H�?��!M�Jc��WZ�6X1~�z��Ć����H/45��ߞ]]]N�TrbC�O��r�\�tt?*̟j�zP�".�q/@g���ήXiM�0�JO�e�H����ԟ|�^Z3Ii�w<fq�,�/U;�TY�ĜC��qɘ9x�S�o�h��;ҡ�_,�p�f{�$����RwM��,�᯵4"�*��Iez�����-Y������1s�q������d���]���xN��Ļ� ���h�8��k�� s~f̱��''U��B|�h}l|)V�I���i��%�~A��Ѡ�$:f�s�qk�CZ�H���e��gϞ��a�X��|ge�J ƨ��j��ԗs��!�L+��<dpa`���&�_X�l0�_6'�4�M"����_�M�a��߾��3��[`����R�nE��~.6��.w�'���2�-�W��_���b W��(�;�߈�t9p'�i�򕮨s=s"��pB�zP���Ou�!�ŉ����A2i����F�Y���̼z,%RL+��ٯ�u9N_T��a?QsA6�Dҽ�l!�̺@d]~���%�t�rߟ&��k>J�?��4�����tuOG���گ=��(/2��#�Dr��˦��\��ѕ�|�v�]P���H�����@�m���8�_]S�m��8��9��&����ez��]m�4X�6�vO���G3�v����Q�a���ǜ�Ed��h'��]�����<���2[c�- ����c��t�?����;�K.lp�Az�Ƥq���R{��g���Ġ����
T*p���r�W$��C
��;$��:b1��C�eK��@(���(�(eo�,�'l n\���ҍ̷�m�Җab�ޠ1�s#ٌ)�{���VU��#e���$s Y�'`x�.�lħ>3�CnN�w��a��Em4.�*�R*:��A�s�G�z�2�;�/�f��FBd�+����8�9d�
��>��󽅧��
u�$��+����n{���_{v�Q�}���U�2��$؈�r7lN��X,�#�^d�Z�W{i�''#�9� ��_��m�8~߳WR{�HB���򵳥&��~��3,.wi:I�*���\{淚������q!��W��B5%Ӓ7|��~҈�0)���ݎ�̋��m����Zi�gs���ڽ&[�D�zI$������T��b�.�x+. jKq�	��\	�`�	�ʷ�dƧ��OF��
 2�V+�*ifh ����I��g*��q�O��0IX�P������v�`Vy�t��c�R�H!P����d�S�H����/��4�����G�����xً�-��(T�_�蜀7�ǰ�8w,�(N��B|m6K}F�@N����� ���d�5|b�}�u3�!�z�ŪM���G� �Kз���<H����r34�5���w9�!G;#Bs{�7�I�4f��$��W���zTQ'��(3�6*���k -�_!VOY[���RΧ���+�5���:�xǸ�R�D��{��o+��K���dM������D��9�t�Q��%V�Oz-M(��4n��ύ���Ё러l��d���}t�teW�Ԇ+�|D�
����pgle���d%�V4U�qw	���3~�#��zS����ک��5� ĵ�0b��9I�Ӈ˴%��o�4'B�db��2!{.FZ��e�&%���q4￬�F<&���4.����/~��Պ׮I�P��b&sz��i�d���K��}b$S���Um?�(�rg=2��X�\P����O�G�w���;:��)O<=��E*�!h�[�[(�P�e��խ�mV��f�o��<���RT�s�fP4����iz�Vy����Mtc���߳��b4��
���r���a2��� z���e޻σ��J3�/�F��/��R҄V���7B.�Ma�%�>��[p؏4�ʬ>]�"�dp5����n�Ⱥ����*캹(��}� � ��E��M�2;_.)E�
� qM|ńع���]�v6��>U����@�F��s�Z���mH�N~O^Y��K�I��`��h�=���c!�?ƚ9�l�=�}u!�������ˀ� �5���U��\����Eݾ��HT���f��[�y7[#��xJF�i��l1��zHr�ޗ��}%uD�]Uk���.�4}ʃ��I�5J�󰩺a.\@x�3M�f�x���:8�eT�_�C��Z���5��R:	�(9�?�(�xU��pB��.s��!�'h΄	�{
��5z�8o{����x��eϹ��.�������R�te�E���
MU��~C�o���������N�'Ks:�y_�sZ� �U�mŎ;���J�z�EK��7"�~wV-��U�w\�xo��r'�>Dv��T,�M�H�d�M�?ۺ.����t_��R@
�bK`*D�����Vz�������[�������)���4aa�?2)��*���[0<\	��1��vj�6����@���%|0Z�X��U���GLi���ڬ 5P!KeKn1*�FÜ�<�M��o�@� �H[�u�	���/"Ao����R��E�͝ʗQ��8g
�����"�!�e�xx}W���O[߇p�"@���Y|�h%Z���k��'Q������}c��Q��c�.23Пd�-@4��Z(G�=
&�j��1��'��=H�tL�T�B���	Z-?o� ⹀��h�K�8�%�;�ɴ�d�$��Ń�}����	`����Jb�r畤Z\���-�n��"E^I��#ޫ�Z/��c���� 8�av�}O�q4V��0	�J`��aR�W����e�1冏�V��P|w|�ӱ˥��ƨ�F��R��,)�^>�z��e.��L�
�(o�+����g ��6�lG�Zu�۬��%�@..��2A�������Ǳɡk
^�7�� ��d��Y�N�����M�>M̿��.W�i=��j�(��
��Gp��M��e��޳�����Gw�3����\8��6�����QY�K`��)��\`-v�Z,�^�@�0�2W����ئ)V�ㄴ1����U���9�i�v�1>���/*��YA�	�RƄ�ji}�{�SOx�մ{ae���7IÕ��Z\a��NV��9��� ��8Ej�� ��K*k���L�{>�x��:���>߲<(�/�3��\ǐ=xS������:�A���e��De]rG��=t�E�,,�Be����E��ޚ	¾�jT�m���9�ϔ�?�: kԳ
�},�Y�?��0���)�L������c�/?����e�cSC���:]����XBRg���*��e��+DL�M>���8!�C�	^��Ӫ�g��6O<�X����B|�N���wO=P	��У�Y�Z�D΃M����|pҲ�NqWc_����>e��\$�e'��3�e�Gs��\еU������":6�nG�L�gxD��,�g>�FC҄��ܫ��r6�i��oIH!�y��Ml�3����X	�d�\�1
i���PS�Y�>~8Y�sC���I/�,C�a��&������n�~����<6�&�'�>�7Wk<R�0�S��۹e���k-�� ���`�8�K������G)�~JېY�ck/���.ڝ�B�ɒ7�~иQ�A�W�r ��.'e8t����Z}K_���}�ujۤ�wY��/���=�g����"Gb�-ݡ����+t@"�0�@n��絥q7c���O6�OZ�,� 9��0拭���X����[��*�m(�0_wK@�� �������q/5�JK��P/+�!�i��X����xNU�DW���}j��/�*_��B��^�5ED� �q4��4�� &5��Z�z�or8*TP��8w>�+���n�����W2���f���F$V>�	/0�S<$4@s�ӊ�Y&g<)_cX�zH�v��-L6{�(�
��#ǫ6�0���RH@�A�)�e�aFF�����%|z\S���2)]������;nl�j�UcK�`��3a�S9� ݽ�ruI�<��Z�M�y+��q�cC��6�%0��w&ۋ;tV�U1�nk
w�,���g��Uk���g�����A��[s��Ʉ	�!Ul�c;{7M?:����w��� 4t�E48�F��3-��zT&S�'�^�����:9�[��>����Gȓ�t���;\��D�T�^|��yE�%1���7�
ȃ,��� u�?�x�|W/�Ծ��.�7�]���<6T��+�����l$~-����"�>�Mh�.O& Vw�"��=�����a=��2�N2X�0=�K�rQh5E�8
)����`]�W Yޤ�b�ۗ-��e�9|�t���Ə��4C'���}�Be��LW�J�6R�M42%9�BC���3l*�O=�aod�%MT��aO�Ν'�m,:w�M���[�k�|��{��n}��")���
�#J�:]�`����W(����?Zpl�DR�!�\� �=�h��l��\[�~?�CA�!�����B�Ü�Oy���#��N��k�	�=���T�4$Ft����X~��/��[�Z��P w*��X�Z���B@��j�?�l�f� ����BC��J餃��*�q�����W�`F<+�6��U����ܳ���G���>�jy��6��	0����b7���}2����~�U�	��B���R4�;Y7Y� (�-���F�Y�$W�7��p" ݸW�p�jE,"�;5����62�h�jAB���k�e|6��BF;3S�-V�	ֲS
��O����Br{��]�a��5�!ۅ����G��;	�_s̩��|2[C�{ٴ��>ǯZmo���`�ռ�������⚊��D+��7�%qb�[�	0N܋T��>��&�h��yj��iIM9���@���R��Qtw��HG��i�J��,h�p���M�U_�.AEQ�d�9�M&��W�ve(,�N��35>Fo��
�[ȏ�����0��7*�	^�(�,�'�tq33���;�
�^]2�܊~�k�tx� ��|a8H^(�Vm|$棝+E"X�Ԩ���)��w�Mf�39n,��k>Z��M�Ӹ�8�Hi�8�J��:f�Q���H��Ŏ�I��C.��Uq��{�`s8�Q��h$�;�*��L&EUp��M�iХ���ܠ�K�*���Ћ ��c{y�-~'�xi������f��\�q�����´�ϊ>� -Xv� Y�`������6 ��2H��6���e�%�Ch�$4�z�=�������*�[�)�X���}��p��M�%�-[wǝ�{�ϰ������Τ���:�~-�(�ڛ�<�R���`�7t������.N9�CJ��1h��h�s��S�[o���^�z�XN=�~ upM�G=��9ۮ�Qw��2���~���� ~��lVkj�V�����&�)����h|�(a^Y/�c�`-��z�sXՁ��O���J��Į�j�O��=�Ƞ�I�(~�Bfu_�2�d��;	��Գ�s3q~�K���r�L�g��)��ʺGR�5]�ta�!傐�\]�M��c��J��	��],3�pi��5�Mz��cJ���%b�������.��?p������8H!�{�#?���ܞک@�������<1
�f�3��h��M�v&��J؝6��5S��+�9zX.jx �1@9��������*������@�Uڟ�jй�!^7�ﳈ�mӑ��+�F�Au��b-A��㨼��~"�����Ν`>@��;����Gz�^QT Ǔ�Y�*'Q�h����_�"�U\?ܿ�!�o�'s�PM}�Z5��'�9�F�.�Ƣ���^�@J��u�F�["B<Q�a�a��p�4&�y�'�������&x�|v ד�N�C�@�䕶W�64uOE���b#`T����U�"sՃ��yR�����,�lS�bLk�G��*-�b9ߟK	�f*����	F)�qy7~��T�ra��u�'9�-����E���l��]¢�#����Y*��?���t�Z����M5����'���O��4���g[f��\�J$د�.~�N���ӽ�[���@��=t��½'����`��d�.a��j*E6����cu.BD�;����0-���_�0(�ڼ'�b,Gk���c�vF2��~�GBN��)�1b��h���r!���BGD�W@��3Q�u  գ��Z�Ȟ�i͒W�����#r��e�?���� "��dM�����%6��E1WPe�LG�.D�BH����WyH�-ы�O�������u����~�yI��A���'�-��9�S8���Su��Ԕʐy������P�$��n]�Fسn�җ�@�bSw��Ş���z��q39����x'�� :� �\��>1�g�;�)0��dm��:8~�r&p>�eO�]
�������c��>T
�\���+I<����8�fTKO�B�}��i�s��qmw�hP�WA�+3���[����<�������fg�Ia�o ��4C�h\��{��rh�bl�������ܜh��'��1���_Ǩi�)<`jе�#%W����#��K�x�`��w�#�)jVy��9��=�.�"���k���Z�ȶF��f@rq'W���Id�̷s7,`0u��"�ۢ*	P�hL��hN��hUe�v�%1>&���Ty�'	{�B�w���g�8����P;���HJ[�*���������