��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX��ז4i�Yئ�=�or
uJz�<|���.��-;֑I���O�L��Gl�e���ko�}$���Dt�ѪL�v�%d�:1��:�6�d?=n�n������۱����7a*G%�C�}>���X�\�7_�_w3�Vv;�l���D?bny,)s�ː �����2Y�z���;͐�,��O��	=�s+�)9���Z1؈e����I�L]4ܩ��U�Ŝ�Kف����:,o�PY>�<={��V��ձ�b��*7mnfC�W�2I�,Z������ɲ���)�[ܭk2����AR�$u���K�OL4j�u]\:w�����}[M�Ѡ&n4DNz�k]��籶�����q�r����J��iX0+S���T�?cY�Ӣ��)͏H] Q5�����bƞ�V�غ(Y�º�nky�o��&��������c3�d��q�#x��C5ku(�h��qh0%�IHyH?�:&ҧ�/�P��_O�ͫ������Z�6S5�"F�so)pɪ�݅om��q"�ݍ���y���@|��?v���Ri�0D��&c�ek������.p��@B�ϑ0�(i|ֳ�Z�%0`���'���r�ɪ�'%����[�X��l� �!߁I��$oE9��W��<�$��>��)Ke�r��,��n�W�G>`1Q;�/4>�>���=3Kyc�ws*��7���v�,&97�p�v(���1��a�Sp�q~0���kRѾO:ů��!*Í	�|���^���1:Ղ�!��]�cj�J|<82�)k[o���q�\���V,��}�?9Dt4���b��Jw;��1c�N>�ȰD�h5��&M75S���Ck��ne�u��dP���z��s�HՋoA�������!�G�`Ϲ��Y�����`�WZ�|;�Xc�q���5�z��o|v0S����)��¬8�.x+d�)C�G��  �����#e�=�gԧesxԽ�(�+'z?��6�(�xb��{�N������_I_��8�x>eB4CB��ё�QEc�޸��PH��5�"3 ���5){T؛��1�@6F�1U�L�^Ѷ���\���˜"�����l���TC��x�2vȋ'��zAh�XX��E�'-4��j��;j:U���g[���|���e:T2�2x�`{����({K�$���^�����G4����FkSm�,ߢ ���@]�( J]A)C��L�t%"dD���&��%��I�6����A<,��6������5���fU���ƺ���w��%5�|G���
&r(/��;Aa�2�"��q�] W�=��MYDjf�ӻ�Ut�\4#f�Z��O;�w@���SjD��G��3�k��w ����&Y��b�s=
*82v�a�7��;��}ǌ3�|�(�j�.� �-�I9�G������>�ww��0�����Y��>�Œ/�(��ۺ-p��?3g/�P�E���Z�\2�s��)��gb�D��wؔ$=MG�1����F�>��e�u��:��D�6�l�?:Y?��^���Tp�f��yD��B^�xO�sN��Uь@�->��?l�'6Z�^Dv�8��p'���K�i����h���#��ؠ�:���eJ��76!���Q���0U�5J0ͬSnj�A��mr	id�0G������O������k1
�|���pu�6e��U[��ϲo���1CB����$>d�`e�W(Gڮ�/dLk~��ۈ6�]t�j�!�B5<\c$U�b�u�?��������y�<s�fH�,T��T���3[�n�d��$�,���'����`!Bt��ίr�3ç'���,�D��Ms�J�e?�z<�-��jh��l�Tz?,��L��$��m#�>'>��SCR/�\t�a�rNt��}�&ǔ���ʇe �	~ڣF[���.�dUhh��cC6�z���}x7�e�w���Ȉ���M�w�\P��/C��>��&i�6>Fl�&Ñ�-��I�*�����oS�*~���:��Cϣ�_߻(���=#Ea��=փ���&��7�=�H�wHޯ�2����R:���ZI��v�^��:Y��Oa1�cy�zwf�*�����߱��R%�i�鰖b��*�����hT�H�u37g��*}��� "�OLƸv�Lh�|0˲kk�����-����?cբf1�Q����I�{er/
(P�$R\Jn��t�����0����y�Du���;����2�&\`��ͪ�D����] ��q�A� �k�E�sA�����k��4*�Z��B+�����>��6��h{�*��-�#A�}6&<R�_ߧ�FjtM�a�]�C�Ơԅ�^�1 ��vf�=]��Fv��H`俢�G��
��sS���#�N�X
zk��c�#[΁�i1 ��i� �q����JK`�q�@���f�M��6��=|(�0t!�m�o�G��`-ON�v���O�<M�0L�`G:�В����m[�k����{��F�R�t%����`:T,A1��ؽrEƽ	]^��]M�_��]+��zĝ��~�h���g��d6_4��,q�U�p�d)�`�㭓MH~̌���W���f��Y��{d��)5X��)� duٳ�"�͵��Cע�ZΙ$N	d)���}����k��82�g��Wd��mrx�@=xye�/��O����"`��KX�������i|s�Q�8U�b��5�s�H��yI��"Bq����	��h�����RA���~؆rX����$�0R�5�\yY
Վ�P� I�J�"�Vh���B8��@����<ߗ��ڒ^����X�\�[����D�D���n���;~��s�����e%	�u��l�ܷAІ�n&S����汧r\MQ.�HL�e6�5MUY2�'3�cѲ��.�tE��{�2��ʵ���@�Ń�&�rv��2��d�@����"�n�XJ%��D�����PMS:���7ReS~� �_ ����r(�p���������[�~/U�� r�����ƚ�KAE��ꜥ�P�ye��!���v42ʆ��~W�f=���p�mq�����tt��$"-QH8����0��b�Tt>d��n���b��V�N"g
�p���x�Q 0�R�G֍��>�Y@3����F�AR���< i��!֚� ��p���=�ǒ�2��֎��S�چ���Fr) �%c�ǟ>�A���<��V��V�ټ�=(ڲ�u���t,�"cr1�+���%#��r�q��7����{W�WJ���r3`���8s��$D�\��hr@��Q�vl��t2HmRS���cJ��p?`����>�T�d�!�w����&�dv�Ѽ@Tݱr�ت��tl%���o�_��<!�i��q%�j����4}_�Ѽ����lv��!���o9�ؾ�iX$����o�?浴�#4}����.����}�(��1���M&�k`BCx�"& ���S����D�S��f�'n��:� �	��N\A��2� �G �7�j���(T}�[_�Kp��Kt�W��Z��;�V}[k��>���zs��,ޓ��gs�&TC<�5���r0�n�m92
��d�n{e���QY�g�g�� �V�qWM�v]�l�0{x=���vR��Sd�a����h��[��>f����pg�es
tEH��feB�		�)�TS4�,L�YU��x��%k9!`;mEԳű0��_;x��rA�o1f�J�LDm�|���9�b�*b�5=j����w񽜸�I�i����<��wj�i�G����"V���UZ�˿�)C�X�I~�����F� ڴ�YqN��Y3�ˊʥ$+!����,
	c޼��l���C�j�l��C\ˇ�=��8WUc�$t����f�B2?�����=E�WV���������v���d�r@Lm�o�ή�Չ1�-�Ts:[q��#a�w0~�S�w[vN�@��7��W˿��������X��J�qA��2�s2�}:Z��-/��i7zȔ��>�E]f،����,����#_�xL�T]-庫A|�饻��1����ᵙ͘�J���]��s(+�D�A.�(<�)f�ȹ�8׊?��g����)K0d��OZ(����¢7гO��#&�`ʅ�P�	_#z����Rnd$�yݦ�AxK�'��l�i����
�t���V����C���#�ƶ"�,q�L�E�}{���^��>�����7b����z�(];�طW�4>��o��/�2.XG�X��J}�F��5�4 �����4A�.97:��15���E��HV����P~��KrH{��*��9g�S�N�s���A�,P��ei�+�����1�a�X�J5��k�&�M��$=�LݰX���m�q�� �"hTXxo������-�p�Mj:��!qT�Á(�B}ÒGh��J�7�&�:�P�J�	y7�NO��m���M~�����9-�����)t�Vu��)+$+��,�"�0�ӳp\��M�I���J2��n��?A�믰U�)`���RD%�:v�aǐ�k6� ��[�]NS�@���ә���}O�����e�_��J�r@�2dJ�D�i �܇�s�� ��&I�R�X��0���(������M�_'i1n_:RJ>���8H������5?���\M߽�S]?͊3��І�-�udbb1?�D�Q2�s�t�c�dN���e���Lx��?�����EC�'�?���~�OvXn��ˡ̘�QNF���]B��2���N�U�	ԍְM�����^U~���#� a���y �:�>�+����zlx���`���6�ދ�{5�tT�������y�(fR�
��:b�:w��%�%.�xu� ���"s S��i/�7u��;��ߪ�QnG���ע�M�OY$m�Tj��<iK�R�>4��[e.ņ��H@OYlyf*��O���YQ���G���PG��CƯ�ڌ�_�w�y�:�!/�Tg�`f�沶Qw�Ѽ?�H�!+Yqn�*�nOiTf�[��F�qZ��xm Y7����2$��(H�Z���9S���s@��Λ�^m�O��94���q7�I����+ؖŝ��"n�tBvp�G>=�|�.��}�m7�l�`s4�R��1��s�<-����cN�f��(Е[#F��7(�b�{��١������ù���ޓ�oD��꼼5��YҲ[V9*�Ё���k���Sa\b5d�k��qg��y�^?
\��h�Y��*�YK�~�
�j#;�#,z�����X��'c��X��式Nb�JGޤU�vsϣ8�J�21V/���U�n�Da�&����1� ���ؕk�%�v�_�1ͦj���js��w[q�?����������uת���/kxλ��yy
vWX��Q�aUH	CY��p;�8x`x��Dn�
 �<�|6�,��tTy�x�ľ����Z���q�l7r)�N�T��/��Zxow&���Y;��i�}�쮍�������R��7w��Xfd��.�I?�\��b:��v���ߥ�(����a� ;e�gۍ�vXȐw����G(e�C}�{i�=�'��j�I���lc@�v�7=޿1��7�<@XDC�%��K��)�
.��^D�#��9���i^�j@�RfV�]�����&.$ͽ�p3+�v�0� {D�I��ǜQ�ԱGX���a�+���¦��ҋ&�Qe�*�A]p�J_�O���xe�e��<B�Z���I�޵Cd��*�ڏ�����s����K=�}�Ծw�Vi{��3�&��Y%p�����o�	yL�T<��
�񼳮n!]~@_���$��)��p�~Mu��~��+�'n�VX����� s^	�O���X��G��0���T��Zf=r+!Ҙ)g�Q�F�"7v�����~����(S�@��Jʤ�0�h� *�Y�%y�}�g