��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;���������!�p}v|)�pB#1�F�hZW+	��M�����^ ��RK��d��$��BB�a�����*(�y󵘔�IYS�0�"8��M�px�	�'k��}2����p�Qc����t���[H�(���H�^�X��"v�v��L�p�Qd�ci��H�z%K�t��	R�Ͱ���1�&�� N�%�ju;�.�b�LO������!l�KWȐ5=� +C#Z^~*���J�J��r��c��B����l�<�޴_o^�`�`����^U+Л/B�t`�&����:Ȩ�'&i�EӅ+e�j�Y� �e��R�Y�h]d���,֡&S�|&�*�J	��A�L����3��w�=��<J -���}R53���R���@���ܔR۝�<�X�����~��e\����n���آ�rr��}s��""�ʬ5��s=��ƒ����gc|��0,'�d�L+N����=��Ik-"�x��&`�?���%4�H��׌,.:�Se��	����%�)�E���@"ɹ&��]�CB���dB"c��_Τ�Ȟ�rr��[�Ac����}{5�7R�{<1e��A	pfqF�^���L#�NT�� ��v��?�l�YH,iQ���_���m*{�nɉ��tKi��\��'���d���g�
Ϛr3NA���Ϛ�A�nN�'ŕ[�;���mF��}X��q�	�8X��*�����3YE�:�X��%@�����%�8oTx����=��O"�G ���I����|��L�3Ϟ���&��ZA�,�_p,L��dA���eJ�����ċ�a�Kj� !<�hzn��O��|?��OV"�.���5]8- �|��Qe����m6R
�����Me��
F=Йr���]��_e�B�Վ!��n0>�	�b���\.W��Je-$���o���吢��ʃ�'Eҳ�<	h��U)שhi8�Fz�06�D5�?��I;����j�V�{�����YH��*7N�+k���(�y"(���SsD��Ζ�:�_�(7�:��܊�c���SeO9����G��#E͊�ԋ6��W<G�D�H�}��6��%�5*ͤ��Y��̯�!����L%� �ˎ����� )��'�du�u;"�� ��y^E��2�d%-E��wp�5L�/�&�0�����[��bo�\�m�3��5�~��{yj��x�E����db�t�c�q�c���#��Tk�� 6W롙������Q��#Tb����3b|!����0�����Íןj*8v���>q&�b����:a����%8��̯U1�5�d�h�O�^L+�X�B�D�nJQ9S56,)�_�m,O�%e8��ҋ8\�-��З �$�?���>�R�%���x$�>wv�i�Y���R����!��~I8l�aj2s,�4=��+������jG���]��=�(7�P��"���6L�PH(��8�M�PU��5;�N����D��_s����.q���5�H/Qj����z��ף��1o7������w���B�b-F�0�!��RY츪?뛾�=�lz__����~˵�p�o/Қ���\�+�x>ʶ��p�^���� e��-w2�k�d��� ��Mg�w�0{속�L�(�J�Ҙ��h��g��<��	��*+�f���:w�z6��6�Y���S���a��EH��.�[r8��ù�f�蛐ӄ9�r���F�U�0�������h,��Z�]�-�!6��I:$�)�d7?�w�s����x<�p�u�LYA�i�j�)n�i#!RGٲ��0�)!��G6�(�[�R;��}O��F��U.3�x�k�zj�5�� ��f��%'�� x����H��K%�)�ŀZ��a>����P	�h��f�D��y�Д�N��,��T7���?��*A���A�o�0�MP޺NM!n࿱�Q��:�aP�'K�b�P'x��N3Vp	������^@��63f6�V˚�o� �K1i��>�����V[��ӟ'5z��|�)��$���\ѻ~�~[O	N���u�h����L�@���J��ҡ1�{8�# ���A�V�< � �ލ�������.B⛭��Ң �ҷ�����b��n��)�����v���X!�j�>S�ԑ��50�b,��	�y$��W�zA1�Kd�$�Ʊ�B�����0K(^�J����W���6$� �S�	p�]^/C���������"��Lh/@����]�I�*8֎�0B�v#�h�P\bU{��C������}����?�[/�P���*���#���'3���)�B�sA�w�G%���]�D�B���?�6hB%"��gM���.����5��G�	A/�2\ElYH��K�����lCy�<�s�I�k����0+,��,��(6;���A�X�:/���<��lU��([LE\�N1��A������/t�v��l��~Gf��DW��L]���O�,�h��뀷H�
�!��k�e9��0(�����+���.��� �><"	��!�a��t*ѬB�"��c{���;3�+�O%�x+�|�����X:��e���?��2w�f4d/�����X�2��ѭk�V-e���,_ة�n��A��)���Z����m�
|c��͎x���Q�G�O�|A�Yg���7zf�������J�6��_s�k��>�vx��D+�;�d>��{m�.�h���z uA|����Lt۫�z�@���Y3�)�;-�����D�v� |D���O�X�g�7�q�Xy���GYM��ϝoD�[�{�E¥a���b���M4d e6wO����MT'I�0�w�H�jߙ��O��R��IO>Ko���}I�+�O��vKz�@.s&�"�m�0�u���Ӝ�ß&�Y��Ց~ˤm�Z���ӌ�Tx��Fv�r�ún�����A����K䦉#�P���Lmu�,�ЪV��f�6�fE[��<�Y�,cJ/�)�x��.q����	ŵ�,
3b�e�7;�슚�Pߺ��3 �w�jڍg�;�⧓���7�=�qf�v��R��[�k�@�5��E*�M(��)W�x`~�X�瘝M��1������Gpm�A���_D6K��ٶ�Y�{�J[�_��̋ܖ���
�$��Ѥ��n�b���c'u��	�k��Ad�[%����!������~���Wؑ���lv�<�L�*/ڝc��-�e�ɭˀY|��p�!wB^���-3����x�<���D��y��;� �P��A�]��]O��fMFU���L�!I
�T�BSA��u�N���/��@�E����؟��A�	�79�8c��D��fU��w^���IG/>R��:E+�r^�R���L=�sCW�8����P�qcʐ���bm�sr<-��/J�2Ǆ�fD�/,�eFn@K�+Y	,�yk,��er��!y�6�@J��@]�u���GL$Ȫ��q�y��1FO��O�6�L?��1o�4�"��g�g� ԻF�7�'�r$3��s[�W2	}>��u��I��ZD*�۳��e��hF�t[R�u�������g	Y�'f%�i��ӆ�{��6����fD�'�

��@� x�߱���Z>N��D�m����tSs������Ҥ055&�g�ɻ�s_3���C!)�h�sV`��^A�-���;��X���`�,�x6��r�]��<E�_����H
����|��%Z��=I}�(��v7T�qJ���"�f�<�{��sY��P'>�Ƹ�P�@BeB��+������e�	e�M�5�\ra���˱K<�)��b�c	g܈��W���l�u�d6\����t3�=y��{en�gf��Ae(}�����3MqoY
�ɦt-��	J�T���0� ��/r����\��6v��x_ˀv����r<�NTֈh�X� w-9�$#�[̢�tj��P�������u��3B�/���J��v�yK�mj벞���d�ʦȠ���VX���Ik$�25(��]�S�{��M�0�
*����Fd/�.��7��
��4�}��ʡ��K�j2���}����QO�>��F��k*	�ִ��$�E�A=��dz����$�긊7�L��2�g^\1D+β���P�� ��Y)��?�����d��Ya@�� ��^���+S���|u�8� �;�l���Ĵ����a�&� ��rpN
@��:�d�p�8cb+�{��	�zu8[�.r�bH�M��7��o}�Ґv�#�w	��
��-�y�P�w=�ZG.Ǽ:��z������}3�{(����h��_$�@T�w.޿�y"g�W���[H^;F�����C(�H�OV���Wr�w��`(O�pV��ZV!|�F:����|<���
�3�-��
.MQM9���5s��<q�^�F,S�d�u����\�� ���V�Qa)H儏Y��-z<��o�4�qY���d����@CS�tV tD����u�ٍ��o[C׽*C����#�3>U����}ܷ����f{$�s�����F8�=N�?�R
)�U�RA	�3%xXY>�`�!'�l�%��,���&��:�7��>��Qx_e�7���6�YP�nKK6`>��cG�Q�P:�`�B�O��U���o	�[��w�9/M�E���~x�j*2�����ѡ��g�a~쿯�ԤIWO���9��C�N+�!l�3�_��_�49�s�?}|����=aɆ%��׈i�biq_]Y'ct\na΄o����w
[#g�-�M��^�4����pX�%�)dX#���3��9�Q�%�ꛧ�B����s�5ƃ`mE�)��9&�x�+�)��(W���b���$o,��m��)q$*/5nvg!*�	8�i�4����f�O*�l�`�w8�?�Y��7~d�7O`�@ �:�$2:�VmoŞ[�6~6H0 �ƪi��G���,D��<M�V��w||�vй�Ee��������3IUX���SX�Q��B���Bj	mލ�e8���v��
�� :�Q���6����f�|�M�@�K�RQ�#�
]��il��P�y(��쮦�t"~Ժӽw5����������鰵�7Zs3{OLj��̔P�t����x�X �-��m}�MdL�N4�����<�.ڹ�{\�2�/��*I�+ ���h��:@�������up̸�a �#��JE�f)�D����@�O�>�rH�J�Ͽy�m�~�B�m�QYZ(�Zl{���E�����q�H�:����)E�DK��%3�%��5�Ii��	˓i ly/06�ͩm�iUϰ/M���c#&�0���q�&���)αw <G���~Ȕ���e�'V�g��'x�yѻ@�l�z.����7��e��+I��(��)vi�ذ�]���P���m��.��anw�7'��O9;�=�s&u��4>���!X�\ ѵ�5H=߸�7"���:�@V�W	Z\,U�}�DƝm�U��
���y�'�����a2���BފZ���KG,���U���Y� �V�#�� �WU��m�6 �~<���c�`��={s�H7gB�J��X�+�Ci��N�P{��