��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���d{Ex�ӯus2�!vD�oa� �M�¨n�E�����e�K���W$�ڢ#QpDV�̻O��:�oV�����E�A�]:g�-�Xf�5�%��߶�ɧ2�<����Y)7����=3ΏT9Nk$!�a�~<��ݐ&��9��VJ-�Q9̅�4�<�m������E���;��K��e6�Y���Q��h3�bb�.�'i�8��:F���Π=�md���P9g.���W��C��t���',�@��W'ЈK��`�ı ��Oz�Q =M�#��ٝe�vH��&��_�J�`����u@h}�J椬d�,>()��:�A��ʕQ��3�N��˯����nz��[8�歑��0��^kD�J��\���P�=s6�*�k�1�+M��I��^��ɩ�<�g@�4���Ξ%f���]����m-�5�#�Vl�;r���l����r��;���v�FqtH�!'���Z "I�q��<|S�Q�����5�W�V���*�:��j����2��
Ʋchڶ������!��~��s�wA�<�6��@��2ʓ��$��@��;,�(���W�`��w�;]���C�v2a��M��ua�>���l�r��� �#?kL{qP�
M��b�ݴū��=�A&.N0�{���V#_ �$���
聈x��tU�=0?��֑�ɻZg��2D���*��� �Auf_˷$ep��
�,)�=�l�7��'&kE�� Q�y�`u�">^7���h�8? �_P{2�n�Rz`f�41��g�pM�n�H��7�]xP�����iM�����?�!�El���D��(`|t[�YDX��m�Ή�/��y9O�` �*�K�h=U�O��s��ʂI�h��	l5�8T�R�Y.Ո��?A��k� ��e��亄]b Z���3.a����F�*��ۂ�ܥq;�J�\�N�,	jx�?�3j�J�)(�Tr᧶lϕ���-�C�z�Qx�&z�Y����H��f�ֵD���%��ZhApd�OtV ;k����AK�kpc�C���h
�X���f8��=Z����ha���e���e!���v�`�.�C�،=�;�Ա�8�����-W<��f��*�Ӑ>6q�bx�ˊG����vn'w��wHZ܂��.���zYV(���J;���wԆ��g��o�����)r�v-;C�-��ڛ�[k{�Ӈ��z{�����S.I��?&ɧi�7 �ڸ��}�~8�ҧ���*#��1N��Z'�#���>ѐ\<rR��&�$B�NU��u1g�w&J��_�d�ͩ���Ҟ��t�p�S%�:���{�_��~�q,�B�7}ut�u� �oճ�Md��(ā�)΀����Ne�����	)�{����n�*��҆�nb>�����n�P�zvk�NL�m-��l�Ǔ���j���@m��:>��&��Z�^Y!BAf�{�jU��H^C��\���/���濯-��f@�!lz�ۇр�e�4Kt�G��D�UH�r�.;���}̽Mk�S�H�jR��z}Lmx�nAk��+'�5< �=*`��0N	�����>��z8�N���!5,�����65��A�LAvG]{*oV���{|8���]��_t^9sB��.ewh6��T-�P9e\��|'*��Y ��$�z.����c���T��յ`S0D��`s�"-�\�����<�zx���B_�J�9kD�h����7���O Wܝ<��t�\
���{8օ����
�s�:�I�J�6Y�[���ћ��^-�KF�X�#�Vu2����~�Y�ҕT7웑� ����z�}2�=��ᛐ��T��k�-[|q���i���NW_D�d��O�+q)ˋ0C�N*(u�1����(jJe�'T�w<O��F�A��<m?g��<_ܰO���B룽��*��Q
z��"|�Jl��.��n��i�y���E��$'8]Ƙ�%�,H'QGs"��`W�E���|'����<a��$;�p��2���q�^֥�-��!�uޠ������tDEb��(�>y�ꂱ�F�oA�.^����> *{i�G� "�6��^Ϯ�=���T�,��)`Z�]XW��PsT� ]j>�d�*��� ���E�&�")�NF} ���R!��2�ݮ"$�]Ā�9�ڝ �\�m#lC\����o��2FnL���`��I�>���y3�������'>�⬈�{	���t��lp�7R�!�M�(��;_t�����1Bf��U���J��Rr,g^0���m��9Y��u��c�iӫK����_Ӱ
_&����v+��e��7�GO*�Y�>����?ٕ<����B��,3<����>�� f���@��#MJ�W8��m�!�Ԩ�
����d��.sSu��6Q9�#<�?��2Z,$���x�t8X�hZm:��떺�/HW������6��՝��5���`����5B�L@,Fzo��o��H�q��/~&LUܦ?���\ri�i>u/����􀾩χ�T�ΐ���x�*S�.��d7�>ƍ��WN�Rj˾3<Qn�*��P#��w��`��<����V���Uo��)T�m��	~���s���D䩎��z��Y���J/Jܧ����A���T��~zQ��KV���G	:��m���c� U�a�aC��
��a9�0�]~�H7�f�qE������8�:��2�����	ƅwZLv�ۮ��I1�`ؿ��> 'J���˞�
�:������J�3~�<��Eh~.6+��.2�D��a1��\@��\���\HD2�w�N��� 5�Kۯ:�#9[s��8�("�*�N�Ԩb@�C�, �D[�-�����m/2{��2FW�7�{�3�P���GwO^W��g/�%���u�~0�G8�̱�:�n��Gc̑3@HWM���f`�Q���+Բ'vf #���Y�ٗ�N�����b6/���������[��Q�HOn���I�����gv���d�N�ġ@�����Ł�v��Z�3���;�����:K�d�;Y��9�s�j�ǖ"h��oC��l��oLw��ҾSdD��g�7b$�M ��-5k�nk��?D.�/m*_�U2Ṷ}:R�ݤ\�]X:�ND�QS b54��V��9f�x:g��c%��.&�1�)�F�I�wb�Gr�6Óp`?�*^M$�sN�V��=�w���h���1-W�t�y�Tt#vḮ�����trA�	�o7sCRʭ