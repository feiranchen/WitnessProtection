��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e��k¢�"�8c��%��ϴ�:���{���h,�f���j���JiY�6����_A1wV���X+�!�V\�Ļ����ZT��+�	d>�,*sPga�V֙"V�I����L����Ą���l_W�{��n�-�m@�o|T���f��ڢuj�R��چ��ǁ,��(G/Ä�>u>����ōY��-ű�r�9�%�C�4��5��E؆�k���)���������]���I�`H�γ�q>��$%�R�r'U\���������do=� ��
�86�رE��W&ܦ�Svu��.fóO������-�/89�\q)�Cp��w�>�]��O\@K����v�Ě�,��A��S&۟�9f�=�@GJҠr�2ӈr�2�/ ����v�Ps���3��15��q�aإ��g:u�E���Er����u5 /�q3�\,	�.�e�'ڥ�(F ��
�U��3!h=	��V$����rZ��A�JA�x���<��ۄ5�8��� l��)��Q'�� ����i�=3�aٞ�Wԙ�U�:������f���?���H�O�y`Mk�Ǻ������Ӓ>=~}:Q�P���lj��<�������.l����	�����{l��X�Y�g�#�� *Ԓ�G�O�҈�$KQˣ/�XԖl��������(�e��r�ބ	���N�E��A�!XL�^��A㗊�i���"����n�mtъg��E����E���h(��a��ԣ����6>�Y��vXY��C���l148�X2�Y?�r�ሄy����P�10�G�KM�/w�0�x��gNڞ8��V��v�01�e�35=K8度g�)�����#�;�'o�8�p�����0R���$������1����ܾO��g��ŬT�,�4՟�Z�X��k5���ĻB�'Y�=ݧ���knI��tF4E.go�YP��TB`zD�t�C�bφ!vy�L(�iJ�_�O�r��G���it���IB�!����Ӥ�A��U�Շ�B�m1{pt:������nR�q*Wڏ��j0��@"��U�ư�����W^���qm|W+H�D��f�M�k�~�JFt�U��F	�%Y�Ě�$�����:v�F��,�W]^�y�ӹL�1?��V�Ύ������dI�HƩ�?���X��g7�ê �����N�ɟw����.3�:��N�qf��X��hp�M��֦��@جT*�>�N犵{6@���D��6�dS����.E�<\��VzR�����AǅYΖN�!y�i���N�i��[rԂ�uSC5�o�o�3���.q��`^�l��@�쒞��T�~�8/�0��T}g�߁r�C(��7��D����F&"b�u˫�F�{��X;,V�RA���M����NB�Mܵo�%I��+��؉X�ap��-��kek��=�C���ڦcq��I^�Xu��}�>�v���Z�AX|'����e�A�ǎ�M�Y-Le/Q�A�y�ŷ�aH��x�q&'��Vd�q��Ǝc���D����*�/λ_�|8��8M�o��q�ե�� G�7[�[0ZR�{�RC�ʳN���KJ�E�Mx�0�I�,y�s�u7E@�!$��<�9��#��7��Jy�0M��ϙ]i�Z�c��UD��繨����J�Dֵ�Q��t@����Itl�5g�ၞ�蔈��,y:`���ҥ�`�k��oUe���H���C8я�i!��vϋ�eY�05�%�l�% ���F�J+�H๦e�T��	q�/3�/�<H�ձ�k�E��u_/��S���Uqʅs��\����$a�@�\P�if�+�.^�t01���h��vI��o���
࿅�ap�
�*��2�@�U�?�Hm�K�$������W
�.Ke���f�۠�����JN����a��%������%�I";@6�e���f���	�	�N���,;���Vë0#~��~�{����)�a1�N��"OrE�h�>~�{��T|Sܭ�2:˳(j�MU���/h �����m츿!�KS^��n��]jMy~͞���l�~�0�����1T�t�����m"��(_��qf��n�)k��=Wc�� f�9?Q���+x:��l����B�+�u�+�q�v�*i�aAy)�c�Gz(ǘO�����	��;�?��,j���]!ī>�f&��&Y�ԡ茓�5���i� ����F`iX`&,��C�zCj3��{��g�^:RZ�� |�B�AŐ��a5g�ֽ�U5������(�&��_I$���
X����� �rdc8¾:6�t�K�����Cm�5��Q�D�d���H�$�')���M�а&�����22$_.}�K�a��G��q�ӻHS��Ϣ�	���Qj'��\4�ae$E����Ja�a6pQǚS��t�1.���r��m��dߪb$�����Z-ǻ\Ϡ���[�t5��8\PF�h�nlN���❆�-8�	�Awo{�%*0��g	�x��j�Xm�B����4�%D�醼d�l�3��"#�8�=
)E��%��Ƭ1��^���MY	_'0qYT<�n7 \>@g�SZ>��'�/M�����r�?�Oq&��R��y��u��|�3� �L�-όՃ|��}��!���{���@��۾V�K�k35;~,��[%"�eO�q���%�饊���5���#^A^�Zv:���99D���m����v�c�,�o��)|u��H>�{S�̨��e��o��*�b�/�=�1���
}���Un�0�^�|�͜ʌ{��bjvQ�4~�v�%]�غ�&QO��h���4�'�XM�@�^f4ً��� �IN�+��x�������a8�ϔn�����J��0���Dzo�C���3Ѥ��Y�b���͓TQ��;�ٺFv;��fH1b��}�����BJZ�_��(,����C}�"\�FW3������z='cڐ����D�w����U`�@i��ߍ?�Ad��ĕ�jt0{�����u{����Y_V�T�������>�!F��-�����c�U�U�T~�7�����iP�{�.
�������@�NV�2R��� ��/��[Գ�X�rjbA%:��y"-��+���5���v�1�N��e�#c�;�)��U[��:s{��2p�ꎺ-#��8EO�}}�	'���v�h���%c◿]3�ieV1B��OU��9L�},jjF�MH?������@��������./H�����IP6x��ʨ�$ �����v�I������W��z�0�6W~'?�;"�&(	��
�{�4ֻ�jq_�̎�{.\��I�x&�4'�	��˶����;�~z�,d�{U�Mƙ��A\�|R�:�+�#�9W���_c��6�$Y��a��%�-�};&	�Q�AO��'�]�k�r��:#!yi���%4UӀ ��;��0;욿�~��ң�$I��eS�}�Es�A@�R_��h�G�B�	"��D$��ՅK	&�rH3-���g� ok���!��42�i�����9�<w��(���ޘ*�Q24�D��*d[T0��z���vw6����_��'%�������	��f�cq�H�}cޙ�O��� ��T[���3���`��`��X��l�ݯBM�-úVy�>�-�ϱ*�!�˴�fE ?`��l]ȣC90ٟ3A��������2���4���­��r��Z�������=���ːaq�߰J�-9G���EDIId�}�!mh*�T@- ?��J���d:!e����j�ҿ�θ�Gh�Y����zu���$�1E9���Eu�A��j�z�^��˷����G�8��F>HhV��p���V�P81y���W-��:jȉG����7�n�S r�;��O\��=|�l\�D{�������y|=�֫^P�괫� ��W�.7CW��#Д@q���*����b�
��e">Y�&������ �����*�FO�ݛҙ��Q�����*1��pkm��T %���G�sE� mP���!q�|'��.������ӞC��#)���̊�;�SEl��c�B1 ���\��j��3����,4i~pw�[�j%m���"�=��Z~M���%8K���z�ﹷ7�Q3
n�;\pճ�A�96�i+�xap]<bd����Y�?])`.	±TT�>�z���M�ݫe4̪��o�RT�X|���U�g��v���3xt��D��<�⇿SU��w�C�c.^vu=$R����d���Nysᤠ��~���M����UR�NkUx�Ug8 S�]
[ϒ!;xYl��w5q�v4U�����J���-Z��!e�Pia�1��i����E��=$�&��I�kE��H� ��5i���>'��E5�On闩�"ل�C�l\�E�d�
&{(��d� {�_�;�3ߖىF�����b�eB��̋6������0����)m-��H[��C O=���x��HT��s�.�f��%-��'H��l��l�΂̿3_OgWٿK�/In�go� ��|��I�����5�	���z��M	�;1~M��k�p�����
+k�(���|٣��4m�<cw��Q7���Ê w��WZ����GD��h���U��σ�Ϯ�:��i{����x����IF<N����|�3Z���-&r�lq�h1��pTg�UD��FZ]��k�K��P���M�b'.$"f��.2o0H��m3�0�6���E"�c/��,ϯ��xgw'B��LXa?��r?���R7����d^���3�͘˲�@[�м�y��S'1$Y����g<���w2�$���ϐ|%�ɏ�T�r&�NDS0w��2� h��:�׵��^eQ�݀�)D���φΒ<E)��v(US�����LY[����&�N���p�6�剚]��� ����T�@N�L�x�-2�j��ve�7��@����c1V����tYQ�Q!��L�`����:C�UwY`i�3�F�Ʃ��;6*����c����xA��V�����`���N�X!�]�-��y��3�,�&k{��RK8�F�S���ZY�Xh_X3|rl���$� ��k��Q�2����U��Uq%�[�����pd~���${��6W7�Ї� �,q���޹���"s2��&M��v[�̶(C�]�]���e�Lk@x7ă�L�tȭ9@)U�̰+1���Ä��"��:o��x=a	�V'$]7A��N?`��/���7	����M�孈� \��Ǐ}m���p�v���/W��ԓ^܀�Ɓ��S�]�_1pH�9pvS�Q=��l�u!)5�����
�#(��tnE��x���E�\L
���'~�E�4�y�
���KB3���g�e��y9z~8���dVK��xI'@~Ƅ�ܟOt-�}ic�{)L�krd�d#���y���e�Ď�P��,;)�P|�

B8}��]~T%z����v��Z��^���і���V���l��~$:��y�tb��SX˕%�]�PT��V�Q
���O�F[��>�S�c����T�C������(C�D�F������7W��;;R]E�ʣ�η<�����˙JyU��9�i7M�P������A�^�~0���nz�'4�W���Yg@Ф�W�[ȉ\����2��?�ו��e><�¸�y ����ޅ�}�آ��]�-��_��"��2���g��&X��Hr�&�=;�i��/@��=[��ǜ�`������w�4j��Z{�I�B�I�� ���ª"qG�Ե˵ӿ�)�k�E��4�{TiȄ�VNަ-}y6�ɽe:����_�U��;!�,��*[99?��1��+��0�&i>Pvq���`�������r�2��ʟ��J�k/&R��F=U���e߄g�W��.�\��N��Kn�F����I�~]���;3������轙����������tIGq���!8ڑ4�#�B^qJ�A�Ɇ�b���p�<S���ж���H��A3���n��#�J��f_(����1��aA�z\/�mK��41Jl�:���-y��7��H�΃>rP���ֲܸ�W=������Y����� ���8
K�G�����ov�Bv�S0 �Εo���-�X�!�PL�8e��A�p�+��Lޕ9�åd%�]�oMD*�c��wm�{���(U�"�c�%^�S���'�Td�W�����E�������Ԫ�Q�%��4��o���{�����OЙ4@�,��֭Rz�Fr�m�5�j��� !�xX�W�ߌ`i�;n�q��[�/V\ԩ���4�sNZr���jk�g��b�I/}W�t�H�˅�ir�ާ`���#��8�7��{rMq�BMג���:<�.�i�j�����kKٶo�h�O��ЩLo$u(w�JO����ֹD��GF�/�&5���v`�0�d�@׈yҬ��@ƣI54ܰ�߲��F�6��Z��4}��ò��� �=?|���Mm��{C4��Ԡo��h7�w�/�>��S<�X�q�G�7��m1��)J\¨e���	bGV�g����3e�M�f{�k���!?%��Q'�fo�<���c���R���CU6
H�a��.=��m?Q
�J�z��I�M�*|�Ns�K�̞U��FL|羦ײu=���|}�ᤍ?�&�aOZܩir�$��Sk:��a���!����S��t��������f�z�aO|�&:��d$��e:�����K��׬�'�����rܶ�9���%E���O��	IC�ݩ��2Ld	R� ���jH6�g,^9	NU����TN֍u #T��ݓMI �0��8~����� OO�O�N�yR��-_������0 �ӊ�V�b:n��R�`�)��~~�V+�ˀ�g��Cd^KF� ����h:�ƣ0,D>9T�vl\cq;z�=�����F~�������.�lm�%���΁�T��~����0�ؙ��<����B�7暕}�^\�a���`T��ߙ��O��N�� ��Zx�Kq�Nr~�i^��G��q�x�v`J��ԉ^C���� l� ?[�����GF$m]�-Ľ(M�t���g�
nV���F�TB9���D��T��>��������o�/�d�^��m��~	a$
�D#���(�0�_�TQ�ip����Of�3WT!
DZ��f�6i�6�� N��o���L��3ٖv#L�T���GUܲ���=��ʱ��dIF]�&���1��~�[l�9FW�F�O��CJ'
��G�ϑ\Y��
���|�j����-�g:3yۧLZ���e�[�x����ɬz�kj7�����xvk��n"ތ�p c���}ČL	���t�:OmC�В5MB>�n�A��_e��L�n�i���%(*?��b�4 ud��؋=i&�"V�4�i�VDy'��O�NW+��������VdG%�����#o�9���,�_��zՁ��9�5�"�e���J����r�8�2N%R�,����Ǥ���� >�m���?������T�!�%R���':2o6ڬ�޴e���>UƴvI��6�Jr�B��eWg��{�����C*' �[n�6�`w\og��H`k�u�'g�ĦחV���i�ڪ���:�M����A[��~pR�.��m2����'G�XS��:�Rx����6��,rO�82��оC���t�+S��7�
$(1�y|p&����WΛ:
��o����h1��U|�R���#�����V�'�dO��������#�z*�/D�VY�2|�e,1z�9I�tq����u%x�d,���,73&햱���"yf�%r��t��]�$i�fQ!�����.��#K_V�����=y�K�kqQ�_�`G_�V[){�͢/z����8�@Bu����3(㰱���k18��{9h��2�/0�Z원So+p���,��C؈�iZ����,3z�D��^���e�V����O�D{O����U
�}+ �H%PIF���c��ǚIjh��1"48��L��Hb#��]B��ɃA��3kj�SW����<'_�6��k�q�[��� 'Ć�R���<I��&$��?�!����s��'��)�p�i��v���|�&�I	����A����b�u8_��lۇ<��s E,[�`]vs":[��KM0$���f\^ێ�=���C���Sh�n��:�N�U��5�*ƕ����K��GSe�hts�5�q|��7/Mrv�Cև�d&I�����>�<l���N�����W��g������A�ȱk畈)�ޔ56������-4�ʱX�s�0��?�!�/���=�8��)F'	T&<M�}R͍q��n�5<SF�b5&1m���-��1#nu��Ɛm�����E���d]�"�̋�r�f�B��vc6��d�F��5*/�h���%4$���ԉ�R������&�/*�tE\��S�����7�wR����e
�ؕ��1Q
�����ɑ�=j��O�98���`�l�j�*H!̰4K�\����n�tˋ���P��S�Mh��J	f���5a�|\�GǤU�l����a����y�%�����7BX��^��!�h��Dk��_!ج��[�iS}��Ϻ t��>���6�SV��C�Lk�G�X���CQU'�{49܁�6��r]}(dklB 5���r��}˒q�I0�*��;�n?@ 0SQR�q����F�4<Ay�u0�8楎��N�Bz����}NA�kqv/R�	�sA��.f�P��.~�÷:ˈW��\�8�qJ�B�7-F#߰����'�H�)���'�9�ۅ�P��x�V7O��S�}���h�ϝ����A��� ��"���(r�ou�{�h�����|]\S�E�.��k�Z!ѵv���=�'�Sx1�{]���\�5*7i�Hc�n	Bv�l�e�n��D��L�ع�o�}Y*�0�:�nh��m��$�,�ܳU]��������d_/"C�F�H��Oj��	K�|��c�R���1�Q�0W�D�@����&�������D�'(;3iT2�/�>��?[=.*�;��'�sTR��#�Q���*�
e�a!6K��7ye+�B�Qp ��+��Oz�>��r �}�'o�m������~���������%4�%���3+z��]��}�C�4����C�;k	���J-��2#%������_*8Jm%����@y�U)���" ^%�`�0�kSU���O��Ɵ���@�W8R�oY{a�]ç��i�6ґ��k�W�{T�P+91�d��R��Sv�aE��K�.�)�7�С.8������dڰzk��ѷz���I�K5�~�Y!A�p2��3U �E��4i��1����(y���S�J�ݼ'ze$bu���.���U���K@�`X%���b��$�U$QvH���
$�&�a#�g7�r��N�۽��Ԓ�C����F�F�GDCMn��S�Lo������)���0`ʟ��!F}U08����lT��4������v9Y�%�*��k�@���=q�6��үL�g���,k?�s E��Xf�D��v�����E:g&������ɀ^6>���s8:𥆯a�<z����f)�&����;��9W��2���Z���؟���t��1w��.�J�� BL��D�5����E������zYX{)�i�i\��� :`i��сVN0�)�NZ��m=;o �q����X�)Q|L1��T��7�/s��9�L��:���w�]1>L=�|N/Ň�z��������[��4\��+gP#��j���Sus]������U�8��AX�C�|:�x�������%����ME2������R{�@0%$���^�?����t��G}�H.��������ZC�
(	�!҃.���g����ۃ3����wr:58�������[Q�P�"��HrU/��~�mSܛe��P�P�;�����#�fc�6�o\�֕+O�G�'r1�i�TS4D[��ō�oaUh ���0�9�8��zG�p�>�4�����I��Yc��)Xk<�ɾ{NBJ�q�<)���̮����Uv	yk��H��Rf�k�z4��x3�?�U�	��Tf�//,W߻�)_��9y�[]�ً��i��u�x�vB4R��6pr�6��$�q��/[sA��p�-_ ���3�a��{Ñ��IΉ5Hۤ���y@=0dg_yո�ǡXёemcL2�S��u�X�|��]�2Q¬V^`���D=�Q�`�g��9�z4�4AL%t�P�� 2��1�tӄDG�q""���I���X���ø�[v^Ȝ�'�T��{⬦T7��i��^�.uq�O�$Pi�"��.��F�e���7%q'@n����9R�^��5�VwM'|��}�	��A����N�m��Ѵ�jk��t���?j�_іQb;&k ����I�{f\�-�9m��f�����V���E��r���nfJꆒ��؜���E�o�ZE�~*�h�T�VT�����W�ip�&�c�!L�f�r!�r��щ�`|3�]�`T�_ك�%��S�KBEP�|�_T�1f�ps8*��:7��P�te*�u�� ' y��S���ZEh�C$U�u�׋�S�3�` �Fqu���~���p��¼���s4ǻi���,�Y�(n�<���T|�}<˰G�%�_�>'���
�_�����y�X��݉{4D�w>.�DU�]���^m�6��I9�o[q҇]�Y�*1���՘,H!42`�,έ���x�c8a�0�p�<�)3��o6�n�ysT��)��nR�;~%f),���"��Q'b/2����Ejr9i�ͧ/na8Y[v�{ �T �Ps7����u����<P�����Sm�����'!ϕ��u2���j�(N�f$��\�% ,�\�,tOx�U���twJ�����
��K�XH{��[ߋ�~��$Ĵx���kѠ'�,Rl�h��T%��^���J�N~3z#���!�q3�Z������w�W~��)�+��A9���ܢ��8S���k+�w�F62`��O�ƧL��yk�.���{4��Rt6���}�� B"�@O���m�sR����e��)d��iǵޤ.��yX�͕�8ܷ��޹Q�; -�<�w� Py_S���kR�[��� �R��'�K��=B+���A:����T�����֫2�re��+	��k	Ta?U}z�K�e)28[8F���*O�iɟp`L��Vm"����C����^O�'#�OKF��/꿱���z�*Z�n���;����X[�%����"�a(����8kAKA��*~�x���e�"����h�n���reR�*adZ2/ ���ͯjM�z�B�s5`��X�����_hn��1RD��!#^M��ۇ���c9�b[&��^�+���^59	 �yXl�#0��w�>#�r��-�Dx�]䝿���7	���e�'��L���J�1Bl��{�o\�D�i�f���N�"��[ZT5��;���3�{��Ȗ��S1t���-9R���gu".Ys7� ��@�L������|'�Ԍ��"F�Z�J	Ӣ�.���!Z�������SZ�(�z�ӷ}T~� �14B���r�ޯ��FJ��3���\[��7��#쳿��k�z������0h�7�<�����ꉺď*Z/Վ{LĬp�҅[�f�'��>M(�n�(��Bc�[�zz��l�q4��
n�2Xw �1�Q�#���#H!�L�S3�(F!�ZX�/��+��6'�2z9�%�ۅ�B���Z�u-&X-�{���	���<�+#O���FGM��'e2�\�N��2}-)O2��s`��sor��3Z84�z�6 >�4�[�͞�IJ�j��kw�iqȬ���<$�X"�{i���|F�@�r��C�56!�te���\T�hj	��BmHyQ,�Dµ��I������<�gت<9��0�F�a�8�@Z@.��z�.������� ���0#�P�d���а�/�˵*�a~0�����Wx*^��ZPb��{��F���(Fo���v���3m�RZ��Y��t�F��`a��@ہ�]��d���[�3�bޚ+�P*�W/�>a��c�#[���� P$COu���
�G���:%��+�E��v��ےO�5K�^���Lc���8<�`S��s18�M�*��O���`�~l�4�ѡM9�>$JX�>m𚀬R����\Q�ݩ�:*��F��+V�,;���&1���z�����J�ؘuu���#L�ڢ� z�V�M�=b��mH�9H�yn��~�ڍ��O��%S��K#���@���dw���f
�Gk�cҒF1�T�Sdq�)A�X+y/ʧ�����9�L�1*�f4��
w�7�{��������l�Z��NG�Z��٦��PB���]h�am_=��_�А���w`��ub,��E��U���t���K� �P�~ ��g6�̋���p ��Is�OQ�S��/�I%{��e�x�6B|!��A$X���Ѵj�O,���=�A���"F	�q�a����w$c�1!�+6Rg��o
m�&H7}�0
�2�9!ȝ1�79��*&���0H�)���<~��i�^�����_[$猸{|���i�Cr����8W��i�!�bB /_s����{�\$�K���#�A9
W��E��ǀK�����D;������1����cMH�t������,��*ï�m��f���Y-' 7T�,�{x�m'<~�2�lέ
�a.�Ü��S��ۨ]������@xU*!~��S�iَ[ʽfD�k��JC]�G�5RIB��?��2�m��E���"�v�� U�(�8'���)���K=[�� �҆%����V��
ۢ�[X�h�,1�>tO��c�l����,����!�����5Eq	�fQ���m*y�Kv����\*��dV�Кn��*Y=<mEv.��Cd�K3!CK<�6��"����o�i�?Cg��Z����LA��`� �V�6��r9����N�Ha�e��t�N_)^����jg6w,��h�B/������w�*25@��S��߶�`aT��:y�90��������m���y���%�M���I��ݡ	00��49Vf�Oz�p�z�q0iCV8����MճԂmu��5f��ғ{F_�&�*�C39f�"˚��IX	ulq�Rv���	�u���;oxO,�Q9Ԣ6&�͒�t�ЙL�#��̽��& �����2��ׂ/ fy���zSL��hgjj�H�����=)*�L�y����n\�xn�G:�yۇ���P͋��W:&����q�O�H�n�-?�#����_�y�?W�hpb�&�<�/��0���;����R�02�ȲAs�?Âՙ�Ԛ���=��=�
�<���;nkV��>Z~��㗃?���ҷJ:�C�\�|��
C��0��KU������`g�F�^d7r_>�mE ���&��V��5\�<3O �<�GR;%'�B~�-�F���޴�R6V*���!�}~��������l�0~���������s����2�X�H*��϶����R������_����7S�b�c���� ;}���wB��^��,������z��䀽�1�!#��c���F�_;�3/���w�����]4v=��Ax��W؛��Y��`#��}�>�<uj������	��	�E�Z�ca�CK7ƒ��撨>st�^<�uD���M�?N3Wa� �r(4
q�VT��&H
#S�Y�N�c�8I�Em���1h�qM�ۤ8�����EQ9A�x��Ʈ�ӿ,����2|w���:")1zҚj��[�H��I+�i�&��/:����k��7��'���V�0�(w���h���4f�a׽��:Ї�d�9�{�
�`f5هZM�+e�ls�OTn�YL�K9�P7���i��4�L�+9墚�]+�~�|;��4V���#�-��J*��� dˤ��_x��fl��Iv�%��̮�i��x�Xi6"��Z!�Yz5�{�����Tش�D��8�أO�x\-#���ŗA���#:y�ow�_��2T�v cCB�T��@��Q�j#*!^�"�}���|�R���V�f�;� &��\�'3��O����F���{�k�r�t;i���[��B���;�WE��D ��hg�i���vR�H�7k}f��d��uQ��]]-ڄE����p4β���DN�^F�d������)� ��~��Ӧ(�/a���BIJ���`5�s�i(��q�ߥ���.>���.��1(�A��*q����!u�� ���a�P�f�tO̖$�Jdމ���^얗j��>�r�!�g|*�����<�9y�>�?F��+���sJ�8����V86(:��4x��V69x���<��c�Y��J��I�Zգ��0�׉r���D���rt-g�(�ZJ�l���f?�4
zyf{��¸y!g��|���XY���`�7�lf���Z��>��������&����I��-|�,i�
��4����=z+�鳞Ȗ~ILx�T؃��f������L�P�4�߹�h�����u�#�����u��&�AB����;Mc[�(�Ci��M򛽿]��$C
E�~��r�� o�憰I*��`��6Ȼ3b#��[���$sd6k�|�2r�� ���,�ٺM#�aV�`*�t�eZ���v �j�$buq?G0�z���텩��ܛ"�@%"��d�g�0������Qf�H�<N�P5n����)�q���P�Οni��I�w����G�5p�YYF��-���jG �m�H�H�����>��%8�,ci���am5�����H�V1�Ng'�CzR�OX)h�&�I=2��0N���4�fVn\���r�����#z����V_
X��n��#t�v~˻�̙�^���dj#sG���*�����O��Q��d u����2ǣ�;g�v@���q�����<��Ru��R�!�~�����%�Ϥ!���*��xq��WY}_������U�d���X!9�C���f=�M%����ǷH`�{���l�gMN���E;hr���u�s�&٭[a����$淂o�+wG��Y�d.�jU�ŹVy��{���4Vo&ۤ�?�A�9���W�hQ�1]�����y�S@.}`�8��ۋ��rh�gI�5���� f&�����p_��P_i	v�N�E�NE���u���?�.&�I�����O*q�������_p��Aݒۮ\��� ��vHe;AеԳlR$�VQOy�#8�HMw�<�z��b;�s\���d5����#��cϮ��]���=��LVϠ��T�j���Z>��h�F����J�7��DQ�����&L%k������ټ�.�a��$+<=����8�<�w��}͐;��;���z�#ߚ��0��/��H������A�Eɀ&�Dsu�.��^�P �R���Pr�}#vViAl�BQ@����Z�h��7��1��	p#��i�̓�<�u`m�-��Y��g�-��-t�2���$�a(E��S�����Z���dd�.TED��Hb�H��p�����9m�I� ��g�A�r�1aE��� �GM�8���l���[}mot�sS`B�p���ɟR���7��rz��ٛ�|���*?u���[1�t塓�9�,Ӱ����KieS~�&���~H��r�ͣ�K�?D(A�?�Cg���>w�=���u�'�8��6-w���yg�~�#�U!5Z���״��`v�ѹ��0=`"��$Sz��VI��d��8��^;�b�.��_&8z�s�qNV���ǩ��{�c	�KPrQA/#��jg5�!�� Z\g�cR�|mW-�P-m���o_�Qg*���X8��tp��c0���h�� N6 �J^H����{pHib� �I��{����m��TE�f��4Vf���K��)Ń�Jp} �ܒE��ҝ#���P�T����Y�s>T��xB�x�D9�O�I�:����骬�eUϑ�a+��|���������j.-|I�8'��y"/�p��S6�����Ye�����|x0��a���������/�wD5_��(�똘O��t�d��x�-r�9�!=�L�|�.UiqQĳp�:v��v��M��HYh����Чh���L[�mFR9G���V���5m��J��诽>-w�����g"��6˯�Wp����C�2?V[Y�?-��ɀ�+�<��H�~M�I�v��Kz�h߶U�>�հ,�喃��S�����ӵ|����RM�R2b'\&�ق3��nހ�����*��D��� 8+$\�Ѥ�I<~ǭq|��H�)�3iz�/&�6Lu<��ב��^��&>��.�Z|?n+����;a����#��<Wz��_D��q���O36G����v��9�
�w�Ћǝ��#����w<ʾ��o~�ǮŒ�O,R^�ś(���wU�"�j-p�|�	V���!c-��2���\j.D1
�G���5��2m\Uڎkr�u͈w*S�"-�"�7���&�N�~�w�dB>uLu1�����h?�Y��j��k�U
.$�[�����8�R_'�K�$���(���$�hx����;'�nAؘh���,-�g�N��<������9*I�k�h�9BO*1��YYR�.�v�J��˧��r3<i��]f��j��拮sb|3�۬4=�:yM>�(����43n���F�4	]`B����|1��:��5T��jR
X_�y��r��ܷ�:	�v/��^�ĺ��"E��%� &,U�C��Va�%�"���WP�Ò��=:��N�����>�v~X��*��|M5B���=y�����'x*����E�y��c]�[|����ԟ�M��}��07��P0��1R��4���}%�0;Q-��ӥ���-���L��niw���fl j��Kp�~�f�Wvhu/Q8��VK)�tU�a�k<���O���L��FP�����	`������lC8�s�6b�A[b�	m��v1oDQ��Wò�G'�JA�����^��mi��ƖbFe����E���X��â!�xu�n�K��7����D#:��V���y���,C	eM/"���c�a�K�<�%���P���H�o3I��{��SD�ܲ����(�_��f�G��Gr�Q�^��k�g�%;�;�mA~T�Q�^]=���j��}1�k��a
x��Gv����f����~�^��'�_�KaT�����ō0�CWX�F߶J�+�f@)b��$�V�>����ވ�X�|���F�p\꼿)��i]F��2�^)~C�.b5ʼ0^}k>x C��S%2?��n�����	#���sCˬl����%�r�i���:gA���Q7��_O���4��A]�,r%��c$�GQs�$ii,b�r��9?*��C:����WT5.(w� ������9I_�]�[����P@�'�0���km��A=��f3�^�I�%H$��8=U�~u޾p#���x��UΥ6��Fܼ�,`m��&d�/]�ܚX �{C�9�:\�1
O���^rVw�~�0�_�1��#�����07���n�~�NC2�L�V\~d�aQ1�8�⤥����b=��@��xя�l�O3���\)����O��8�w'�T2}qfK}@�Α�����Q!!Y��T���L޼,����+���-�-u�k��!U��{_�G���@�M=Y;��y~��I�Jy8� �^�i�%�kz]&z𤋮I�o�y� �0i�q�x��n[�R��x31aC����-��0�ݯ~b��I������`8�*����De��-wM^�<&~H8�x�#4�2�q�[�WzOi��������|�y��j�c@���	���y�df��W+7e��g�ϴ�`��}��Q�Ž�:M��%)��>&_����q�����o��ݡ=����C��bP��t��d�W���(��|����}}�~G�P	4�`�)L�b�2���J�<]_�^̊jҊEu�Mh��C����p���t�'�i�Ò�+p.�/�1�wh��9�	�h�����y^�v�5��|6�#��yI1 ߅BpP����(��T^N�B!��!0�sϒ���1jG{�������5�U�c?Yv��� �*�g�I����XR��f]��ۣ��𮠖�}�����6�����V�:��`��_+��H�jY_
ݧ�մXp�=�Z皜ڲ�ŵ��:�77�QУ�_ڔNş(h��	c�wz>���t�+(t5Q�v�9TZ�=M���]��z�����{�̂����~�\!�蠽��@���zQi?ŖN�X�U[���V�j�Pt-�(���\�I�9�0���Y#�k�|��)�ц�C�(z�*�x����>�l�gIG=��W.�r���J(�1��`ԓ���{��k�S�$�ں-�j�������3sh��K�(��26w�Z��'�������X�T�W�ip��^5�[
<�i�Y /w+\@?�����2��q�.i����:�iE�{���X�\�����z�%�y��pm o.��$�*��]wu����el�����������i�-׌>(����R7Tn�V�@�~�ܛm� Ja�8�(Q��o7~�`6�»�����a�2-��6O}*�����IQy���
��Ey��9W~�3����}�I�@�¡�J͏�m6���Ѡ�|���n9<*��Y�P���-�#Gtl歼��Y�~�Z>�B!%�ΩH�[2�SȠi�sn�
n���@,�s��D��zx~���?[c��9�́[~x���-EQ���K -�H,�!2J.f�5��h>=5�=�[�:@D.r��u�U�7Q�3�`�� �����uM�LѦ��Y�X�Nh%i�M��&�U Q�G�/��Ih����B�=�bYH�X�e��tL@G���a��S�ת�ڤ��?sJr�ی���J�mwm3�,K�:d�5�V�b�����X�W~�0�u5-�������s^}�\�#��M��jN�;ҽ׫(#��*� �A�N):x#v/�9Ho8x���G��̉3�
�6�H���0W����ބ@�a%!h��x(�ǫIHy^	����\7���T�W�N�Q!X2R��
t��Q�1Bō�O\lϻ`x�g<� ���|�$��*��A#=�jR��ق��ħ����(ߚ�-��=�h
=�Y�̬e�{g>��
�ߟp��O\�+|x	��Փ��T
;>����Aޖř�b_�c�ǜ���N�yB�+YL��Quh�;R����e#�y�i�,s�,s"��ea&c?(m�dG�[,��ב�D2'�&psQ���~����?�Jw+��/ "|~�x�k�1�O���n�۲HF\�T|U臰A�!�QYAhd�f,��)��\�<U�Nۙ�����={ ����;\Lt���*���m�|�����T�(�{�~|5X�ȯ�k���x���*E4��f:Ba{N��c�Y�E�B5��Z6�.2�A�J����h6����c5:��ƋnZF�˷s�_q���^��ؔt��l��"�k�U��.*[Ė�,�Q�:Ǵ�@��h����5>3��عf��E��)ۦi*�kfy�O'H���a���9}�%�EV<�. ����Q��=��ŗ��fw�Ɉh�N�J�i��M{����Z�n��[�,x��8r�A���
>[��^+�%���9���n#/=�����Of+�w���U��}��-ː��`��}�>c�<l�ߏ����[�f�w�$I]ޱ1���V}�@��>���1����Om'.��� OL����;
�݀(čp։�� ��b�Q~?}�F���~���h�P�}����UV�?T咉�x�:mѡh͐�ľ�S7;�T��-{B�7K��dF�g��'����A���4�`�
��B�Z4N��E�D��dd�IU<|N�8EHol��-�8��k�)�	���uh6�N 0���?���b���ۙ(����4���7�J�>[O��}�5�_]���oL��6��P�����	щq��٨^�Yz��£��#~F�ݸ�^��)-1�ZT���%'�NwA#uZF���~%/�V˱�~����� ����4��AJ�B9 �{>���+/�� \��	RY׿��\��V��S�1�����.]����@P��cT�l�N�5mZ&�H#�O���ܺkkD�!���EEy���u9}e�Qޒ�4��w������P�%d�F�
yo�PL��>S(���咳��D� �FW�j��m�q�>a���,�Y�Bc�vh�n�Y���kb�CW��i�W��)�yl��:���F/[�%O��0��v�º{A�>��0zI��x
|�g�Y�&����y���CP4���~0}�ξo.����׆�"�Bx�����^_&��/~g��ը*�kp���������O@.��e��9��@m������,$.��A�LL���@�*=�V�2���&�iU�1��|q鈃i���Ik�N��l�줰.���b������4g����7��|�_��L�q@ЧZ��N$��N�?�`��ɸ&1
ЈQ���	j{��z��><AA�x����5� o
�	ܶ����.�mΛ��]��?�#�ԉ�/��;% ^���{�Ԟ#�0�����,µ_B�^!s�Ɠ�~0HY�n���M�UL�h�Y_��b��+#�8����l�h�]�m���d�H$�dS��sb�ч֞�d�	]����u���BzVJ��ί�J�r�k*�:S9����?��J��\Crp�7��=�i���ˊ�V�=H]xy<u���2����Ql��>Ph;��b�'��X'��o��0�����C�|�ك���=i}X"��f՜Ρ��f�j�\�>�mg7ӣ����ظ��/��@4��0���~�u����D�ȇ;� �9���o���X�v�����Y�(���kM�a�6��|F��#�'���W͇�v������,�<��E��(��fd�m�,I��U'
��E���"6�gQ��3�<~Ί^����9���� �"0_��	+�xk]�B'0���=g��c)bH��[b�%d��x�eAV�5�8(���C3��	i>"�{׉: q�V��H��\T)�0�E���8KCn�7K���}���xw��^�Z��Y��R:(��Q���4M�$���^��V�'�>y4��F��SkO����|��~�T)�9B������s!�������4S��[ˬd�����bm�U��5(���x��7M���*x_��d��h\�������٭	)�{-
�	{�;�q��_�k�7=�vi��VH~��#^�	*5�/�un=y�+X��mv�O2�9a��G=��%l��y�qa�L�F��1�Ť�����`�t��g�����Y?B1�
5�C���M%�i:�R�!�������l�f�^�Lq'x,+��յц}PT
d�s.�1fc�VO'�?&T�i�@��Z�)�xʏ(zu^��X]O2��I�=Wu��x����B��w�P���9�׉�Ь�	$����C������e3��72C^���Pـ0=�*̠�9�A߲�̭���͎J��u�0�Ұ��m��.d�Dz��<��Ğ%�j:qΎ�?8Np��nL,"��7K����2ȍD��2�ΙL4 ?��P���Wo�&wI����������o�M)�6�j�/LO�(��|����b�"�c�9|�l�����[�X^�]m"X�_%"ڹ
��D��Q�s�x;l���X 5�msŠvt����&2 ��s2H 2x�7-��`�i��<�
.v�<��sq�Z��^��"� ����`��#GM'�g{�����kH
��"�Xl��׺r�^gA��.�1�̹��Q���A�~Y}̜&������]>q�ʲ"���`�Z�&�����Zv^X��Z>�Q�s�2����w��a$���1�;��O0����b��?�&�^�����,]�A^�&�b�L�Q*:�^̖�f��)���r�3���o�hV�J�DŎ չ�x����R�g�������qn~��dj�����	�(�p=�|�����U��.�0<P��u5�7�L�l>�2$u,Qd�] ��
Y���bNB)�pw_��G|o�	/*f�sQ_/���I^c��e2�V"�ؤ|�l|�R�B�*�O�^EYU�5�]��$�n��~p�xY1�i�d:\'x���ճy��1�GwVֳ%�>���xJ-���/N��/�Y��.})P��RBq�p��vٰΩ��u&���`s��$�}��2 ��o���sӎ����Il��4Y�ݔ��	���i��"y5�]�48���Ry�Ĕ��h�\r�A�-�]*��פ���-c��?��l#��L���K_�g-���׋C���M�����`3WXhr}����/lm�B��%{51��ͺܲ�sDj��A>F:�#{Bzc�Xg�nuW�Þ��"���1�+c��������b͞K�dE0`삌d::[��]�')Q�9��f���\JԾ(J�2Kb)����e�45��(p����ħ�uê�ML���#�5}W�˰��ބn5��o%ݶ�½��q-���F�z����\1�e�*�N|�����Ԃ �D
ވ�Bu�Q�7S�<C��O��T]T:��'��S��9��؜����m|��N�2�@#����!�UÇQ�e�P�[(�=�&�ȞJ��ޯ6�l~Ē>`ұtxy_�q�`��D�qO+����쭯c�]
G�٪uuX*VN�ixX%[h�_]��s����O ���4A����5��򁨥c��MLg�4��|*�|Ug�pԂ���g��||E���9:���۳6<��-BdrWgh[yt��.����e�I��0�=�����[܆jT�P�}���Z);N�﹤����Z�+A<ӯ���\��BmCQ�D��F	����8D�ǣNR�GP/��p�~mφJ�(�M��Ήlk�K��[�V!���r��cm&ռ����=�W���R�U:��C��xЍ��v�Ǯf���l��M�k�@w��D�7��7G:����l-�d�,s�>�{aj�(_Q��V2�E���m���V�U-�^��[
F�ؘu��8'-Is�V��NLϰ>�M�����t�>]xJc��a��9���3ٌߓ방�l��O�p�{�y=&�߀�
�x��S&����e$�<��q{�Ïp�o���N�x.B�nh�rSww1\��2�m1�l�-�)�C���\������X�G����V�1.éhŅmt-+��Ѽ�.�ܙ&Zc���qb�=}ޖݰ� ]a���4���o�&�\5(W�v>*�g�P�#(�B�g
�G�!7�Ȃ�o��� ˕B��/�F�J߿	]�OX�ġvE�<����<<j[Z���7�,�_Q���&ntq$�+��*8��Z��|/���D�h��>�B���-�l�Y�{��� �"O��x�y���J�>&���쏉n�\�0u:�8ajA�����ǳF' �$���@�M��H���te@�o�x��,���	�V�7��YG&6��j���5H����9Й�>A$]�Y�y�$�gA8b�:��-mU�W���}��&���8�||>y����3W:5�F���시���Nb�@&���-EER�xR��3^-�ʋ��1vR�8�ܨ�EEE_��1�A�լ���2j\©mŤ�Q��(�Pk-~;,je��ʱ�3�Ι���Q�/G\"g�2�%��Ý�J�f�E��.Rf�)6"L/�+�H1{�jxJ�/� ����e�&�Ou$��P���)�>��<����D=5�}8�%Z��L���
�����F���Geo˻ʄ�9/�(J%np��jp �#kf�u�&�� !o�v�~ã��l2 ��܊��`�D�f�q��hL��� �4�/�5e�\wѠڧH�=0-��H������0��{q��
��ȝ��:2/h�b�UQ��U�u�/�ҁg��R��`���=��O��;�;�TZ�=�W�1��>4�,��a�	G}�
���C���+d���V�����|��nm4�k���H	�E�|F�肢D�Wъ��B�f�1��1f-!E�7 5�!�x^#�۶s�R|��b���	�P5�g������<�g�3���E��a �.����R�q,���4fJ�9����0O���n�6-\5��?�&�0�oߤ?��pj�/����h%�ef�E}��Ճ�"*g�!�H���T�բ��Ua8e8N���%�[>�Bܚ]\������Ш�x	� �}����CHk���K܊ z�Kd�ʧ�Ok����Ig��F{�ܐzs]ֽ=2��J�Qf�M���bcL26]�A�?2�s��0ȉ���?��N\?edy(?l��C��d�Eڪ'��B�T�L�4R��c�p�����m��z�����4¸�S�jҁ8�F�ǈ)� ��'�u��g����Ɨz�ȷq���_p2ԉ9#q�>�xa���˿:�Ply͟Wb��3]l|ՠ2�f�y��|m=F�|0=������`�K�ς?uь�_C[*�O��-|>�n��9��ֺRÙ��{��Wb��ɰ���v������/S��mf3�=�n���hqK����@O���P��v�4�=m+�N�o��¦�&o__F�+��Ж�og�O*k;�JH�K�7r%˳*/>іE�쉠� �sD2ظy)�$�ɲ�D��3���V��$p���W[���./��S�#<;�ȡo���z�*g�lO�]W�a{:��pLy2���TI�ĬVkT��^P���p�#]�����6�i�XCi=�n�3�d�I�.*��NN����f|�#�K���<���,[�^.����tqz/鄄ۙH�_i�P�F�J����r��L7a;�\L��1nˑt���,�<��T�귟�0�����W��^�P�l1��u�,�����^16�e�YA"�W��}|�j�E�G"�����*Y�#�mO�� �|\�i����i�?�65}�Y�՟�(�vv�`�ӽ�%K�D��~�ZO
�*�g��gL��x��9������l�t��N[��w����P��W�	YN�tk� ;��Z�P�3_ӎ�!@��]��X7;�]t�1f�#bx������"ܤ���=�"}\U.mB[���%ʵ�L �dy��Ļ
�r{�,h�ם���{�� �F�.�3'�����bn�^�f;6�j����qk�֋_ц�ِ��}B�߉�-�D\�a+�l��o�m�8��ӕ�o���k�4��h�NT��{��|���;�E�b݀�gv���t�9��aO��w���R 7=�If\�'�"���~Q@S����cW%���y8Rucfx�� �=�FZFx�d�Y�p�Lѫ�&�_�B�#��9����>UF�����'ZsAА�J���i��edji��`!��#�@��6Ԓ�冧"��3k_8NqP���:�k�"�wY��i�Ơ��h�O��R��Σ�S_i��-Mo�`�O�+ђHt�$�B��;���}���6�����\K�c�עG�O�)(I��]BOU�,�k�+uqj���<���ɬT���tt��[��FZV��d��o�fy�����oF{����M�A}�J�[8�~%��Ԇ���V��Zkҕ�
��������_6��v*]�GN4T��e.s��o{�����J~��O���l'�+-��$HÄ���(x��ʝ�+Ij���PRm_������iwW'������)-O�'����I�)�9>m�d�Yhp=m���[��<\`�UN�Fwb�a���~�����3�l���`��Z��9��!9 
&�87�)6�k��X3�zYc�t?*���n��>�\�"V����(j������]g�3��~ɠ����DT��Ɖ$f��6gj��*���9����w�I�z!*u�,�*����GR�7�L���B՘D1�h�P���!�hq��	*���Z�sw@(�r��N���4�&H��-������a]�(V�a����M/�E�Z�)��څF�8�
֑tE��6!�4&��kS�1�T��En�E�� *]1|An�w	��$��Y�1�]�X+B����[�>��&i~�.�biZ���w݅���VĤy��S��4xri쬠�2�F?����Kq!�MXu��(��Ie���!Mv� �����/ugQ4���k_��]H�ސ<eV*��[ʙ�屺?
&lGAkJ
 �������,�}I���l����W�լ����R��H��� Ì`E5��@�#�5}�#;�t�Dos2J!1�1�p�����12r@DT�`�������Y�6�ž������/F��Ւ���B��قd<d0�e����e)�7c�-I�rV�]�cU�C�#�,�"O-�(��þ"��S���Q�Ҕ�?��֦n�qź����s)�D�T���6ϊ�u!E:�$[#Dn�9#53��lOF��(���gZW�F�6(��/�t�yI!�Q�С���VM��O��m3فQ*��e��,PH�xX��I�N��s�a���N�R)�G��ۣ@�����9-�/�̆�h!�k?𬡼ִ�04�*I�["��7hI�b�@2�0~DO�]�^�	�� �X��\���!N��TT��CVJ�ՃI��9ʓ�2�\�5��R�B;)푗��[��,3CJ���UJ	�M/����P�����;�"sܱ/�lf�-"9=�U�W�X�"xW;]���ç���ZU>������N&��	%@��?��̈�1�z�Y�۪��ԩD���Uv�QH?ĠϽU7�xk�߫�u�	W������q٫N����B����Ģe��0��X�YF�f}p���Ff}ؒX�U���暂��N��)��pĝ�|��ܭ�2`�d^	����<KQj���5�;#/C�,܅C��V��0zI�~u_*"O�Vn�%	9���K��'����Z�|���X���� V�5���`e����KR:ZFӕ�z'y�,������e�pg�bi#,��xj�!h��Yp�z}�9B���G�Y�d�?�H<��\�e��������L���}:IYs{n\k��B�v':c( <bZJ��-�F
�d�OͶY{a��<����Ɠ׭~Q��Q�b	K��#���֔����{إy��6��,h�헎2����T� �m�ؗ"2�P̀�3 ^z_��!��&Io�0��g�u�YI�R���hk=��$G�=�mX�&t����H	n��:�h+߆����R���/�R�N��7u����G2�˯����Y��1�� O>�	U\�ѹ��.��5�w lC��~��KSR���D�����D��=����O�X��ϱ��X0�'~��s��O���k�?���A�Ԑ"� �7)u�G���`p����ƫ��] 9v���w9{i�UO�[	5�(����o?�F��vs��m�CX�d�e�}�\1H����7�u��t̿댴�Q��y&�4�D�h�܎���רJ���k9���1����k�~�E'F�7���\��~*�y<�oI�1@�Ǿ�&�*o�����;h�Ȇ<��Mim�l6�F�	(l6K3'�~��6 L#��d���DЖ�g��ۍ���H�C��Ȝk^Dq��C����}�� ��F�g�,��°�W��z�G �Ţ.�| ��!n�K���oF-�%�c�8cSv*��v(k@����k����Fq�W� 5-R��؆aF�>:Ū���g�J�oы�D�|���/��5ݭl%�_}�?D�B� �	���d��u��[��zQ�d��bcJ�P�v�"j�3RaC+�'l�;6�Q�A�Ȝ�Ns�PZ2�WٖP�|:I��O�ǵV���m'�\�A�!��=�J�<z>��� \g
R��+���b����z���,��'wH��o�`�q��?׉�m��Җb'���o�����?�@uoS�15J�QG:�kKOd붻���ժ_���1���W�����2�7���[]��b�u[�Pډ�"b��F��E�B�!O�0��c�����&��VY�1K�̝W���/��J�����n��2u��L�¤i��|O2ՑE?����}TS-���"��
�B	��l���3m-�ˌ�eM���R"��V{~(��!�E�(���x�D x�@�cř����'Dt�
��U3b|4�N&�+�4NcrfmIw?��Ѹk���jp#'������)og�>C��R�r$~��p�F�J�	y��f	�q_'1���-�_t%�R�臤C��i�%99y !�΋�켑�k<(���P�W�_�Պ��fs�����:w=0b3<��[�,�qu���#�fN��[��q��08����%	��/��	)�A��"����M�Q�a	�y�;�N5b��?|�2�Z�����je$c��%^�o;�bٖ�\���=�~�6��m�g848mQ�#1�$(�TG?���2Y=�y�|��X�6҈C񎠀�ԼK��&0\����>,�ZG�����L	�'s�"���Z;����7"s�xU�KgX��V{(�.);���'j��X��?���G��)-���:�	�2�*Ba�Ow`?���
��`To{g�Vx�Z�Qx3�Y:��Y4:
�CR��L�)�[�O\���puT"��e� �e�:�� ����D��D�
.�[Nv�P��>�£~L�ev�{=�V;�x���(�`��k�a��H�l��{߁�����N�#��U�.=�!��]�<4C�!C~�(`�C����'���A~"PF���7(L�0?}��o�#DZeyF'�8�A]t�%v�D���t��B��, ��]�O��;@��h��@�a�MaƓ�ȗ�@�c%%����&.�@�v��5*�tY��^��e�^�_֭���1\t=.��>\��i�!4���NJ�h�f
��tM�?�X����茫~K���I��[�����%!�lT<SDx gΜ*��9���b��BPW��oy����~Jln�l�F{�s `��î���G0r[�O#	U�^�ø�,���?�}�?g��%�X�W�A4H�-���fm�y\]k��h�%s�lKʀ��|P i����K�e���^�]�~���[^��������u�C!�%��9������u�8կ��6.�Ow�Z��ʋ��Ѱ6�&�R�Qqa���	�w�4��>�^��(i4����qhg�J�VOƻ���MPN���83�� ^�X��Y�r"~�ѧY�Y�\��"���t-��|���{�^����Y�Z���D�9�A�e
����=Fw1bCƟ�ۯ+>����mZ����_�d���K��x���*�/�k��.O���g`�T��r?*�*�}��U#?y�Z�C׺���׀.��ʜ��(�Ez������w.u�˃��?r��qh�ܻ�V2�4ܧB?O�ϲ��}����)��0ǉe���7�A�1��4z`4��l�F� �=�q���w!br�ܲci�*	}�N��Ǹ��c�;���Z<���Œ���D6a�\f�I��Rj�o��Yܺ�1� �º��33��I�y���L���#9D�E�.�]�զ*���p��!�A�h8]_�~tm����e�ⱜPػ���03�(F�fC��oQ���I���V�R��J�~F��kw\{c�#~�H��\�q�`����s\�c-�Q�G�=x{���/���]C���du�X�Q%�^��-�\6�.���t�~hy���`�fI�z[> ���0�l6�|E�7s{�oKX����J�5�����ꖕ@_����K3�#�_zA)�'GC�SɦH'�����ĉ;�{��6q!*�o��%2aa�p�� �ØgK���JC�e��Ŕ�B� �&��IΡ[#�!�])�i1t)A4ܯ�x��5����ܫ�X;�Y���w6{HJ�����b�s�ߚ%��GW���.x����LL�x��f�bZfc2<0�	ns0#NB��Zq��|z(�A3�f��8�dt&mY��l���)?�e8����d+����ѡ@�(w`�h{�V�sD��"T-�V��N�Rf@s���}
O��:�<j��\л[re��'uQ���z���)��܁�a�-_�n�#2�
�@��b��T��O{�R��La0��|*�4`H��Ԗ+��c�u�%k���<a�pٍ�s�T�	0�0�������'E��j�S�Ypu��\x��˰qG���=tHyx�h��z}6�+HG�_g"GH�-�`sX8bL�vBɓoyc��P�[�t��tæ�^����(��Z}'�ٸ1<!3,,l����
n2���|~��3Q�F/��E­�m����r�h��&�*�&r�j�����zI(�л�L��" {!�7�4(��& ���C�i��vS�� CcVdJ�E�2#
�Ws�����.�DD#���L_;�1c�Z��J�/� 6!V��}�G���h*a��`Ye�����,�y����}C���S����湸�Y�>'ַjwe��G�W*�Jb�܊��[�SHơ�x�a�������dt�r[Õ`eP�ǰ�
ı�핆�Ќ<��@�Op�
>1p�4S�qS= ���B��z�R?�D�t��)q|Y!�����J�!�2��K~EO��pćKnN��D�p��ή��̖�:@�s��m"l1?O*��E����r���A��X����i�4O-�GT8��	�*tI�P�~�����Ɏ�\>�1Jt\#����Ĩ@�����i}��`�i޻����J=��L�m��^��eB����̼U(]u5y�&O���UEڜ�����2�+��^�fW�h���|�$)�>5�Z�kҏ
�������9�.�g��zl}p廃͵a��m�ܜW4�MTyD*k��ɜSL7,���7�m�E��̡�h�����Aʐ�L����-q��M�UA`����Xq&=~�����E*!(�S�|k���p��`#�
 �/�-ٔ�GT��a�|tf���I��!{�^k6w��$����i�j1#�������go�X/	,;k -
 l������j�921���2��7z��FK�
m���0�%�w�����r�\ǯW֕B��l��U"U�䯟$*�+!!����E���X*�P�"ϓ�`X�����E���.oQ��HIN���pOX��8;�`7�����F�'�\�����lO���]TA\���۷Q�:��~�E0����+br=ь�{���;��M*o�炼�p,
2�ˢ�L�q�	F?�1ξY�g\���f���O������+��7g�J^1���/ʁjg��90<d�������9.���-�<I@�p��hJC0�˭�m^�06eߕuY��&��~�erp�eCۑ���&�0bJR����=����I��M7t&�'��,t7.9��A>2ë�:x6�z�3� '2u�QL*�%�K�N8.�W�2a��g$z��G�GR�d�n��K�c(�����K��$7�(�~v/M��,��P �w(v-]��h<K,>�-[D�1�U��ݡ�H�e�,�&_�+OP�"�b���pr�%N���p:�p�q���R�r�g�2ߚC�w�z���Ȯ�8k4���ߗ��C.�d���ӝ�V��E8A���{��Z��地-�֖R&إX�C��/C}��-3^<o:%��kJ!��Q�gm�:���Cz( ����U U��Oyf�*%�`;vP�x��]gIf� �{��w�!�Z|i١�W��'��+o`����J�1ŬDkld;����s��x�PD8w����\�r�P��]ʥ#y��&�_~G� P��2��S��`CMe�'�M��+Y�fh�Y4��ݰ��k��i)|�.���Z����N�)d�ٖ�2񷓪�~�=��+k_�m��6���$���
�8{va�7�ܸ0y�����I��BK�5J�1w���`�9#'�`�BVN���"b��xJ��5����:E#u�t@!�G̋!�.OZyA^�38.gm�]�&d�^A�PC)6굣��=c�3���9I�F���"�f�e��]K��O�3�@7 �`�z�(Kp�2�R�;ނ};��hX�'Y<�\��B����LDot�X�pD���@Lb�5d���z3��pW6��r%4 Y�]$�#M�]x�}����?KC�97�H6l���c]����s
w�GWx�MaB��U��S���#��u�~e��ۅy���>��� ��--,Ȟ6:�7s���v��0F�+k<�PM�8q�?�%��5�dq(98i�`�1f%��6/b�S�9\�E�t�����_�W}Q��NeAu�5�3� �]�㐭:I�]�/��5~��ws��3Ҏ�W����D"�Q�K���p��<If�i�ĭm���;�b�I�R�E�zZ�2�tNk�{~Jg|ĸF�ذ�^a	 ��{��C�*�l��t�[��Y�lLD�Kna�c�v���D���9��׆�6Ϊ�F�w�wEٕ�qDk~	�M�"u6�k�*iw�dl�_�p�Dd�eT���n���
��>�)׷^J�1��l��u��T�2m�B/�}&���x5��b�;��)���ƽ�it�~1�:7�	P8&�x�\U�9�ZE�D�&�@yu>_� �
�%䭏�i�F�t�g\�m�r;��t�E��H�O7���s��Z����3iI���x�U�%Dm�ة��{؇��N���=`�ҢXdy:iOk��b�]�����n��w�	%���D�������k��+3ȃ'��^�1l�?�d�U�f*��I�)���eЏ��:����m�8J�7:��O�h�c,=��jJ���ryx,��W���;�������� ��ArYH�PS��O�� �˙�w����-	-�v��RE�q|��9vQ���-��'�З���a���#���2��8��G��8�uHt(��'�]���<�hZ�Z�{�jW�m��mV��ʻ�"����D��^�<��y˞2C[5z��M�*|3O,�֨1jj�V���Jw��W��:���d����D-ZZ�d�_S<� �t�Vt�ʢ~9d;_N4�!�.���ċ���[(��T���B͈w��$��FF���S�L��`�>M�G��b��|�^�B��M�z�8 ���@FU-~��Z�WV D��1]nMM�c�Z��$H$s?�����xd��<
�2����9���noT�S�$9���G&��o����[{?�QW쌲�)<7��`����fb 9��+�a)#�ǲ2A��4�m>(ؠ����9[�y�C��'�� IfvV�3%��J���&�@���v�m�������buEh-FU]�p�9�ǐ�=�����?�����������>��uj�>��.�p�d�7�Gؙ��f�P��r@�Q?���~�y���#����n�-|�b��.^2�`�&}e��V��}�T�0#�ʽ��P0=�,�!��K*�ߪT��̭U�)��!�	��d����xe�u��G㷊��os�Ęc�us�_�[�E>�n�Xd�%��U"<���m�H�y��}:�LM���m��6�������j�����wO������C��g�AZ�d_L�H�G�%3���%R����r�ǺDۺ�Z�Z^#����8t�&4(��v�%����Jmu�v����MGPxz���H2�Z'�bĄ?�_ 	{�}�Y��1E�.g�%j8�3��E؟�:�"��&��� �\���1�
�}a�!e���mu���)CUH}�I�_�v4�r �qt˓���n��k��a�����j����aE8�Xkh\7��l�w��CZ���P/���K�E����<�Ű�~b��4Mz	M��*��/��mfY�Դ��_��b!���'m3��ga߉s�h�	n�t�.4����ˢ��j�,AJb��O<�V�/�{��I��rg��sٺN�Ig��g	G͔8��:�y�~��o�#�`�݄j��=Lz�u��1m�_�й��4���'�iK_��>K��m�F��)ØuQQ����a�*1m�:�M'�����twܚ������$���j��cb�1y�q z��[�E�A(��ly��V�=_EA�	���8F	S0�-�IcF��|&GE�	�o��fuN�45~߸�I���%8����"�	�QKW�u�s$X���Y�M�{$���BZASī*��"�y��T�u#�$W�q���� =v�ͳ��
T *j�����n:;�����\�)�3I�ȭ�!�ɲ�-�5L��%z�R�(��R��|�iѧa�2���.�2#��3lY�,K{��E=�_b��m�	`�j�2\�奒��8y�Q"�p
���L��3+��6�.~v�b�1r�C�_����*Q�
1�^X�m����~�%Ō0�� ��KC�#�(7`w1Vl�/����!�C�h䊕�k�N1�=O���-dS(Kux?��I���"��u��{T�E�B�y�L�i�	��(��~�߲O!$�VǨ���O:���z�G�Q�+T^���"�*B2�#����s$��^"�O�Қ��oj���[}V�AF�!U���T��0^t)eN�N��=^P�5*��\������+���(5����F�2��RT��dp��������:[Y>����wUSZ��)���w�8r�װ 1���������;����+]�"���3�=7��2=�I���:�璐X�VS��V�Be7�Z�+aϒ���I����z.�.�=�����EB��L���
�������8���� ����3�KP |̯�0����)?!�؃h�=���z����L�#�5�0����3��rrn��n2֍w�`!�`B�d�Y8f���MA����=a�㐾1��Li�Z,e�*I����ݠ ]Pn���HjW���*x[��� 	�&]Lz�y�"�,�GB4ѧ���*;`�'v�cbE�"�-�����=���4RJ�}����~<��4�J�1V��k�?6�*�?�#�bP��
hVq�\���Xu�u2��ݡ�{O4�A�{\�^�	<H�2ya���.���ƫ��;'S1���v#��G�qΎ�����m�>+�R�P��*��)��ɶ�z�$�-ڀv��̦�j�	3[h�px��B�9j�ӎ�/
�9n>�G���Spa�E����	�!U+6��|���l۟��[9�������P� M#¤��TFS���*�0���D �����TG0�9i�$w�ख�J~u������p%�f�;�Ӟ��}=�q�_.��a07Fb��:�'�O��X0��$/�\�դ��[���7��p�D�G��=�ן��!��<�H�$��iw�J�QVU)��ł�Qv3��s������񧞡ȥ\g�b��D">X�e$��c�S)��1)�Q������[��Kunj�q������m� �j>:�0�f��^*���� %!T'SIVsmy~��>��W���w�1:��a�πaf�������/�=e�ի���HM�p\���-���>�=�L�}WP0�⊁��쎲��V����&p(��X(	����>�*��.��LwY�E�w#m�I�[��;9�Z�qPvG�]�x�:�"i�4�PIRM.���Sj�M�4�s��qa��>�����e�7ǋژ����=��o[- ]A0�w���)�&;��Z��y�|�T(�Ś�����p ���1ަ #��P���g���x�Ood�b��A�|�B7��[i�|��BA��5�
O��u���xy��
��8k?~'7�u5����s��n���B-1w����ҫ����L�3{��Ky�c��5�W��yѢbp��C�`�Xy*�Np��5��8zc_�������(��g���V5g}�����O�PM��������yע�E˒�����.\�C�^��Jf�o
������{�v�R����Y�r�X����XO�e��K��0�|��q�����8R�����"Z��Q�b�� BI�@����$S��6q��}�LŪ���_��DQ�)q����/h�րu��ܪpI^��
Q��OӰDȲ8�5،,~ʬ��,�V�Ħ<���&�+R��i`$�����S�pk��tNCh�7��>o���p�T�������ӕW@)�mK��a]��r	�@��g�>D}h����v�6��|�隩$�UE�lC��KJ!X3�G���3��}���FƦ(��応-���{aW9S�*Q���xO���l?-a1�[,�j��HD�Q9�S������0h؊�H�A���βJĸoX2���w�c�D5���u��Ih��p=�	�k-�,J:��l�ʪ,���B��{�*f +��O���^� �i��|�)o��4ىy6��y�xkXw!$@�y�s�P���k�$���%�U�JƫһlŬf��C�/�������w�ı�����}�c<g�?�K�R�]1
�k�S���%I�<}ĘV-��vC����("��~9���g�t�P�J7j�(�mK>��"!�O�y�Cbo��������BSû�]�f�p1��S�O���:�
u3t3�M�Ϝ���:0<N�Y�X���\�]&�]rj����_o�=Z�#i�1�W���p�N`1u�U��Y0)��q����1�e2�&,ʋ��k����L�ʨ�b�'P��3dx�D��J�믴��E�p(Y�zt]*�:.��d@SQ��]��- dp]Y�8z=�9+�N��.T��$ug��]��c��6�p��� xy���Τ0�<^,n4���5^��\����Dy�У�,�S#��V�w���O�-����i���;a�{�d�Q�I�4@Pg�1�N�Β��`G[��;ݸ�ѧ�X�7|�������r#�&�������ܦ�����Z �<d�������Y��w�@(�{����HW�&)�}V@�mƅ�SJ���.����H7���";ԥ#i��l��C�R�GeZ�~Zl�.K�}��f���?W=ƨ�B8�4&�(��C��b��Y2�$gV^6���^�AE"fiJ{�[�͏�R���w`�z�" �t ƙ�[j�X�.�k rs��x�d`4:֓��jp�)�^��=�c~�d�<��]j&�T�>�G6 ʰ�cՕ?��\nJƉ�x��#�W�A���L�5��.���nPK�����������d�Al�3���)�-�g�]���=�������)�3ݙ��i�Z침��K�Æd�z��v}�R�W��2�?��x��F���i�tˀZ��5d|�!�[�]B{�p9��.�[�~�VS=��&����ı��fwo��=�Zg���`��O����T/��.���pgy�I����G[ޕ.B�R��Hx��! ���$Xqڊ����Ϊ�X E�(J��c����xs�ٸ���ܕ�D[V�x|���9���In��+����=������q(��m��h���łA����9	B#����d�N��S���8�F�b����G8�>4�K5������c{�T���Xё��{}�UX@�ݭJQ�h��_��}~��q��b���D���r6�f��GsW����$}��a�iI=RcQ�k
l@Ƿ$ܽ�m�m�v�z�܍��l���ǘ��u��������w���~�pN�"?t��QK���`@K� ��0c���B��$O6���5�����Z��ן~��Z��-��V��И�ϛ6}�8�W#�m9$tc|�^ �c�l�L�N�H��gB�$��s���05�]sm��4o��KF��p=]����cd��Ϟ�"�N��y��vE���=կ$&.�&�-*���ɑ�1�J�~L�Z�N���M�ѯj�����1F������`�>|>��":�S��^���� D�k!��?���A2�M��D�gU�|�'�ȶ��UiUQ����hVyz���G�d���e������ppK<��� ���%$.�ќ>�7����y��p�c�G>T�
���:s7*�/1Ȼ��ϝʄ���LVy���8Ӥ ?�.�'��C����&��N L�GC�,P�%:�ZL�y"�C�~+���Z6�Dk�t�߃��w�<O�hE�Z���f}�f�l�����k��^x���VF��qQ����|/.�D�@,+lX)K�[�,��8�q��rq�C�'�%q��%���Z��64��WV�X"��HX&����a;Ǉc�1nfO_���͗h�6X���׹`[V�;���\��k�Ek��	6ބb��]�� 3]9�x�O�S4R2-ŗ�/�
<�J�v������m-�F��ۥ��W���g�x4���iu5�/Je�d�|[�qĞ��Wg�)�7)�4���-tw�ع�9!fq���:A�T��I}�FǿӰ�]B"b�;lm܄����k��є�)Nٰ��
��I�������z�'��,�lv��w�Ң�ұ�j�:�۽���oS�H��S\n3��\���[�r3�B��j-H �8���h��&!��V:Э'���_ҏB�(�c[-$���4��(7jK7y��)>�]Oӷ�NL��=f�ڰ��:����pE������"\�n����!%�1#��l����W��:+�(�Y�ѱX��t�Z)�4�bݦ��y�CQg'�r����q��_Nj	�L=;�ë~��_5^�������2rK�l�}B��j՝>�C�MBbA�֪e\T���,
�Y��@�T�����c7�rE[w� �.`�1�;1��ԁ$\�̷J�HSͧD�����8P�@��`5l�dƒ�2��q�s�\ό}e`ڀ������W���3�W����jD�=�
C��=|A�/.���!��{��(��g�;���(ؙ_%�w �@�Ιc�[��8���ťƧ�m�b������Y����19�F�I�v�����-9Ͻ�'�b#: 5a�2v4΅e�gh���N�w]+RU?^�U�&?Q)���wQP��G�����þ������*�5�T�����X��D/9YD��N����I���Q�K���hd����. ��>:�ޑ�I7�/��m���APA�'������������$9y�ӏ1�����Q� ��J�2f��o�C�P#�@�9�M�Yu��/�ل�>�E�F^��Щ���`Ss{|r�5J(�8n���\��A��<N�nMHX����:t�!ܴa�(]M��,݊���ȹ�v��2��Z�� g���-G�a�Y�=^�B��~����f�����������T$��8y�8�B����t_��*����������$����up�`�_���W�;Qu�����B��~�F{�h^����s�?�� �˭=�&¦��^</�NM#����G��D��{�j2]�~�17������8̅Yb��|QF�U���\s��/钒fdUz�� l����(|+y�d��E{q�J���0�Z�t�Ĵ���E����ck��		Dup�x�{��о�E���[�f19�R�B�"�"g�a�o�5��<"�rW��9 ��_CO�� *�L�J�X�xi��[��5o�5��B�j{OǊ^��(�]��gH�b��S��k,	�A��.>_�l����s/l���'��J���z #��a9�]�����J�DX�3:��K�ӟ(���EA)���IWMsd7���S���� �K��ܗ�MQe�������;��ī��b߀z�U�;%�w@�-��@x������L�,&�/y@��D��?@��ħF����`��iȋ��!�	��������;�,��S,������S�W��~i��u`��yp���h��pǣLB[������z�pӏR_!�n��g��
X("29T�`�JC����&��J����'o�rt�k |E��a|/:�qi<"R\?�*��Ȃ7O��QYp�����F�f��fM��t��R2�ȴ7�dZs �E_lۜ�zY�j��[�]hm��v��͸8�aNB@�D7{��4�^[��2�A����N0G��ԏ��N0 �����d ;~G��*�.�T΍�+�*�^���m6��}�t�͎o��9D,g6�L{b�q�.�P��f�`�>2������!w��@)_\����u�.)�9-'}��A_�q�ޖE���N���S����4�m%�y	�R�z��äW��{ɹ�,T!�E�W�G�C~��ZЙZ;Y���נ�r#c�)�����t�#��'��@�;����!"�L�XS[��D��e��
F/JA���,|Fm�h	Ʒ%�*��7ǵ ��-����N�4���J��LD���jD��ś�9�l@z�W>8E��#sSV6�CHˤ���&�b�ȴ���~��%�:6���| 	�1�g�y��Ǳ����o�Ёƻ�Ý��b,�� 0�����)���<��J[�'�	u�ɟ��)%:ʂ��=#��$�/��(%�-r�{�J�;wE�2�O�0ǎp��u�S9B�4҂��g��v;�O,��7����G4�V�SEi\�0�Ұ�!�7��շ�?��F�e!�"f�|��]T�����#���Mc� ���iz�����.��z�耄�M����$r����ݨ�/�twj�ƹVb\}5L �UC_r�h����Z�k6�_�� �?�W���r��s�v`�>L��{�����[su�,��
E5n�N0�s]��릔K\�V	�4���;%tT%���RKH��$�>Zk�(��z�4�K~�ApM�		YQcR���R��������:�.qV{c�y�9Ϛ��������^�x�E��D��Ck��ڮ���e�״Ϗ`���q8�� \�!?�Z����j�o�[>��n{��'�����~Y��	�Q����s�\Z���@.&�a]�+��穸_�[C�t��{�+kP�@"���dO̵� G6���y�1{m�v�f@��E��oT�2[��
6E�F/�
}�b��;[����_�j�9�Z"?��Yq��8A�,�����`4�[F���Xf&�;|���>n� #��B��{���>���+
���T�?�3��89M�����W�v( ~�Ί�*КWb�A����P+*���R���0�W��o��g�:�) OXV�ڐ�=���꾋��As�Ͱ�+�����ET��j���p^���RtAHV��z-K��{'�Q��t�$�9Tˢt��?G�Y=�������i�6_*�a���Q1�dʝX������D����Ty�u+���d�;X�b� tƍ��ϰ�71��E�]K'�%Q��SH�����A�0�Y;����s3Nwv>�_��Q��1?���&{�`�+��e�e$��D��+'�f��QP�"D���"uL �{�RL���џ�&A.��l$eA������*�3��}v��j�.Up/!��б���p�c�䏊Z���g~����ndqG����KQ� �w��r�I�W�y��������$����!4<5�
��H�Ù�u)���	٠)l���Ӫ~�y�B܌Lq���V�2ӄ��%�ك=�+i���X�@�4m�n���Y�yy?�{���bn����Ac�r�ۖ�{�u>ԊÌ� ���6y".��!���������T��߉�.wS���8�w!Ȩ`�Z^F�p���Z��o�y��V�C�#fƅ��=)3.��Pܭi;���4G�<�!�@u;,JK e�ƴ�c���h��Ҽ�vf٘�1a�G���U�y�
*I*um��x9nQ�Dr�D~[��(�����y����&�(��k�>�z�_7�oMT��_bh��/�*�yG-�2ۊ�n{RBoj��)�N��
r��)�{$N�6:���@mz�!Q���,4�L37-�؟%6(O#�/5q���a���֑��>4�`v$?n�B	+s�K��`�ϞR��j��_�1 �֑�%Ux;�ɗ\^���BD'��d^�[%������Wf��T@�R� Ef%�)\]��q6uQ�xK1�Q�͹� �U�VO����CYa�vW��JJ:4Ŏ�0�������U��G�z��m֓l�BOþx;�[�]{<�I��KDP"O�5��%�?��nmp�����Y[�U��e���Y?vC�e?4>!�ɍr���2-��[�4���ض��g�k�~0Y&0s}�ͮ�O������
�Z9>uU�L�C 3����	@+��G%ԍGS�<���W	�k��a[(��ӣ��a�`tue�Fy�$�g{��ތ)�8aj<ҽ���\��8�k���Y ��O9��|������
���G&Tt�Kt3�?�̹\<qu�Rz-�֯�F��|?b�ѳT��F�>L�_����-�1����p?�Ͽo����+£��Z�Bob�Ƶ�)�����l��Ax�R�ۦ�ؑE�	)��M!�LYCy�Օ�k�b�ҩ*����\�R��ـ�u���T+�˵��][G"�ِd��K�4�<���f��w�
�F�ہ���l�y���(��W[��N	U_(�,�ZPQ 3p*A6(C��	1V�'��SF�[d����&�����W6��U	/�jPhJ^��H���c?����-�AF�?��5B�=M������^neS���d]���Z�k��|�1����\O�����`[���e�+���r�a�E��q��y��m �SD[��$7J���������P��<�j�%��uO���B~\����d��7⽧B���D�X2�i�.��4����o>���e��0^o���E�ݻ���]�q�N��,IFWG�fv�+A�X"?j��f��M�d���r�.�MLv����[��	�F̋EIaꛂ��3��6l��3�%�v���V<Z9d�鞯�=@�B!���qX��0�y���`F2�����藏23�{�;�S�k�s��?"m$<��W���Jad�ޠe���\�s����j��Ebz��9-���=��o��k��x��6CU2
t��zq�B!�(�Һ<jD/�x�0Ec�=�%nF4G �#���j`�`�Ȣ�R���%e������X{V�/{=�;L��Ω��� 50�B!��c�X��9�nLp&������t���ж��$��h����0I\T&�| ������)8��<Q�dSL��{�|��A���������w�j}����-�X+���v��C7�|`����Z[W�(�����[PҀ_�;d�q�1�`WT}%m�uKJ� ŋ�־�M�Vڨ�[��|����*�;Y���ZB����N�_�}K_/�Ѵ�U���~��*�m�f��F"�D6<�o胶<�j^�w9�c_�=�4�ey
��+�\���6sZ?�æya/x1;��N-�#�kA4�yh�`1���ò�v�1�m�fk<æ�Mm��P��zjڕ�],p�����[�/m�J���V��`t���(/.�ǃ`�4.w�{����9�҄ �`$ �[���M��5��
On	|�A����h�l�ԁ��I��<��֗���VPaНO�Ҡ����88+#�b��������czu����q}�S�x#���޽�T�z�zE��	\UI�F\�׃U[nt�=L�AK�B�[��I��r�H����~I����1(��0�\7�����[��A�lr�TR[;a���
��:$�Hz�-��0n���n���5B�vp��%-F�h6��=k��8�^�]��y��/k�KP�l-�ސ쓒�H��$!�@o�n�"`R�Noy8t�T��쇛ȹ5�7�w�z�Ė���&؄��4����#[��
1Wv_L���L|�X��	���_ȕO:���^��/�w�g�^��{�>qGb3kn���Du3Oe�$a�(���0	����' ��s蚯XuW��6�o�5��2Q��"eL�t�X��,��&4f<E۞�8+��,0�`�*��i=E�qO�7���~r��i�n�?g6Iݲnȟ��.���A
?�����@-e�^��֭s��Ur���%�{(�{�EYy�;�ÈBV�9�7x�j���zt�+����\E۹pǨ�Z'f�r�z;�5�]�S�y���̗Yn�nYq-g�ӿw+d�-qR���l)ǳ>�G����*��?Z�܂������wJE_Jh ��|���m�H�Jѓ�a<��1σ3�z�쓴Ȋ�UM����|F�>q��(i�(K���
'O�[][W���G�u��eWv�v3�e\)�x2X�Z�Ն�W���(�
)@��P����qXww	S3mjW|�,=tbѾ�1�����G��l8D�>,�*��( �v����J&[nx����;<�]RA@�u��i΁��h���}��)��̀l��%���(���S���E1�oU�j5�1�"x�=��_[v꿼Ѻ��V��ׇ���TM� 3������� <��m=W�fہMWľ�@��4ekD�<d��� �j�����P� 1>��!Y�/���/�Guԝ��ПXDrx��&�WZ�IOֱ��r#�����}6q��0*�������oB8o��Dƪ�yi�ח�LB�=� �r���)���K�I��9.�6��1�,�M*����+'��S��lꛎg�l�<S��W{�`�#FSK���
�N�Ŀ��J�#���N�CC�.��W���ܥk��K�ҝ��z.���=�=��L��{�iFU��ʍ����=){-ɾVx_W"�9U|=�+��br�n�(yVb��z�n�i�ǫ��y�DD�Yj�no"�%�O�w.��󕅴����6 X�tv0n�����N��=?�s�3�9C���P������߉8�|x��;����J���'P�rK0��`+�!��R��%KF�H;�}�%,m�&���(kj�i�wZ������5�FH�[�%SJ��spܲHH~�}� s��,ɥ]N��vq ����V�̜���w<|G��_�5�i HXu|%P�.�By�_�� ��8���-�>����o8�X�
�t[Y3߾8r�V������/9CkA>���f��|�:(L��KY��fqjZ�.�k+M_;��ɰG�����Z:����=	-Q�A��@�b�yr2tc��c܃O��q��"��0R�����	�n�	��!�p-�p�9�����z:m}�h2�)ӈ�p�%F�!��>���~3!��s����2x�j���D�Z���+�Y���\$�o)��������,��š� �PYUJW'���ȴ����|T9�I ;����WN^]4GF���z��.�>>�H�/'mX�Im��D��pd"�"E���ǲT	�V�;l���iS�O$w�<𓡰 p�)���T�ڦ�p�s�O�c���I#�(w�w�
�{�^7�Z���0��-���3���E�Է_Zv��b���!����i懷B�7x��W��j��v[�\хO]PT�2�go��Z�?̜*�Ww����	o�Wm�Vs��Ú�Bϝ��[S��2A�4�L��`'t"��X_�ȕ��~�[SQ#�wB~�ck��!��a�<�)�U+j_Q�Ƨ�e&uRp�W����cI�вK~\ֻ�_b��!�������t��>�m��4Ίw6� iXP.�����+G�M"�m�מ~�}Y�T���C���O3Ci�}���Р>p���6ц���� �_���A����e�5��w��pRŪ��G����]<���Cߦ͒g��*���b�t��ޢ4>���@���ʉ�9�I(PuqH�G9Y,x�7M�\��1}G��$�߭�{V$�M�ˇ窩�\��\k���bz@�,&ZI�IV���"�hH���;8^��p���+z@�O<(���H�I��Z����[s��P3�F)0w��D�+���)���<�Wr��,n�)D\�8:xx)����WI�T�>�I;����u\[��<�H�Ĉ"`�6a�:��v�ByQG��^a$��Be�p�e���n�Z{�3~=����y��<�7�V=/�\B��gߍD������ �S��P�gxM�{�?�6+�۹��-��}���]u��3��<$��d*��Mi��*���$"��9��?Т�<7!wq�Ø�S�//�Γf'$�-LC��w�f��w�,&�3}k�e���F1�?�h��bhZ��K����C0]�} ���q�t`L�FH��'����X����Ł�٣�����O�pڥ��%L��3�:&��-�w=J�c��F�aS�ʴ����O�7K��U~�
���!�������$��	P��ܯ�|�u�B����=2���n�^>��%D{�!���0;�x9mp��#Ac�b'��ԻJ�rNUx�9��ẗWCk� �Lj�g���k㊥�o��6v���nf�8��H� �%6���'��Yl^DAv;���K�?`]�KܒRcv 7��p�8 <]L�q����x���v���e�)��&�Y����8 �)>u�'����.�yv]Sya��$Yh/C�߹�m��w/�Yasa�w�qL��σ�VJ�����VQ���O**�Q��_����	�M�wa��h�(}t-x��G�xw�C����{]m��BqU�HT��|��IƂ����Hl�0��@�'�$��vR��3���=G6m0�h�/��hl%#
D���`s�d�sq4!�ي*������֜����U���	ɒu�<�A��)$y����숡���F�s)����yH��T�Jh�6ÌP�k��x���ou$,��}��9�C���M�������/���scIεi��w��E��l����%t�ç�'�)���j�>��������g�|3n�G��/l$b��%$�#Sd��P�+��&2T~yf"o�s�t��X��}�ܙ��=��L�}Ն�ft���>W "P��"`w$P��'�cS:��#�q�x�ڪ���}o<�P'м��P�d�Y����Q>���E��=<$�����6#��gz�qc�"k����������7f��w�ȳ6+�i��ih��{v
I�h��#Vq1��!��Y�+�A��`5|����K�ň��\��}_�N�&ݶ ��\^%���W�Sh�������k[���d�˦zOe;_�c��������⨜�R'�P��V�7�y��%y"��;S.]k�ݙw;��JK"g���X鴮�򕁨o})����-���N�.�:Ϻ��S\g�d�r�Z��Z!�$�w�Ѩ�{�)�0�uP�m#���wt('�X�F���^O��(�u���A�Y��K��wV�\nΙb��C�q�.�q���%(�>5�O��KS��vT�����Z���J7;�������K��w����O�r�=���i�3~ޔf�w7V�u��>G O1H5]��퍑�(G� M�������إm�R�:��pz�^e����FǛ� ������f��w���	|��Y�������aݲƉF;O@s7���\�
t�dG�V$��b�X���P_�J�C���c�݋[{X$�4ἃ�|}�UI��s���B�N*��3���>�R����@�Z*}5KB�f���`��fj��`�ƃٞӇ�T�C��]�ϣn�L�L1�NHĦ��8��%,Wl��fP2I��P��Կ�����{�쳋���t��2?��_�S}���yiR�r�ƾX�S���[��&��ߢ�����l�d}2�����Ҽ�U�]��6�\/xkrJS����b���,�{����M6��	"��bc�+Z3������$�l�{?��� F	ydP���8$M��u]v͕��d�v�u˹�I��\���3N���j��O�,�=�\��f/�U��sJ�՟�X��g;VW#Om�rd@Q�Aݡنb��Z�^��ӂ͌V��rm�'2�d� T�I)z��bd�2����j��G���x ��;��#��Tv7�B���B����==N�	Nt�ו��� o/ϖi��+���ᶥ�j�ž`��/dH�sY���Iڃ+/�Q�X��5�|�o�9�2��7i�:q��Jm�u��8��d�c�GA�[���>n_x�/1�hfL�X�M8{��
�ż['B[��~��"/�ɴ�Iw|�)I$}���K�
i�KuwB9!�-Rv� 1�f�Y�Bs��]��)h��i�4��\~Wq��T�nǮ4l[W_e�R�,�)���L���T����.C���Cl�y��c?$�u�ΰʾ�4��q,�y� ���I���U�n�֧���l�6��N.�i����u�_��"����Ea��
�G��x��#�Io\i�U�I�U@�g��Ǉ!�r�.{s���b�L������c�uk���C���L�|�$�zѺ�VB,i"̓��+h���a�,�عh̠Y_q>���
^�%�5�?��zw��F�D���5�|ϭu@�����[C��z�Bƚ?G�	ñ�|f���'�:�@�R���<R*����@�0m/�t�ͨ�&O���k;��\�G��+��=G��\큽��C����ZM�����$���b�h�:�Z��5�����9:�B����,�ِ���,! У�ކl�z˂��7p�R�8�C����p̐����џq��_(Z|���*��������sugF�'׮�����_\�̻N�]� ��[+�h�U>LpT��D�\��G1�L�pd�<h�֙�R���@ ����6*@�Pb%�H�[�Sp�wX���ӿh���SȀW�m�AP|H��~��e?K���_�Ȟ��#��E>_h�_�`�d�2MҀ!i̝r5�
�DH�|n��R�#�P�Mc_"1�з���ސ�i�PTv_���w�j�CY����o�;ȇSPt���ߜ@9SE�#������;�P
P����eɴ:{g����������b��~�a蒴�!�3i��GFvFD.o{#u4d�B̕R�5���T�\�/�����]=�`1�0j�/���g��6�u�[��f����#��;���@Ρ2�k��3h~��s�fF��6��#��X�xB0�̦��{��l\E���`-��o��������J�U�ڙ�6��Tv-���'�����=����+ԧ�o��X)	���vdd]�73����ZDG\�ۺDM��=��S'�K<X�aݠ2���7̣Fc+3p�������..�Nd&٠��Ը�UI[��,R��R?�!�7����e�p[w1�[ȞƦ�D,_��!+F���[���E�/]m�%ь�V��{h)�s��nC�+�}�u�4aI<O^�@ԡ#
0� �t�E����03`�CL]��o$�I���U$�V��9�w��%&{hJok��cx�*���o�nAV�B3������+�JaR�R��:G����|#�HxG��?��i��I��m��n��[��;ҤNQi�T�b�;<�sB<�a�r5XT�/
�!��,��ã�Sxgڪp��iՃB���� bC����{p�h>a+ح���1q�d�C���QW߾��t��d���e�������|T#A����I��Ucʋ�	�θ7�$Ӏ�����?r�3���8���t1 +ޖ�NmY�*n�@6ðh��\����/a(v�o�r:�,��+�h�9`����p�@*{��h�";��t�^C�>���>���/���\�ۦi���Rw8�e���(�GLݎAm����W/�G���r�K��~.����j�� CN�`��:N�3�j���g���F��1�����AJ�V�;�����;�{��l�P�t^c�R� BIiV�*|-z�4���/��|ܸ},v�>��?{�㖴9=��M�ߨo�N��e�zP��L��b�md*`���j�W�&I��Þ�ţ�"�~�"�� ���Ke#v.]L�f�$��M;��q��(�tӈ�?��&R���~,�ǋ]3��d8e��w�ئ�#�ᖩ�r��ɦ�n�s�T�
���C˭��U���ʩ)��+���+�͠�[�JG�J����=�m)DY'V`��T�L���L��Ƙ?��>�s���,JY�GEs�(83�a�i�N(c��*�>���L\E��q��;����V[Ӿ]ꦣW�
 �edeQ$����8�~�"֞��;�=&��v����q�׸Լ�U����;����M��&Lƙ�+�t@)K����9_�#%Q#6�x�S�)Ү��<��R'�
������i�U'{������&E"\M6��{��?ۏ��f���Z!��1f���U-m)����'iުeb�h�9S�4��
r�rv׵�yq��q}���ڒd7�֝��'�*�Tԭ '��^�\�̮M���4�󒥉��"tHcE��Oo񩍩[4Uj8�j¿�wt�`M�в�+���Ӯ��^-`(	X|F�t�g�@�2���t|Xd@���_C�Ha&ڧ�!YDО(�ݦ�n��:Ó8�g ����t>ihݟ��֚&-�Ȇ��_�A�廦qO����qd%l�S�ƽ�.|�w\7��?Z�`�}�U@�~>p<�̧d���Ɇ���6Q��k-�3���~����Г��AɦKKP֨ӶZ��)z��:�<� ��2���	+��#g�h�T7 ����D�+���O�J`{r�r�2���x�Ӹ�Xl�􄹈b�����(��a�%QX�b�09u�Zu9_�C���Z~�$�e�d����\a�BՎ=��C�\��N�n���U�yq�4&�&���+���BE9�,�K�b�?��:�wO�a<`��^w�`����;�/���+���r������w�����c�srG���p�z��/r�[_��e����
�n<tTo۳�=�?NDl�
r�d����>m�m���[����+t)a"���ٚG�s��籘"GHD�� g �8}�ѥ�A7�&�ⲷ�aW�^��]����*r�,n����;�gt�h��(��=���U�>�g7m'o���T�O��l� ��bHW�e�v�W��9����=�9O���h̉�'�M�&�¹kgrz�u���RPԵp�b ���S��%�2�˙^>���y�Ó�J�����B�k���:�@,'�Q2�%�.�K�ء��F��0$vdo�b�S;-�Ն���m7q�m>�_�M��e��l�2R sr���!��&�!�����#�_)�p���SZ����'��(h���Ѯ�{?��]�?����O�Tj�;gڄdz#
3�D�ʾy�P���D����r{�0x...��ՊU���=�8m��%#�s���X�=m�֠V��f�����O����o
z�E��+LѷJ.0d]���cIO=�M	����]�D���1�^�ɝc�F��n����"̚<�)!�~
@	��}��W�Y��r1pJ�� ���F���AN�]G��.Y�
���)���&��䐯���B�6� �
������Wx3�ו�IE���g:�|q�>E�����z5j�<���Ss�=(�ŗ��RЕA�A�pma,��|��/0���~͗/�@��BR>vj� ��n�x�j���|��!��	4�	��U���J�ㅫQtR��N���ߛ�W��I-|2��"�ԧ�	��2��x4fF��\�RNLLմc�Ŋ\�|��d��x�"��U��;rF��EE��o��%5�<H�� ����C�������AN{�K�vl�行)l������
��HV�wmb��:�\z*U�fV<���^<)^� yu!lm!a4�&��1@>��zET���m���d���T���@��T��;+C[I���^&-�2<��0u�\;P*���=.y~��2'��=}���Zm��%��N�ēM��`�Ui�6��	T��s�ϗ\1qi`=�)�zԐ��¸�(L�����W8l'���D%�Y�&x�#�Q"G��Cac8Ӡȏ�8�:,�E 0np]_L^uŏ�!��J��~���iW��$F�V��@�e���v=Q�:�}�mG�h���'KM�"~���:\�ʫ�G��25�	[��S�ر`�jsO���P�o�U��@"o6����I=���Mn����NCk�\`<=���| 6.q�V
��/��1S��ȷ#T��6Z9���p�xp�W�$Y�p�z���D����O�G4�pf�`oY���o��3qэEP|$���o�Y/���%E��@�q�U��"���˻Q� 2��)z_mpq�2�Kˌ�_VK`9s�� �_�����75E�~*ڬ�[bU#��Sn���$P�} � Q��$( [�0�L%�J�W��"�8XWKS��0]-?�L��倆7v�#��[)�]�_D�0�- �8t���F�Oi�>�&��"�NU�U1�%�)�ȱ��IW�Y1�u��n��3$�0F���RI�#i���V8�7�w[�OC�X��5�m�^�!���J�U��2K֝xrf��rA�OI��Nxj:D���o�_9P�>��e���:���/,w,q�;��c�����i���YE����V�9eO�h�@��
d.�T����>�޸���lf�b��-�0jV�ϐG�����r]_���x��t�F��IzA������ZRom�D p�g��̈�+��ߞ��p�k��I:�������Z�rDd�����b(Uڪ|u(�Ѷ�¦��������-��Rb�ebf����S_=І��N�ñ ?���Fp�}x����{~��`�JG������[�5�Cn-�f��#�X�t�����+s�&0.�v7���d���Cc(����(���iE�1���Q��rF��]φ_�^��J�̪����*����A���۸��3�^�׈)�S�2�kIwξ}���MG-d��T*�E���绞��R{�R�axP�Y&o�^�˹;��ٶi�=�k�.??�d��.X#�{/��8%�`7�_��_#N)�����>��cCt	��A�$ҠW�	�v]��
����K����=[�LhF@�Z8_v�Ar�/c�X,��֖�*���!_�9�{+�����4r�R�����;���6OGb�13k]���U��zRit~���Iߔ��M�K'��o��PB�CK��UL_`�����f�j#�@E��TUԦ�C}�2�o�K�U��k)�
��ǜ~�W�9��fjYh���)>
XcR5;�~)�$.�:�/�����a����[��ǔ�^�;������f$��m�_ڞ�!f��*
�Y��-s*)��OӳZ�Hk7/��j�م��ycq�X�<��)
pТ�i�N����c�pnm��S�W	�4��޴��m
��|*?k��NvĖXb&�ߖ�+��i�Fۑ<�t�Ư ac����<S��tyN��i�$�ʓ�\�T�>�Jn���Z j�>+}�?���0�RK���w�J��W�d�7� X�NO\�<-�;�U��7��NKX)q'�cŶab<��$�#�zW�{".	@&�_<�2�6�|���z4Ryo6�v�X#�N�eĘ&�w�_@\��Hxc������?3�x�y�Y��B0a��B˩�}Wf�=/�q���_�(�B����a�T��ADr𠜚{�d��嚶�r/�8����Œ���k�R�׫oY/�'u�w|z�Jmm�<��4�!ס�׹%�M��oW�h�޹9DJ��:�f�	oe����7&-� .���-%�t�������$�*��4���EF�9M�Y6T�ӝ������a4���Y �#B6��9h��k��G;�©�۵�����O�����7���# ����%S�W�sg�����w�A��{)R�B"�6��flW4�^}/��i����A�. ���ω�J�<��G���mV�:9^m�֙߯n= ��a�t�@�%��rW�Ɍl�e��9N�p���� ��-xU��o,�:2�C��2~>yg�����z���Q��	I�ͱ�qF�a�ѲF����VOz�F5�=jؿl;�)��@��,㊡u=�QX�@��$gpJ�5�G��(�>R�R���$ P1��9F8gm��\=��W���/oLo��dZ�cx�R' hL�S,V<����/
������+�wN�Kb3c�Q-�
%
�|Z���X8d:��������:�e5k+�H�?��!2��캓��퀛�\�Ǵ�JV�w�-����{*�@����]�Yӂ�>X���X<(��R�����;�!��:B�_��D�䠨f����DBK��qٮU�葢�n��z͞�G&����&�a�k��I� ?���̯�����E�,]ܠ���q�Yص�ğ�NRd�� �$�u�1����d~�~�lF����pp�Hwl��.!���Ez/��<�S��P��d��VS�!���N�(�H  ������-���nֆ˔9�26�#y�ɟ��W��4�HpY>�|K.a�aH�b�uq��?�֠�X�n	������2˸X� ��Y�W<V��H�l:wL�c��Gܬq���R��Vq�;p&˃��w�u��S��DDD\gIr�u�NR��5�\{X���3TM��d�`�?�����$�!� �(U���?�����8I�)��O�H�`����f SY����P���YϘ*o���'sH9���ي����Q��#�nx��/.������2�c�F���[5�#!f���[AmƏ���5'+���Z��?̡/�*B�tD� K�N	uBΰAP,���$���qk��x����q��j�8yx�q:4aM@*B���&����m�b���Ͷm�{��.f�S7G̼��u�IrFg%+1���?ۼ���굿@�.�4]&�Y��~Mw0yj��ܟ�D~�M��V$�Y�oEo
ic*�p��%Fa�͞��[
�b�t�~	�d�����/y޺����ń�%>���8Ta�e���G�3��	��QвXኖc��xR����e�6^���"
�2
�(�K!���&�/Yk��V�F�<���ݘ]��a��|=�]�i�%;GL.�%Q[�YT9k�sz@��Q�t*�g�EՐ ,O&�b�W���w6�L�����^���~����3(#�O���0)I�,�vE�Jx�\i��s�
�9����Zg7�v�ۑ��y�����.ams��yQ6�� ?g�f���T���:;���������e�h9O��0_z�
[\q#oF��'%X�d ��Dg�t&3S�Pzh:$r��0��*~΄���a�v_�-�њd�?b�=yY����H��h,j
�K������_9�9�c�Z�g��$�#خ˕���Ke�q�lG�� ���9�3��4��Ǻ۾��P����Չ̵w)���R]���m@ک�<����a���J��������}O�^��?:���{C`��wۓ%[U�9��iB�ݓ��H�E�x8^��
�������6j�?ܝ4������d�xD���=�N`��Gi+���!�2�yk�DlA!X?��)�8}#�p�T�rھ��Kihӑ���5�6���Z⃁jĐ:za(�Dv�r�tS��;S�I!ӑ{����"RR��%!���:}�H��fug����&�v���^M7�(_�_�&l_�!�4�|����ّ_�)/�g��2��� A�?��?�fA~d�$,,_�(�"y�������%��Lᑸ�ǲ�r6W�zw�'�Dx%7>.��uN;G��jW*�}̃wG�_��ZX'��3 �b���Q#�b%5뚎�3Ə���frK.�fn���@�%��{��|)Й�Y�N9-H1̦�f�*~<�[� �a��������{p�/�v��W�����x�h3�>?�
��h�N6��^����di�ʋ���8��x�@X�= Y�+�[�]R��o!^��a�������&A�w��[)���� ]�w�	��^���/t��0�~���Z�m\���H��eyr*D�;�c�yy��
-��B�Pר���ϫ̀���9����߉���Q�D����F�x,����.&]7.t9����>�n6���3f\'�4�
ߩW�^�� Q��)�Y&�34����A�yKxp^2T5�f�7�8���]۝?*��&��~��[�f�¥b�F��K��n�	k`X��C$�FANv!���iE;�D+ON�6iDA3���k�#���a[�&�v�B)׵R�@�Ô������\���;qg�����Z~�UVs��D)����〚x�M6|������8f��7����'����+��@�Xx��	��07s)���f�,?����S*����W�W�ư�cL������q1��R���(��dLF7R��ؤ���a���d K����5��0@Ҋ���BI^�k|nw���c/�!�_��A�)�M��B����q���c�qEH��VX�h��hZ ��Ь(m깒z�%�c������I�{̧q�Gi$�=���Y��H�#z�E���Ac9��� i5�5M?����qC��#��H<������� hE�'+r����פ��]�nQ�i!�l�n��t��;�����D�)�z�������-��(���6Fq6R�6p�z�ˎ�:;���!%<�xO�不8Pֲ,#s.���8��/9�掮}��M.Ӿ���lP�)̚S�&dy��q-ʑ�g���x2�%�[�I�j��A��{��W��e�5��«� �'�k��ICu�����j��F���5�� �y�Wܓ���bSF��7�Ä	��Ɵ�>�'Â�\x���
*
�o;n�=��P�A��5�'\�������}B�"��+b�	}�P� "Б؄�՟Y�qUIbl"\�+ �����-�����'Eou�g�C��C���G�v�YV�^iwXZ��L����7b;
�.�E���uS�xm9���_u��<�d�)��� t ��t���)U��ygBN��0�O��.�����>��M:w�*�MD�Laݾ��RI�����[�w����p��ߡ����K�S.��8Z-���H���Nź#�,Kt%~%"e�q؆[�y��܂*^�k�iI��.}��z�Y���l���"����E�y�Ԩ.�����NM��V���l*�b�.�`S��YJ���kT�+���i1�.�7̣�5�F��'ۥE� m��M�V[J%�/r�ǉ�V�}�n�+�����~1|L6 ��r���40N�!F�	�_�N���ӟ�C�<���E_� q80���O���-��������4�ƤF�B˘�Q�F!z���O0'	�R茢�9l^?zLF���e<㧽qc ^L��{dt�Dy6���MWb�e�(�4���Z��2�~ �)L���E0��꓏��P�z�wܮ�T����N�
����g�Ԙ�:���I
),Wν��4��V"ˑ�N6��+�.�>�Q�c��<Z�ò�P���'�����"vrQ��-�!]|W�B�e�[I=&�`@��_��N�s�o�NZnK���P;y��H��<��O�R� A��u��s<vKm�w���.*��ɻB���|z����QX{�k7{����N�y�YƗԀ�jC�����Uj7Ay��}�����)���c�d�Sƚ�ZSƽ�0B$1�ɭGdz���<��j
ܟ��-᎞�T�'Fϝ|?�#�{���T^�l��r� )��<<�<v�� ��t(�mb��2+��k���;^ݍ��ĉ�Y.��$fn����H��g2� ��_�g̅l����9�BdpWYngz� !�	4������kp?�a<�A��hq��$��T�`�k�����x��~1�����Ԭ����ae[
����k�\S�:��c$�"�C"яh]Ũ�u��N"C��gKg��J�12ߗ85$Ͽ� �k@�D���z��)��c�5�Zxl4�c��f�	\�=���J�H������}�U�cv��RyÈ�����zB�r�w8$9&��9@��3S�M)�� D�7���r.�>-'i�4����X��v�94k���5Y���"���<ى�2cϘ���)21�����ګ�u ��b�R��m'�6� _����ҿJ"�����i5#�H�;p�[�:j�)�J�}�h/͑�J��1T@�W.���J?(���Sޙ�7�@�*@32g��Ĕ�L���;J^��UQWۤ�+��W����b$���-6��&�:��L�Rg��鲍iA;K�f7p� ���װ�Qqa�����<
��O�)V����c�a��eO�T�Q����*�g]C����H*��w�RO�Қ����J���V��M�^�>�$�N�c�CV'� [�ü���+v�)%�D�q{ sr��:|*p���H��9�Y��n�>gw���7n�J��Ɍ3��0��Bݹ��z�1��I�ߞ�V^{��ζ�I���c�����g��$�`��f���Z+H����@IZ�ih\2g�U��V�zx�=k���<n�����;�+�\�T��:-�܉4q�Q��=�鞦 /����Ka:�n*��L��Im>G���o���-���s�~��9~�L�q�\*BP�^֙#� PҺ� Nd@�Е��|�!���P�b�;$Cw^�#�/�°7'��Gl��{<W4��[,Pr>�3���؎���K�k�Q��ʊʇbZ9�vZg�i�=l6��9��0J������4�Ji6M��'�����.Wk��t�R���6�.���*L�8��6��P����~��ߺz�[�EZ'J3ߒܓ�8_	�N3[�Ҏ��l�~K-d95��+i@�������2���b�&@]��b@Ne{Q�p;��*�BǠ�t��4�轸<]5}�Y���y�A�Al��w 8�Tby�z�jS�4��lӌ�~��6bs#5J��N#�+_��P�__����0����Q�1�Y�,�{�b�89���WN
��P��!�l�+CC?�����>���g��� �Lx;gѳ è0X��Bw���+��g�A�E�a��,]�K�e~�`y��%�ɮ�p�>p��Bw1b�Vr�2���2L�򽶟 ��I��D�*n녙챧rYB�!�`D�])�r�=2�)n�`��r���u{�2����U�)�\�����atxK�A��3���/��d�~�H�KM���[u��w�@6'� '�u���XjeR�8�e�A-ι7>�ϲ�aK�L N!9�����kԴ��p7��ݦ��l��峥����g�_����8�L9#k{�J`�ι�V}Y�"�����Q����R��S��<RZ�}{p�!wDWk]���Z�/3����	��s^w��5yU��`�]KM�����&D���xuK��=��%k
IG}��$у�A��m�J��;0�A� �QDw��1r?x��0�B5ah\"$��aR
N���;+$�J�-��I/��z��PE��\�G��Z�IM����{�g��1�I��[0�p9U�:�ǻ�`��E;��g �"��>[�=~]Ft�z`%xHRp���_0�qnJ�[���L*$�H�q�*>toe���]D�l��`��M��|Mûg@�����v<�]R���	���6���b�G$Ə�`jǂran���}�'��7����Ìc�%H�o�N-I��qkW�G浠�޸gYi��Uy�s����M��E��\C��:UC)!�ތ��a��n�2ɵ����᡺�.ݖ3Q�r��n#��@#�������aw�f����q��1������xMα!���h����T	�Kn��H6׋:�XL�es��;E�����eio2P�	?�k%����Ɉ|�����UC�*�����_6�#:��ŵ'GP���@��|�w��Wˌ^�@�̌������[�Wΐ�!�KLUP�4�4J�Ԩ�|o'�.޽�����]��)]y�Z��[�b�3&��7���@%�fB[YR���Τ&$]�߸}v�߄��t7,�Zz|wh���	���<�|���yj�Қ�Q�Y:V��zsM6��ѴK��g��4Ax>\���߁��B$W4��$��J�V1J�x>��O�4&p��ԋ�7�����V ���P�f�v}0����C|�c�s��Gk�Hg�Ж�P]"�\+�J��eTd鮅!�����l�#M�n�~�{p&g.}�p��+�sZ#���$8)M���Nj���p1���~]sl�XxM���`�PƸ���-w�)� ?P	����n���4��N��L������p�8��ԭG���8w��h!;]�T�*#���ڍK2=pG�
@	�~�n��M؟�ܷ�#p[�m�, h��3��K�O
�~@�}&�$���hu���W�v���g�唊yܳנ��#�n�a�FL���b�,�,ܨ &��{�>�t����n���3�2Q�baK#���R�$� 5��}}��%)����Ab��<�����ݘ����o�� �"_��{���������Qq��Б����/��xS�1ً�z�&/��4��4}%�͓����Bz�ù��~d��,���7M���Q�G�ޔ���(�M���t�ߢ�>oUG�=�#ˁ\�If<����q�Bo�Jܛ4���!R F�=�l2W��n��
��s��\�4��,�/�@Ԃ%+��⁸x���b=	��v�2ѩv*5C=��S�i˶�&�4ŕ�f-�Ҿ5-}E�~SMSK�\�+���V����(���H	n�߾�Z���I�+pF����Z�",����H�Q�ڬ�ar]LI�Ol��0p[R���<�[����F{��jRy�<IN��9���zq��>ܷ�P�㥥/������A���q�Ix
^b��� w8��g~!z��z�:~E�*:���9�T%;cfJ�4����9�*��O�/��@�߈�����Z���,��0��v-�ͼIT}g�e��
o����& ���\9����*�X�ƤTna��B��v;�l��x/G���ɽ;��$j�υ�$�ı��X����CZ�,�*uE2~nГyԖ<�=���LQ����]����ꂁ�e;�wW4�e3���W�����s�h�q�cF�ݾcD����?i�f�LRz�����+-���\����V0��a�
A�u��xnQ�M�~�JxA��\W)����\�#�Jy����@uA���ݽ�b5��E1���G��_��h+���4�;�"p �g��a&(�pi"�û�����c/��_�9�W~�xa]��8=��+7k8��X<Q�*�'s��`����z(�E���q�yu(ӕ��IX_~���%6���F�*'�����s�sV�o>�W���m�FA���u<U��]k��<f�G;V���IZ��0D66>6���QQA�1��lM�}�ojEp��ע�<�³�>����4�Rȥ�1�H:�F�i+�E(�?v�*̓Z��<�������� �T���c�0�G��]�$�� "�Jq!����z��B����!|�Oㅷ>Ң��==��	/յ
4��@I�Ne��g$T��a2�^><�_�ۋ~?�LS�1�)[]4a�L﹏:q�*i!+�׺NX���#�*L&ê�M%���~1Hd�Z��m�/U�n��Eo�(>#ܻ7[�mY��̝ ֶ���1p���v�
�iq(�>��j�9�g�'Wp�����}�!��)���<K���K2���+`+5ώ�7fE����{��brXR]M��5��*�Z-)Q���:���x����~�Y6���-��\�]O�w�'�k&��n����'_��xyfja�.k��ɧ��<�٘>w@i��O\����hu`��?����Sw��~��@U��s/��ۦ�u��E��5`��e�,����MaJD���b����U�c��o�d?����Q3�*
�H�/��D�PP�y���,_'��dk]��R q�[-���И��*��(=��ȳ��2���'C�jUY�X�B>���j�wg��.ܦ��-� ����$��oRX6��b�,$od�~$�}���i�^�Sj��>,)�7�s�bk����U�8lHJK^�#kW�0K�e��tw2s~۽�us>E6����7�aj� 6�g�7�_	,R�P�Э�e�~�u�ԦA����mB�5���"!&((v����UF ��\w����~rR�eo;�������J�2�5��J �I<6F��;��p$�����ы���ꇈ��n���H͇���*zO���o �������_*�&f}m��H�����R�w� �;�"�n�N�A����
���kW�Iζ��J}�ؓc�Ѽ2��5ʸ}��Ia�U��/ڈO.�[:�u�"��m�����ܙ��㇉]@�q	޺7N��{��h�ƕ}vT�ݰŮ��Q'��n���d^�ȡ3�W�zg�2%�G�̻��ޥ���X �yӍ�R����:`�\����9�щV'�͛��c�aLkI��I�t��4!�R
�(�"9a� �DĒ�-%w�g ���Q4�vz�� o�>�C[�d��s�avO���K�V-��=0k�����Q��~l�"G2�>���F��\:���b�ke�Xh��..��} A����
�>|�m�烳g5�5X���W�?��4�7���l����u*�j8]S�����n3����	�+M�����5i���꘷�M	�C��ny��1< �q�"��r:��.��¥G;@%�������e"�P�( "�m�r����CK>�Aī~��+��'�κ	��:�i:Aݧ�?=u�r�W֑��qy���ħ���!(Ӏ؅�~�S�n�G�ҖD�3�٣�o�!��$T���j$;~(�)Ѭ�#>t0o8�ܬSs��{{�gyR�����tK�~���>SsnHf9�䕄�6r` ��y�,�И��u���<�դP�PMH~xQm����}P{l:�|�+��(�� �����2�N��� ��|7z�[�����Z�2��O�Κ&����s��F��dR��|�o1��.��'��sd���c�nv����@-�5�C�=��e��'�?	�ID"��`,���p��_���RwuoQ��h=� NUTJft��Y؝S�/R�.�t�3��l��M>J��]��k���k5�y��Ӧ�7��*�
�����b)P3�(�� ���,�vcn�,7_7l�'	+��6B-V�����"-�w��~a$�b�?�P� vN�qss-�ʒ"�M�=��9���~3E�8r͖��gh���"�x�E?5E�����ɨ�����r����y�~��s��~�'�g��ȟ�a�-��c�l|���kD�k����s��(H�'D��B Q*�����z��v!G�����]��I����C�a���"�	���ɐ��*�f�0�DA����:� U��qB��u|7�Ț��Hז3@��g��4kq̇@��j �	��XV���5��Gyr/؏\׹�Y"�!����j��>p�ʃ�#�W��kO�~�\6˶-����	���mn��� ��=Ϊ��s��?Г_o��aP/����^F�}�/�)`��p��Y��ԙ�	�A5����l�]^ç�՛Qv����tF�x�!o�<�������p�0�cT^1�כGg���э�����J�ƺ$���L�����;lt��!b��քC9�����*����a����� �����%J�l�����w�,��1BK ����g��^��5k����+���YŴ�<���c��`ބ���'v��Pl=��o��O���J�����T�q>2՚֣�����4X�Sh�z��wm�>lv��ۓS�IM㛷�S�]�
�V�ԐZ')�Aq��^�����2�V��i_�m��M�z����y;�'��_U��AX�᯵u5�qi��� ��DV�=If�/����39Am��nN߫g�#��j'�i� ��䁸4m�`[u�Zd��٩��넿H�Ct�g����0lp�E��;��w[N6�y�j�4��W%��2�TV�G���tD� �~wo�T�+>����b#�s��m+�C�f-�|^C������~;ج0=&G3�
�^����o.��B�Z%՟p�y�V���~����l�P�~*���E��r�x ��߶<�P�'�Щ����cG�P��z���V6���+L��� �ŝ����&o�	L��7i�>y�{�ӜuUZ�=���-����~��֝��B��)
��\��b�2��F���-��1_\�FX�+���Bd�C��16)=ȑq��Y�"�X��.&އx��{h^�w�X���չ$�Ͽ?�B��ӵj�K�w.'���,yN$�l���<Z���O`�ow�N����
Q6w'���t7��܀ʶ�=�fb9���h�f�;ߣ1�w��5 j����׶���)�޽�	�0X�9^r&�B�-��g��e�|{��5"��j@��G�Pln����g�K�Rh���O�ō\��	���	���O�Xfǜ��V�!�n�'��g׼�F��Z�?rOU�ȟz�^��	�}#AGI ��X���_����Q�è�2Xf���SB�r����@֌Po�կ����+�p�%�v����:� �'X�zПf{��Y|!h�N y`���:2�hgvsa���0)蓕�NT��^�PT�"����4�~]�m�.��3X�S����<�W���+ۺ�dv�$O���$��=U���tGdaE6PlrZ]�WF�0�)�~C�uW��u��`%�u}����{���c�H�DM��P���/�hu�y��aO�o�'�Å@9�zX+�Y|[T0�㿌���w�ý�����>���@���?7:a��4 鑵v)�������_Ց%�R�}a��Z��-�yH��i����'����2p�∢�i�'�뚟F$�:���� bFWuT -����wg۔���������O,��*�I�҄���.���^��%�L-WZ�"ܻ�M �ݴ�X�|v�~�&�*�(��[L�ќ1�1����&�^Fl�o7Ej��*�㕢���wfD�J*6&�'����.m_Z~�1�K��ύȲ����[�n	���~����CCT ��)r����D-��W�v<<����rV_&W2�[m'4��Tx�h<e��C�.�]��}Y�{Ԥ"�&���r���Ld0�z���?�����oF��e��.+��=�F�P��1gC�u�q��@�D<D�ҐU[������]�V���ʴ��H  s7�SA �4ǵ�Y��;IeK����q�Ra�X�)�vn�� Zq&F�ils�,a���
�#�v��=���D/��C�^8;�k�XI�ڀ�$�*���_؟ȃ.U��	��.��?I���<H�+�ȳ�j���E4�C��X7;3�_2�ʆA/_�n��{W��	���:���w�F�&.`���iEk��7���X�H��Ц^[Ҭ���[b��pb������uyA>;?`�0/��i�`��O�IȯBq-͢S*8�b���o�a�a�%�7A>=�^�$��(��Q�ᓂ-�h�u�r��,��1� $�76D�#Q�Ea��8F#+�)Tõ`���e�ݿ��k�����M�Bؙ�¡*����C7
|BC�����Mg'�gS�0��=.�R��h�>�lf��ʚ������#����=@|���u���3��>,~s�E\���������t��;���9��d:� �QX�T�EGk7�h���;.%���-��(�"���i����%7�<�F���/y]3���DGg[�!u9|P[k�ӿ^��0i���wQי���#�X��������l���#��0���͂��KZ����D���b����2Z�f�Q��rM�׺�-e�� q��l��:��^�OY���\�4|(�����`�@��'�I}��w3�/�I���̑�����'��COz�-�qǢ{J��W�ro�����OS�8@�T�����i�l�z�T�0V�!���A�ظ�����M`�RW*��G����&3��)*�.\�yWyvflf-�g��������(��֛7R$/\M.A/��m��5C��]�m��v0�u� NGj~	��\�`D�7�bC� ��E��e��u�,��P����'j\X�%n��!n�A��E'�x��M|�[���)�3�����j��>�6�b��X�,c)�-n��=�H*���U��_N�N�^ bv�
�,7��y �v#�u3Fo��Y�]2��bW�r4�겖�E��_%�Z#�{�u�m{{�L�zyn�x��﷘�Yn��#;�q�`�b-�,��*$�{�����[�Zi�K�)ؿi�E��<������C-:�;���ڈ+0�H�sY&5y n..�"N�*ܩ�6L͌8�^���E~[l��ydUF[|�{�k�2�d.��ᷠ�F��0Β�F�-�f�¶T��I1���G!t�د��M�H;�_�&�YGS��ۯϰ{E,�\��u�ձ�av�9d��\+�Si�&��c��VZ��BV����3���m��ؙ�7L�"pU���8�t�V�:�K;�g�����㈬GǺ�g֯�+rX��-�+2�_���H����A��쥎�JG��H��ä��P%ۣ����M�!��{)�рTV��KCu�GO"�,�����9F�E��C��[�f�cg^�Ҭ����T'�f�q�t"�1Ķ?Jkc4.q92LX�:���E��R-���ɹ��"�WqTP�v����E$�(k���7rąK~ŗ(��l��f��{-dW�*��ϠU*.������7�����Nd��/f=�6\RL>�j�P
�~7����FnR�۸���c�E�Otb?�?�Aj� ������I1"H�EF�^8��y3�Uk�`*�����bX',-�wԧ�"5�RG��:��^��smڏ	 �w!<���=XR�%)/��'�kr�p��u��a����gL$��
vJ��	V��=�λ��>��&����6'���m����@���O�HC�N�+��wInqb�e}��<1��%O��g����G��)� ��AK1�2��Թ{!�Jڵ�gӽVǤ&am�ce��G�w��.W�ӊ�fn�^Y�5,�~{���ڿ7��+�[.�7kbIQx��1p�J��{l��@\B��� ��/w�����2 ��H�J���N#ؖ�|�ұ)\�dCC�i��J�5R����̅>H:�? �OJC���ٿ��q�����"k8R�X��$���l�4�eXsvp������ۙ�q�c�霋^.��ʽ֓R�L_���j_��"���`3f��J<j�Y0g����Y9��Hč�������r�Ȁ��Pn�]��������������æ���g��V\��PG!�!��mɈl\��jr{�&=;ÓBO�_���v�+��ȖC��)Ʒ���͚~��'؋��|��yN��6þ6PV�����f���[<o��D8Ld���<mހ��2�j����M���)��=�~6h�DY
\�����[7aWi�Y*��qZV]���xD��EٖŪq�M�r���!�z\�,c|E$Ρ�C����ɨ5o틈>&]@�c�U�G'�WR�B.��#t�	�.\��I�S"P5-M���`v�lᤱ��X��/�2�\UW�o!hl�B��>��Xt�~�$��ԫUӜ(�?F��U:�� Ɍ#�B[.l��~$6��d�rA�iYY��ƀ�����qf�=]�f�S�` !ƮQ�� >������]�ASG�qJ5^E_�x%����Ci��Q7�!�a[N���@�T ތ���>u�,�4��ְ��}�\�o��3c5[�WC��8/nI���w�
"e/�^'4n�嵃���۱%7qe�K�
�X{.o2����v,��v�=����w9�_��cWY"0�$R9X�7Zir}�6�H@:�~�8Y��������f�h}F+ϯ��'۠��;u�{Y���6y��C@O-�ˆ"}���w�/s
� \��:%$����=.�ܴޛ��S'��u�޿���-ڕ���0Z{�2���j�A8׭��C��8>ႏH��Z9��7I`�	t����G���c:�]�����$C6��
��P�)���U�5h���eMn@�� ƕG��m�Sd)3&�88� ��?=���xj�_��		L�*�F]�v��Ƭ�f�V'�����^~�4FM�7�B���w�	2)ܯ���Ee���Pz~��n���:��M���G����v��{qa���j�AI��$l�.��V��� ���-�N���x��Ԉc,��D��5cfaq��wȌɺ
��.�#*�3⽀N���f
Z�� �������,��Y��U�d�Y��P�v��Z�h��u���L�I5d��`BV �Ei?H�qHF=�B@�fn���rVJx|֒�S;�����_fw��D�����h(���,��S�Sh�k�no���gK���� H�&�m|����k��)O�'d�$~2��V�r
�OJ��R}Hư�om>���ZxN��1���ɘ�_?����ID��a.Q�B����%� ��;$���.
�HqF#`�$u 94�~��DΏ�ل`�A���	g}���y���G���`-����<?��?�"MD@o�n��{����T'l2#�B_-��#��uq>J�N�\Guj�T7u*��e��0
0"��=[Tj-j�f��r��|o;��(oݠ}H�����VXNfiM��&�N&�D�Ow�@���s�8ǰ�H{}/CXl���{5R�&,�\�o$�R�l�Y�?����u�t� 3�����s�JK����`S���H�&ָ����[��u7;�̽���a*��蔡���V��EZ *�(��>_��!�����:}c�.��@$Ul�Z���R��6!k����v|���?ba肺O�	�)-U�d�L+�\�[e*�Ѧ��u�߹� �~�F������ȉ��6�=�?c7;��t��D��3����C�1S}�+EҐj�	��o�&��~�������6�]"�![~��gg��'\dN��'7Π��?KW�:��f1�)߀��O���h���1a�a�Q[\iW(�
S���tgL�[�+��5��y�!���|yw���xlG6�Q��:�hX��6Z>F�Q>��F�W߹o9����ɾ��uT�u0`����?������v��B>�ë	qެ�[������lt�s�_�,�|�z�@R���ǖ�X�R5C}��V������H��S�CIHNԸ�%��n2%���P���5�����'��MZ�fuC�QR�̺M0?^H��O-�)�h�Ja i�x�6�6���N�I��oH~�������^������̊��**X���.\�لF�|�M�<5����%�P
i�	N������r���[�K�v[c�k��"o�)�f�hC�p9,���U}9��>מ�Y/�� ���m|X��i3���Cu!t�}ݚ�D@msF��!K�=X��TW�׀�.��%�H�P��YL�d�mFI7��%�0�]�)���^Rы�5N�pt����z7EX�
�����z9�]��lU�(�Qd �h�#�#d80�[�f�>�O��u{��t��.d��x���a����~�]4����r��c�gI6���LW ?�H���g�D#����+���+��K7F�,d?��VK�%�.^��-��W�0�&��&/��O�?�E����|0��^��4p<���&���	K������/�㱂��V�z`|���la:�YW�LY뼔*B���j�M�n�o��0�.āߦ�L�Ţ����g��º�?�l�����b��?�QPsb+�^3�}3�4��cK;�T��XW��.���o�,��j�L��X�%;G޻���cWMǥ ��kr�/0p�����A �DL�P���ze#�P�/1q2�Ǵ6�}~��ɧ^23vm�g#��H���uf���$�V��|lF~L��O6�#��EV����X�=���o�J�>���h��Mix����"ӆu0g�)3�E�)����������|z��!� �a�[����ݟ�Yo�
]�\�`�e$|�|�	vcE�߲+���XGM3\Reaa�[)"��>	��g, .��ޓ��,:������^RGk�}|����qfC
	L�(.Ot*!S<{��62��6SE�g3,�S*S�����'�`�-�}��F	�
�.Z2eN|F�NE�(��c=�{ܑFu��v�I�h�	�d�ӎH���rY�q
#�W�	��xԔ�E}ݸ�9V� ���û�!���>��{�.
�ܓ���hF��/��f�ZW|7eA-A4R�Ձ��+��as��y��0�.U�T�%T�,�|���$f���1�c)��l�:��{óH�~<�J\�~�������F�_Me��e�N3y{��`�r�'���{u��Vǋ���5��ђ?hEXq��L�;��A]S)�=����o¼�^=���z�G0V��b�;ok�o�{��e=�oە��n@OΤǈ�+�X�|�;��_��r�����U\O$f30�V����
tO2��hQ��g��3w	|Cm+1�������f��L��q-��5����ɼ����_�"�� ]�Ŗ��Z4�IQ�ـ�Gx��5��1V����0�p�} ��BTyy5;��xI�a���4��IX�;��~4a6�	�l`4�֥+ա�'�G�a����tJIy�),��19�pX��ŷ~��U��8�#6�/�{�8]E�&@��X�����ە~3���g��� ��i׹V����V��eo�I�h�;�3�� �[�@�}�or��jX�g�8�zq��e<6}[l�ȒK˸��T���G|��8OE��)�v�Vu1�j�7,w�������BwIX�1���u���~.�3�U��Qy��[`�k� N��X�,�e�ZB��;��
�&@rTE���A�~�@�t���ƚt8okjO�K�Mj�x��r��U����ڠy@��vⳞ{����R(�"9�|�H��t�2�GH|Z^���^�\���Y�	Z���r��������ܹ��(c��y=8�B�oK||S�t/����A�S�S�t��1��eHz*�ϘI5�2{*|2�o��������).q].`�q�c���h3O��X��kX�;�1boڶ�}H���c���/�q�4�:����+����T�%�If$����O���xIy�7�a�heCy����IW��Z�8��3جD���)�D�c+��<-��^���b���q�b�8u�y8��pĞ�����f��N���&���'�>�M�H��̩l������"��Y1XF���A=y��kC��_-wۗ�vǢ��x#WZ��Y�tt=C��ϴ�z�A1�g������jP�!	u�ٿ��.q�����jD�^J�6v�D���T�Ԓ��Q}-�L3�jN��r�����j3�D�t$�j��6�*��y$�"co*��J./?�z���9	s�Q�#����`�,:x�}l�I^�oL�}^�4�i��, ���A��'�5P��;lp>�ӱ�Qs��L�����׃)J��H�%�r��Ӂ߭K�-�&H�ӿ�����}'�?ցC8����BnQ�a$��/ ��|�WiSs��֮Fv�N�,1) cCN��	s!���)�vwcH
�����RY�=�D��;&�~��N�~r�6/&B�lHW�!#1��9�޵u��P��B�����i����+�.C��,��!�`�ם�߄/Ʌ{V�F��HhM+�;5{}I�P�Y����uS��U)�򟄕e�|�c���Wʹ'ir�Ua��b<�J�6A�<�4g�౓�2H4n���K�g����4JT��*��\�O�9�b�sM(4��l����:��8OU�����㑅6��A�/f�S֋)\1�����-�9�C���04�N�2�?Lg=k� [�7hQ����й�g� V���/�q�,JV3����?��m�P�
���M��$�BW�џj>��\��G����؍�Ѥ,AA`Q���8?TD(
ְ�uvB�}|�o�y�@����c4{�T
:��I���7��a
��=6���!䫛��
kVICI_��+��?�\�
����K��V�k�:_��_LU\c&d�e��A��j�H�r�Z=��mxL�kDG�Y6G\���3�AQ����5�G��~��9������%���U'���hBˌ� �9�����;3`�W���*ԙi��c0d~�P�~�3q�����uj3Dv�b(�"� �1��jG���v�_1��^�I�m^f����Z��ۅ�X�o�$H/�#1�������+����x.�UX@�jF����Ŀ�*>�r�.��I������/y߉Iȩ~-�O"�lW�sA�r��P���v���iwWկrY��W����
�X��y����>��`�􃥇�`A��^+��l�w����n������u���H�_'��@��?\
%F�Kh(6Y4�i�=�E���.���c��i���o:��n�}�:�M)#�$��0�B*���D���7�[n����L�.�gih�,oD�¦����oAS�y�C�p0fs�$S�����������~�J��U�� ww՚�%P���"sbA����!��[�!�A���i�`Nog[�X�"ػ}�&��˙
]�ѐU����Ln���祣1�i-�����g�����/ S�
��/g�F��,��,,u���R�v$�@f�Z��lb�_�w�/���d��{�6v�]C�Q����ٛ�;�?�~u*���Fw�W��U_��Ϭ�R��3�	�7�{yp���巁�]{X���d�P��*=����z�;�%n�M���)���hu����)���l���4���Y&�z�P���X?"�L~�K���?��ܸc"j�y�"�H�%�>�LT���U���A���9뗂t��:M�w��K(_a�(f�A���uv��!Ϭ��Y�]0ú0)���S(^��Oa���X�Ƶ��H�u*����7}-3���g|�4�}�:ۢ�mtwP�>q����&@"�nu<��}����<4s�#q:z�!΅q���k�����3~l������6��u��B�(q�`�<�NS�,*�Ok[eXj�����m-1��	�_J�������ԗ�Ӽ�󁺊�ҫ�� &���󗍐�q-�^�M�+��r�_O	F�$+K�މn���2 8����'����w��co*WR��t]O�~s�J�9�M�I4�����7w�֔N W�P)�S6c$���h�i���x��q���੫E.�P{1��ԤjzHu��(S �Ox�<$�$����u#��q�y�[�HҌ�Uip�f����ʍ�rW3���)�V��D�F�	���@[F���Hl�����4zgS��p;e�������FƬC6����'�uZtwv��r�ί�V�}6�d������M���g�&��ER�{ME_�9Փ���3�~�R#8/w?ݘLW�O���T�=�t���H�1������S�,��NR���V��vd�8$����j�`�I���u����]����$(iX�,��Z�i'_O�iц7༃�v�0��An�.�ML�|��5/H���Q��ܽ~+~BD��7�iD�l�̀�������t��k
:pIyD-Pu��{�����'���1��@������ȡ�E6� �sǉa�tP��$�Ï�	xa�f���Q<�<K h�ٔˆ�BqH],L�-9;��r�l�({��Lل����\��C�+�̸١�^��r�V��em|�3B;�e4��N��uS��6�I�l��{O���o	�h�G���FX�h�
���G��j�5�<ۓ�~DzB����x�P%Y×$�X�e�ح��:��S\��H�Ћ�d�i�T�S��-`u��)� ��ơPm�V_2�j"\��jV�� Xص�>y=�%Z:��k��=�#�~l�v�qh�.�Ʉ�ٟc5�	D�6�cYS��@9�k}��W�nKC%0,����XJ~����@�z��!��y��峴mOV9* ?ҕ�8�5�l��(�TbU�غޥhBĻ�o��������V$�]�el�w���{+f��:�7��_^5Kkd����7_ę�Mif���7:U)~o���G��$(�5�Z��ȹ�X
����V;}��Z]}�����B�Y5��O��Sh�V�⼯S��ѯV����� 0�0i��v78`��q���鞓0+Ɏo9$�&�x+���O�>8X�;�B3�յ��l�Hd����iyW>0<��yK<'z��0�|�&��@E�Y��հE����*��Gۅll�JM���%$AjmNUq��^��wf|�ъ��j}�[�c�<��.��)9o�Sh�vЯ|�{��8ź4��ě�,�W�(�ʸ��!��R���]9<mTd�7b��vT�c	G��l.W���/���mqk�|���x-��1@� *� EU8Q��O����h���_�V�m�`��Ǹ8G�2dS��jʅ�(�*x�����L%9?���^`�̻�+@
�Q�jlط�i���v�q3-�E�}I���k��̪��'�6
b����5Yz<�u�b��>� �����b�u�� �H]�Έ�y8Y{��Z�JR7x����+N�)E��Uw|��p��w<��g�b�T�Ð��<8�_�ٰ�xPݢ�5���B��7EU����O����������d�^��m�u�� ���hh�p��W|�,�`lN�o[�V�0��%��t<�9�拈tԤ�Z�夞��
�z��#���^�V��	ғ9�+�>��$kyKOvEd�_����d�n�Z��B����N-��溜�"Z���?rY;m��O�#l>�W�)���_G�-��� ����XF0̡�7f�����9�U��@5�}�e�Fx�\�@���=�����(y���ow$�����'�0Q<�ay37 ���z�ˣW&�R#f�ͨT�
uS�	*�!��8Q}���̍]�e�;;��ީ�H�E�;�.����Xo��`������	����Z\[��].�zN�`���b�93��2�:>����0*`/)��<�<���\PK��b�v y���0z48�Dx�3�@"J8p>��<e)fG��yk�\奻#7�ё�pW���+5�6۸�x��z��n�`��v��*b�3��nW6�ཾ�9���㪳J��c$'���@���TlJ/Rϓvr����e�՗@�2�W
79���)6���`;���%Z�=�C�]���Lڲ��:*��:��SQ��
>��YH���Z"��^�L�ݶŋ8�ɛ���ڛ�O�ڥ}[���@�E����F]�6���Q�|�����K�<�4W��(�$fD@��:��K�d��������T�={�X�e��f�ވD�-(L��nVQP��s%��q��"�G�2��s����r�E�~���2Ym���w�w="�	3Ŭ'���5�bq9`"�	� ���b5�lA�ʀ�0��y6�ˉ,�£�p�Up�AM]�U��!�J`_�]�jP����Q�ڏ�_Y�-y��rtrҺcq�+ǚ����y��[��K=�+-r���N>�?+������$-F~��?�����=Z(�G4E3�W�$3��b}�S%�{(#�[>�4e6�!T�խƽ1�F�` ^{����[��ҎՄ���e�h��vQ`M#���aG)��	R/��U�1��]��.���Q����mwk�	��Gɟ	��L&�F�N;��8[ҟp�O�e��C5�%�7���vs�/V�〿���
8��>��������5����Ӑ��N����ZZ�ŏ9d[cb��ɼC༶��s2��j�䐹fH�0��f`��F�X�^\۽N��f���F��T���@@S��>[_����i}+��ֺ"�cQ+�Z
�- �8Y}0+���X� �R_�]�qY�1^M�2��:�����plʤ�v}�G����Ԇ�&�=�`�$�N�~��s��O�Cd�_�Ā�\S,a�u���6�OBW�X1������*�QX+j4���3�%��#����¼&z�Ҧgh0*��B��2�r��A�nd�#ڞT ��e��t��������P;���d  ���2����^D�d������8����S���������9�4�����#���\�x���wK�t���`��!P/#�6��&?G~��E��&������R&\��#B�D����gG�}�� :c������:���9�8q���RC����X
Õ6h��і��vs����:��.d0�Lm����MP4ӝN�_�`��B� �g[7x�8Y��*�e���ޯ2w쌄'��nH�Ƚ��$2+�ZX��~��b��S?(Uo����ݦ[��ء��K���zX�~q;�(�
� j�V�|t��%=d:o� C��!�1��;�!E��ݪ����D�<���,�"紲'����k/��B/(�Z���ɫ�p�'���MV�Anio4KÚ5C����c�5Ћr~B��p��{������u{�ƿ��M���eI������Hæ��s�뻘�O��A��{����Ŷ�x�E�<�f��R�H�`V�O��`u�5ƺ&��|�y��.���8c�sU��U��0,y�-��%:��+泴����o�K��g)|��[�jR/V��dr��N/�������O��@y�~G������Y ��ڪ��C��-�N@�	
c�NJ�E��]����^O�����1\�Y�?C���T
%��+�~�Q�]�9b\��������}�H\�<t�a(��N8=�+%�wzC��k���� ��ɲ�ff����^T��Q�f��|�DE���Ay�"l!�Q7�rHَr5����\�4$,.������0�碷+Z�kH��|lɲ��ܭ��Df�u���CDp�%	�W�#�	�9���љ�� ���!�e
EKT�$�l&���?T�h��s
~ �˪�@��]�mjVN[��')|�v�����j�����oS18�5|i-u鬶�kq���f�l^M)��g��E�!U>D�1���"�~�"B��R��v��ȫ�]d7����#�b�->K>�����W�(�N��_����k�v7?Q[鷚f����\k�06G%/�\�"TEC5F�ʮ��M�1"�e|���,xK����������?h���Lv���
�e�pO��Nπ׉�H�����v㈜Y�. �/(C^�Ȍ}gvUm���]�V	;g�)��	E�:��������_S*��? �49PHp�M����x*�D�\K(�l˨����B�:� T-��e �&O�n�G;�Q]>k�5�z�*�##i��~"bm�޵�����H�}���Q���G:�������o%7���j��í��&x�mk�q�v�H�nʌ�Z(A�Yqn�_��� �g�l��;;�	c�-�0���sGĸA�ܺ~�l0B�R5��`���sK�d/ɰ�Jw���co����mU��D��G���T�KI/^qSr@2R�6v�Z%v�[5����j;8���eh4ʛ�G�C��a�`� 1��T&� Q��Z�������5!�]Mu��1��w3\�Q��"B;[~\d��`�O�pH�9�x� ������ZD/ҥWR(���N#�:�"2%{P��GLFI����+����+,�jO�4�IS��3��zO�B�p��r�"!^���g�h¦c�.dY�iG<n�[�QQ�v�j,\jjH.�u8��U���y+���6�Ŏ�!��o*��c��ͻ�c���x0!��{s��z`��B��O����$�J}O��Bd�u=o��Ǔ��^+�t�PK��n���eg�5����ޮ{Զ�{R�ӄ����Bc)��`ԟ�WM(�{kZ��.�_�	�Llz �_[���pWŝ�� H[.�LaW�3t�s����,����]q/��q�~�/��'�o�gǩ�}�ǳ�7H�����}�܌�|�ԃ��աg�%����`�4���QA��] W�nҽ�YGn�%��%��c���H�4ɭ@�TDR�_���4P�0l�VF��5�A�|�	5�.��.c/#k�i<��s���	�g;��U�%��n�G)����θ���ƹ��7�W��?��=GE࿽�f�`1�\Eo��S԰���
����.�Yw^Y�D��k�R_m�B���SO��?��-ڐǟ��7e�d���U��(�`6Szm�qG}��� B�-A��(�٬O�t)��PW��-� Sݷ ]���5�T�띆�y@L��زR����
~���v򢢯���/�]f7і�hf@�@cn-݅W����y��%&��eq'	R��oO�/��<��~�-
��=���S#��)��8q�;-U��Jux�e/����P�¨��>��k�TJ{���1���/8�ig�i���fȃ�y-�(�E�NԙU!�Dv��TS��� �μ�6Xm���X��-%�¸��t=ɥ@z �&�d9��i{p�=�kt��[�y����'�y�9��y!C�؍�Y!�Q9��2&��.7�)4t�b#s"�$�W�.���z���$�͗�p��`��l(�P,��I�q ��Cuu�D]�,��_�n+��Ti�	��+͹EqȘ��!���D���W,n���14�"m��v?F����Jd�\�ܪZ���Xb�lݮ���c�5���L���׾�0�&o�v�,���1�9q5���2���S>[��.�&������o�t�.�b?��S�1rh=��_��9�������U=���x�8���@ �["�,C�����ֿt���OIeqi��?�~����]��P�b�0;>z��j�D�_�jl}6�``n�AT{�K
);'�.�mÄ��,�k $H-��\u})�-��MVJ�ERe�5��ȍٯ0��wL�2���-��V�ʳPߔ�%� I⁢�E?�2=�hಎ���gn���S��O��,__��O�m��"�A;Ӵ$=�i�e�z��m�4��A�}>��$���0�F���m5���I9��%�B
�-++ZO���ϊ��Wy��Hl����K��^��%�S~G�iL��@�]�6���K�,���T�����˃��zĹ��㻼�	����#�.]�G����zu���ϣ���U����O,��/oG�-��eOAV��\��n�Y�vQ+`Ii��=5�&��½"���g���E� �ێ���A�� �ctEnx��ʳ";%<P�g�H(g�UlAah�)?8�Hȼ�L��mO	͵�U���|������D���O+<�t�.��iPbp�5�巖w_'S�@�y����8����kR���jx���W�gɹxظE�*!?��bӦ��LY*��!
j�
�]��([�z%ܾ�u+�G���=�A�=��!��Rm�Wr�u]�G�����Z	��e`�͋��N�˕}j��űN�?��hX�s�:�g�������b�ve_:��@�!T����ޯ�������ՇY���7����(��<y��4e�u�
F�ǠvS��y�Q���YX*SnqO+�uyU�}sl4GC/��!���-	��ӧ�Y�C��i�Gh�z�0�UB-G������XJ��~=���f��É�P����v�o� �QeK���8y)z���DO c.H"��壟R���@�-�aͦ#n����5D���]a?)���H�����jM.�h��G#�+�h�r.��3�W(�~���UyV��;7�ȉ	��&�j���W)�c�Ɗ��p�x1v�@*ֽ����������u9v�E0���B�|��k�f3�9j����pq���J��x�M�.{��V�.N���z��O��;���\��P8���كyx���G��N|֟�l�ȩh���r�tF��O�_���,�s�\]ȃ2W�0֔����Y!@(�R��L�W��9���%����	�̶�H�E�Y�9�_Ň�~���3�P��G2#�0F�I��1�Ё���jʷ+1�Q�2�4�߈#�V3�{E#��>]f�B�)�KT)�3�R��ŵT��:�1���A�S�|�#��Ta����?��p�}�D#�n�
K ��Q�S<��b�U]� {�}N�l���s���s��@��	z�|q�j�m]&������xd�D`���i�bw���E�� �}c����@O��L�'A�D1��?/��-䳁?ɯiy?s5�����αB�^�o�2#�ș���2|�O_�y/!�*�Śe�A�R�_�Qa�{oC��&D�����V�gM��qR�G;V�@�P����t�����]�2��H��-`�_M���Wc�%�+I��-���:��x�	�CI	�@o������݄?|��RD�ל�ǵI�Jx^�,�߸��d�{`��)}1�>�Ǜ�Qr���}A���a�0lc�U���"�/���C�k�%�����qr&?�Z�����N֞"�������Giu�M���pы���~�`�'���5I��q!z��]J˸DN�r���MB�ظ���ª.�Һ�(��~�����YP�dl�F\���s�Q�y��^�m@
����r侤�δ�M�ɧD>� ��\#�V2��`pG[;MS,�{���y=Ylv�m5#x8�+Z�q֚\
m��$��X���#����Y^�K��s��S�,����x�硯?#�c��_J��s �3p0H�Ð��^��d[��<��t~67&����Ͱi�޴e���E�+�h�������A�
L��}�	���Y��˳��G����;��^�����j����ߩ�Z|t`�)�=�`q�:H�v�օ;i������z�P ���G��0���JW@�%%�pD����?��`P�:��!����B�g=�e-���'�2}�V���)
�7�q��.��Ӷ\S/d�%�}zat�Hz3�F}6�Z:`?D#��b
A1�'5�烉�/�����	(O�$�p-ƃ؟����(FW�w�m.f��Zݔ��%b���2q�AN0a�!�q��k �gZ��"�
��<�8���Q6Ij������Uphs�g��������mdϯWT�xSܬ񯨴Q��ښȆV��c�a$>X>Y�h�CR�G �MAa�N�����<D�±���g5q����&��k�mI>����9��5{�{��UR����ڤ�V����N��u�	�㤌�A/��C��P�Y�t�J��yACA�H|��F�����V����w��>��w� ��)�E��Oh���L �*p�񨣭+S���"���~)���brd)U�a4�g5�
��/bO}���������u �Cî�A��/� ���o���[{�G*�pyNg�����n�z�q�Sf� :����`��O?�z��\���l��������	����C�x��A�F���0�Y W�{x�����A����H깏�^a�[���'
���f�D$�I�-�1����3(��X�K:O�k%93r�L*���#i-��%Zy�7�Y�Ӈ��hư�6ķ��^��"����TQ�FV�Y���������ڲ�^~�؞���f���I��z�ȊW���z8�~z������#*�S�!�r� ��=�����!̟���a�g����ǌ�� ��0^��/+��AK󛇬V82+�CSy��6	�[���6�`�J&�U7�	�g��I�%�����L?�Q0��U�M����+@�Q���YG�F���F7�W7�I�&M�9���Wp���ӑ��.�
��:V�<�x.��o�<32��wM��ou/n���]9�����'���&�Ḅ��îj��C�f1uCR�:�wRHM����}�n�#���yn,Ʉ'�t�u�L@Ƃl�D�.{�X����ʳ)�'��ӎ�!���䁦�]U*����+��O�p��x�9~h]t_ 7�[��ZI�_���a����*G8d,��'Y�%Z�����}�C��Rb/Tv��L=e�:K��ΐ�b�����Jӑ�.9������P�����W20���l�/0�,a��`���L��N�W�Q������f�c�����f��݂2� �;m���Q�yDL�V����j��n;4��A00N&!�XN6��,�����h�j�,NA�3u�W�� j�nT�2���;��-|jng�H>W��65�7rW�����jF�P�|��z%D�^����@�s�F�
9|�� �@�f�d��g~a���J�7��̛
[M��6Ad��\j���`�#6Y�sN}�f>�>��s�v�b��5
������~'~���\�X�}�eCg��W�QK�uʙ��~�^-�T���IL*�n���x�,O�S��	���?��A�3�����o��L0O��%����'ˇ7�����7�l�g�ՉJ�H�B2�;�÷��i7��|.���SIR�%_đ��~�~o�+��My�H�χT�}�%�(g��}3��5�04��e��`��ߓ�V�J�a��ҿ���kѻ�I�x?G=�'���jj�@��c�l�������]�d���2k�2&*�%�m�ݰD�tI�rD��^���M����4Ƅ���[���Et8h,�:<$�K=6�c��)��F�%�$�3k�3;x��u��jC����ܻ���`K:{:����.J�����푊��D�߅�i�7AR���c���$���\�Ml\I#m�8%�b��}�����x���. �o��=�.J"с��ݛ>�*��q9�U����>X�K�U����@�����V��_!
[����)i��M����Wl}�xBS��T׶f��[�*feX�u��3��B1�RA�"���F�5�W�(3�j)�N,h�L�-�:xpp�Q#�5�Bo�1��3&n��{\k�|o�B�'ه�Ӹ���|b���9�cj*���`
*���'S��w�Q�&S�5'iK���*���X<��`3J1U��U䥰��O��s.��T�Q�4"XOu�t�n��("�1�:5}�^��Y�-��U1���ĝJ�?�������e�7u�.}�-�i_�26DX�#2�^�C%#8lQmXq��IOP�ڽ?�!z�1
O�T?	�E���v|�Mv�V�%�L��sI�~����Lhr'V����Z��ı�"�^��#9���۳f�vt�b�;K� ,��6շ,[.�A;		p� �ԉT��6a&�s�V]�1I����HG��N����.�K��w:ؘ(�\p�Ny�l����?����I�M�]̓.^=n�De�\!B�c���{�Ut�*���z1�4v���ػDW]����"����թ��-��*���Zk�~�0�)�>7�#�˜�9Yi\x3c�0Ze.)���?���T
�0�9��wsr ^oEW+���BF	䃪A�*1��)���``h�d\C.A3���!q':��"�	��ד5�&���{\�7�kX������PTv�,�Ǐ��R?��	�kGD���by�34���`�|������>2��h&�S�F��e���Wڋ��Ά�l.뺅C�@n���W��z���p����qؔ��OB�6Z� �nT�l��p_^M��
�bVOrԦ�L1%'���}{*�������^5�`�(�/哺Z7�W~���x�\��@�������g\/l���i�Y";�Zv=�e����HZA����0�Z���5N�����N�)�$��G�<��>�"�V���	�bQ�zK�z3-�{v2�.6~��˰�u�_@`�c g��Y�V�&��n�1�O��g��)l�t!�: @'��C��Zq���r�t&�҃�Z�eEm[Y�KK�!қ�jB|i����&�����
CR�\j�B{�Z UF�G�u�.Ւ�Ū��G��<�O]�+�;�ȵ��s8Vp<.���m�4m?iz�~��9k ȑE�ß�>ap.-owZ��0қ�:������Q��	I��<F�4�չ��+�k�U^�oC�r�P�'�w�n����/ ��T�_g��9��:�]>6�7�(U�O���ױ�����82���41�W��{5�±#�8^��#R�r����,�% ���V�6��?�%�
���@�^@@����AaiED+�hׅ��[o�b)� }���&���˷����!�e���}+M�.�ŏ�}�p|��oT]�'��_PF��̜:>كWi���n���>r./m��ap����QR�F�BZ��/�:���7y6�Tw�F�E���k
b''ȄGI⟧���K�i�+ti	�VF����B/�N��:�����e��ܙq���J������:>�4 ���(�X�דl�ô[}���c���p�@t���G#�)ʥ��cm��!]��GJY�U�*t�a�l`��\� �ݬ���.矴Ny,�� zn�e��`
�Lz�&@b�^Ø��m�B_��z�K�eؐ�HV�?�M������tڊ�T��ˇ���a/�>΁	���u�7���]����4{�IcNfSxm���	��=[}�Q����R/`<�����C����G�9V���cY�Q�kS���Ϛ�Q֒l�� �a���T��z��X���M`�g�;���,VWvJs��M�X�ʃ��[DC(q��-�Kk�9ӋO�T��2��������VE4'�`�*!��uu�ѡ��»��Co m4�do�%�+���2�	)�D�	m���y�N��O4#�k:�B��Ǫ��R'"�J���䁼i6ʬ�$�����@Bl}?O�wboSp�Xw膹�݁���P�r��n}pݩ�Z~<;����.�W�&P�t�[R 7��ʗ05���T�f�7b�t��/RN�%9r鏋��b�v��q�&�G��g�jE�dp�WGs��������c��fѠX��&EE���Y���|%HH;6����
l�	5��;^�� �J����<-6G�U!tv zR�׻5[ԈN5�,�]J��G�R��D�G徶��R��hβ���g	e�IIs1��>0�����F{�b0���� |J� n�9��6�<����}���_�ȳ$y����&+�����j\+ខ �Z�_�`����D`��,m6����r��-�����:����H�*{G
��{k���f��f�,������`&i��l� S��.�d�|4;q!�а�b_��&����UۈSc�G�����_K~���*�Cy�S�Zۻ�f���<�����L����eN���hM?���b'W��W"*�ҋ���g(1����:��P����'P�!E�Q���>��/t匄2F����]1�/<O*9d2+>x�$<6cM�^������Ͳ]�=�$���v#�o�G9	�V-��]�آ�`�L��3׌���� R*�<�VV����ECX�l��D���S�CX?�MCk\�Y��z�u^Oރ�pz�Q'Jnvɬ#����BOX[Ң�.�%s�E�`�YC�zr�*���7T�!b�����j��_��ۺ݈1EJ�Z�@�
� V��q&��;Lu�9&��Μ��	�"������1��}�J�j�]�r"�2]��m�hVǈXL""�I,&��n��Ռ<��(���ʃ2�y�X��U�/�D�:�-�:*Re�e��x���4��UJ�I̃�?)m��{�:Gւ́�
�
��E\f��h]���"��8H�%� =��_��֌V�B��a���L�� ���^>��8��3�@FÓ���'
W���7���6�Z��x��B��)o��]Į|�ޔ0�������^sL�NL����X�� `�g8���XX_�傏 P�pd�!�b�8YS��uG �#����>��t@Z�	7�Y�����jH��G�p�a��ƀӣAe��S�T\�KpP5E���%8r���Kc	��X<Z���@�l����TP��MitOV������`���!\pK��"��8p�W'qR6!��-ť6=�Q��Z��)�bɔjz����(�\n|�C��l0�Ȅ�z�}Mz ����I�Sv��n�g��~�8�/�q�k����V_��.a�I�%�#ի�� ���H���Jg��s�'+r	��ho״� /�$�t�C�.�+8y6*_MbM�񡔻���w�����A�X�nbKq�M�K���#��X�.���G�|&0��	#!g�� }9D-"�C��B)�ᵮ$��­_	bw�N��H+~0� �%����cc/������&�L4]NrJ��gK�$�<�e�QE��T��K���ho�U)A`j�.��V�h}�/һ}�u�;�"����\x^��}u�	�}���[���'nڇr�,\�ߍ���}Zh0V��j�Q�[�'�.��7h���YQ �a��.�# �Ľz�ÅH���MS	>p�.f�%�W^{�e� �(T5a�kD�����j=�躛~��U}�䝋�z�ūބ��䠠�R�C�|���5xit0i�w�d�B/
�#}��"z;t��4Q/�˞n*:|6~w�;wN�����v��L�W��c
ڝ���;QH��Fl�I/G�'!	���ݭ7�j��gO��~غ��FQ���+;����[��>�أ����Kbl��2P���s�D����ׇ�2m�w�M<:i�}�09J��l��#X�ac�����P+�%�[�$mj���;����/��
������I}���+�[���U���t�&�/ ��
��L�`��3����4���T���Fzة���l� �H�'�e�&H����M4�l�M0Ň&���x夔v:%<�8�׋�Z���z����O7���(�15BiKY̬\H�f.8B"�@��'Ƚ�I��������#h�T�XD60��K�I��:*��_�:@������8-�M��h�-.ѹ������֓z]�y&�'n~�з�T/=,�Y��gT%�ލk�A�Dy�)��Z�ih	b?X ����YLNr>�P��m�)�K��pQ3U�2��8p�6����6�����	c픔v*:�r����N�i�Пz�L\��Lq���~��"D�Xge�Y�\1˘k�dz�,�x��%?�F\�?�^�`$�_6ޓ�"��L�c��m�e�G8���;8L�vj�f�\�ek�s��r�Qƴ�T�ɭ�`�+�f�"�;���OXL��Vᚪ�Ɖ����X9Ns�SY$�[�i9ێ�V�T�-���� �P݂[	�t0��b2-�3���D�-|m!*ey�0yI��	��G�+�q'��~-"�����c����)KC+!@��������qy&���SE'��[6H:�U�����kV1{�j7���+��츋$�������])���m���%)�����Ǫ3��8�7ː������ �Ȥn�t���%�A�f@��͔����q,z�w%�_ӟ�?J�=�1�����k�����>Ɲ���I�����rm���MO�1�ܘ�(�f����u,/L� P�
�I�	�$,� ����>eу!�%�>��V^b�f�pE�d�.�L�?�P������fiS��_It����s�1�Ј�̴�ou��qWIAXU�'C��Q(/�&�G�D={��`T��	;��6 ���T��%�':���_)��H΀ݑ��,1�����6*[R4�I��6�Y��l��k�'@�bv����p3�������I,����1�jL�Y<�"���P"�l"C��t����� �ߦ��q����}�Ɋn5��9 �1fj�H_4vv.�\y�o�h�ɻ���@���S�s��t�E3�m�� ����ũv�q�<X��4�Va�cy����?�v9��E�P����[�w^!�y*&3���&�4���]`)���2�X�ތ�c��я�>�q��G	\��p�pq�6C�x+�[sU�G糷�����u�� �}�fYZ����.Ha���@\�DЧf��TӜ	�� د�Z��h�b&��-�T|��+oV�ܼ/��
�!)�)��&$�4��Ƃ��
t�#�M��������X�<�9栐PV�t�b�3i�T�ݍR� �イ��+��#��N �6�ס��J��ӄ�^'�&��u�2�� �B��������P�F��n�f�Le�=��p�F,B/�sG�(*�������;���J�S�"���@%F"b	0�:T&y��;���n�=���ۅ!�t9�R���Ȥ��{!��#����%���/����䉷��\K��B5W9����g�wM�XY���Fȵf�P�}��G�P��u��} �eɼmn�׽V���)���Հ��Đ�i�*��l0���M}FO�(���Δ7ջ�K'�^%�b���h��7�sy*���~�*�����O|</<�ѓ~I�	D/�F��4�<b:�Q09MΒme�F�\��.�c� ��[Z8_���ّ� n��(�	��1�'��rt��C+ds4q�8�����i��IZ87�}4��/liL�ҙ�$$:�P+1Ө����k������������?���sl���[�Z��zؖY,�h��ξ�W��>���H��øGer�!�h(o?[Q�"�ٶ�%��ɞT%G�R��������PS��i|�h�u����)sﯜ��9�L.�*AWc���,�IA෭����Jz�F��"4L��yI$��@����г�H�S�~W��5u��c�;�{�o�����u��
gE�La�ധ`[�Aľ��o6��恠�UP��s��9r�Tٰs�	�t}�K�:6�-lѝ�©��F�cmKH��|~� �O�'��]u�=����r{A�-H��S��%Z� _����,�gb+sTs������`����ڏ� "[��4�9�n�Y`^;���l~����������@'Y�����w�A���w��0<�
�U�e'��3ʕH���^���Xe�q�q%�)u�#W��&Q����w,g��~k�8-(�r(�2����q��6F�b���~��偳ɴAn�gv���ۣ��U���ez�W����S�GYc)�W�V'�B��,�W�����?`|K"z����h�w�vj�p,�yj��	ׯk��8fA�;R�ۇ�|�p�5N p����3V�t��� ����@ J�@�t���.�I�8�F�\<;�-���V{�����G������z�U�x�'T(��uypLU?�F{ډ;�{�tܴ��|A�| ���hl��E�eș��.��x�?4���K�UH@��[�(���K�!�A��`04���]3r� �g���B�z�ih7B�|�	�zgo�&���9�˽��5NF�ςr$\HGj�q�q���-��14ȃ�D<�k��NjqX��ׇ_�Q���mkY��b����D� �<��ƙ]z��<I�M%FZɜ �Ǳ��%����C"��<�����Q�����,�Z���aa�@[qA4$���O\y8��Q2�Iv�+C��KCL���J	�]k���2)}��b�V{/E}��8NB}d�8&A"��K.��$��K��x����D��L(����u�5G�L�HY�B����z�E�D�9ŵ��և�q����\�?��Y緅ļ{	��<rb�}i���s��ؿ&hv_� e�Cin��_�` ;�����(�8B'�)0r�0�3�����]R��V�+,7�n�׊�3�o��o�[;	k��+ ��2Z{�-]!�K:�M���N��K{	�P;�b!�?���~� ���h��Z���kL��x�j�zn��.�Co�bqS^��l�$z����P�0��������s���y%Ӆy���S[S����r�^����{:��[e	nqk�׹�3t.�>�W^����#���K���6;��"�VԳ]�g�/Z6VK�<|�*�Q���bɸ̥x�K��O(l\S��X޶7o�NPs@ŌM�@kgm[���b9�w=q�R����m
����)�-��D�4Y9���ږ����>2�׵;�/�R��01�ׯ� 0�����:/+���!G�bQ^�,��BJ���:{�[yfa���~"����J!m ��#�9?ڽ��8.�[jl�uSj|��W��"�I9�r�L�g���㼄�������bBr6N1⳸o7�Y�5�w��V���i *_7{�l'ƥ�J��-&^��&�����pVcke#���vǤ��jOЫ��}��4�bu��<Q�Տ0���*�x� �G8��.�d�}adI:˯>@��fr���w�����o�����[�8Г�RI���d��$�~���\Jb}�0�U�@������F����F�o�Dk��Z�2�i��v`�ޗ��:��ԫ!�M|�Xa;�BP�Ŋ[�d�(����u1���ND|o�L~�}��Vs��.�e�� $�p�h�aR_�p�k����Җ�6��&G��	{ɹ/N"�oШG�U�U�S0\�E�!�p�ܴ+��z��n����. �2�P�+(��VG��zGѓǽ�F��r���Hו��u���m���a�va?1)��)̡���	3��Դ�~�;uS}2�6r��-[��NYv꜏bɵ^�*_Ė�M�S�N�!� ��'f�9,�X�����d)��M�b�B0dԌ�k���S��/�6L�A�j�����q3�T��O��#�f��sE��ř�S�n|&��Onm��JL�9����X���~uJŗ���H=�z���̈́~Аj��DZ��_uR5��o�=˝̽Aq�;Ed�=zn�*5�ʟ�|ڠv8]���;�Ss����r���J���t�Nj/�4� ��I�y0�G3��.����Ր��/�`2��*sD7���U�DJiVe�"�,-�ஔ��k�֛WS\:v�Xq��~Y���K[<�Ep΋��)�r?Z�R˹�>�M/�;|�:pH��XM�7��U��Qr���	EQ�����.s��'s�`��GY5~�%�)m�e��y���a�AJ�Sgy/̐3�y�� L�)���PL��m���3�ON#FI�x9��0R}��νKh����츃�@J���O����c�<���c;o9��O$6z��r��;zJ}�|
��s� �zm�tX�����t.��'5�Wy)�d��NK�o���gֈ= q����G9���oJ����3tfX�xA�P)�q簃�����]�(�_M��=��9��9"���2fO�|fy%��,uZ�ne]��.:&Wڻ�UH���
\e��H��N�np�W���rBxq�����Њ|�w�������ԯ�d� :���aY�Q��$�[�喑��E��GD�p����?�1'}������ G@�����Xr���7֍$c��o�~����:x�9#�C|�a!���a,�X!�/��d7��޾�O�Gay]��+Oe�dD�����R�L��u2���Mx�0��
�E�`�B�4�-�:�4������7b%���A��Z'�)���� q��.Vw�s��k�YS�?j����s�� �2��� Mo��#e����b����?�S�v�ڀY=��8�B/K�H��z��4ޗ�h�'�gB���JE|��fA��
�lŖ��cn��Rq�ϴqS�o���997z�%^����,Y���B4���)����^χ�><%G4UT�m-���.M�|���K'�q4ՙ+���"��}$C�������ދă"k?JY� !B�x��9	���12ue�Ùf��PO8ӹ�7ӈ�ؿ�e�[��㗒��Y׀�moQ�������z�)B�ģIW�{=��לQ�A(=A�+��}srf�����πAND�&J���c)9J�@H�g�Y�>c-�M@6�zN��	f�t�e��c�u���+��aR5�Pk�c�9L�.��m�	�������GT�׫�����Qn���9-@(���E��K	��T�GT���ɣ�9�$H���N��,����-R�_��P}��i`����x���"�,�F~)Dt��~,wQ	���&��s����be�0v$��
���M/���lB��x��щx-fJӶ-c���=�����s��vS�p,��a��G���]~�?�a/Ȁ�+hVWH.�9�3��w����X��3����4�O���Um!ŗ�u0�~W :��<> �����ψN�{ʺ���1�s
0l��g��$Pt�H� 8}Ƽ"��0U�ڟد�V0 �֝{���8Mw6^N��>+2�Tiypvz�ĉA��Ym5�W��)���h��R?'h��O�z�1G�m���9wF�uS'�&�|ZH�^  �Z)��T����=��8K$�	��;3tz�y�)6ɧs��[�G��#PY_����&�ڦ5���M��v�Ǐy�s�2p��]IoD�Z��>V_=A@fA�e��,e�	cl����?J0_�0�[U�ۡ5���#���	|��	���X�[�Vf2�[&~�B���6��1��w�r��W��3����~ m����`��ֽ��wB��y}��B��ވ־P��u��",?ɪH�`lã�Wˬ��.͈���ʁ׺�Ƀ��)�U�o�l�IjtV��Wn��=�A��*���5��#!�� ��N�.�dbzxxG}O�=Z�C��3�kru��<%v���)z��[���I{�ZJ8�h�	ܞ迤+�;��b��#25�tU�a�7��i&v�1�h��eX>�0�ɰ�g/��72%����/�-\k.�/�#����c�׫E�૮�鿹��g�'�ݧa@S���9��i���k0�i�z�+Ս �*�?����P���f�pc�v�ච ��Dz���qGa�Bt{4_�.6�-	�v�F���@8�>a�!�p_�Xђ�A�}<������缑��Qͯ[�k��VI�R��+�p�~�� ��I�U�F��r؇A M���=��ōUo��S� ׆jͳ�mr݈3çkU8�c���\u���W�w04��n�'��3�����!�Vf-�^X���+�<�:���7����٪��Ư��=n���E�(Ę���^��rv"�Ĺ����KπNM��߱��!��>	��*&&���LG��A&FfU��t2�[�x֠�(c�����'W��J:$��/��p
���Ȣb�$HDoT����nrº-�s����Ϋ���͂��>�tD2�X9,�;c�f5jɔ:��KkZ��{�z��E�=�H��io��o�Z6�����Z�fu�{ӈ�H=1Caɵ�c(6��Uh�kE�2L{�%V���K�!g��t�l�����Ô�1B	�\��`�(3y}]�ɭ:�Hb
yZ��AΗY�';�vB��+��,��ߥ� ��e����/���/Y>��}��w��[�F!�~U�BPS�;�M�0�g	|��*΢p�y�M��5�	[~���(�->���%�]7TT������6&�\㋸�9�!���v
��+���W���x����q��'x6�n��	�dY7�3���l��q���jJ�][K˦5ҵ�W�Sӗ�ε�۳�����������/���	Gy��y-��$a���KH�vH ��� >Eۿ�Q8M�7L�Y����z���o�1e>�q1r��e̞������^L��#�O��f��yѻ��[�"1��1�C�L��Ma��űd�Pq�A�ʿ�.@�C�Q{ݲ,bg�E-n�a��B�^�Ȳ�� ��ʏ='|bxU����8��T�Ĉў�S�f��Q��hPZ!>iIDm����[x{\p��^;P�}��1_�__e4����t������o�F�mKb����]�1Û�_����g����F���;��[�(����(_&L|b�Wck�Њ������-���'F
�&(֋mlO��|��ץ��đ�w�4�t���
�E�W�hs���s��r)�4��xŌg	��1C1��7����������!��X�nl�ƹ��m&�2T���O�E���D���Z�9e��7���3� Gd��J�,`�����Jt��8��_���#<����J	U혃Lه��2��W�ͻ��
�j]�j����񡭄�"�"A���>YFX��$K�l���ހ��3��;�޺��|q���:��<̳.yJ_=��-*$�J��vO���4T$j���~��̠�����\���cSY�p��8�*��"&���0��p;�#_�+W�w�C�N�اB��0I��_��C����K_T�a:3+a����?7Ȟ�ȵp$�˺�|�+\���>$b�6L��a�#�\Kޫ��v��LB	�����pįS�\{�^�a�m�G��	�:Kso�n+Ik�)�J ~��&��ͧdh!�P��u��d��g�s�:m�VbH�ԛ��3��8B�x0_����'
�3i0]�HM$���������d���L�Vh��u=&3��.z�����X5a���v%� ,�F��%t�F���'�j[�3���}ء
�~������cEB�׺��-�2c$�)`��P�'��F��,����έ�E�r��#�%�m*�25u�=�|P��}|��2HcyYr���@� Sm\,7� �*r�E��[{�}�W`��Pۂ������8�����d�iTk�2���@�ueU	���d�n�r,=��ty&u��F?Bu^ɵN��AP�@�f��q��%�A�F�VS ���7�^���ۻw@K��>���rfU���߳5�J๱%��@��%TtF��Q_����{�'hY���t	!n� �a�"�����N�oCwB.����9����'�$u�ův1"t�s�h�s(�xPN�i�4,=�¥V�@�ص�E�E�ǐ�x��	z~�%,����F�:0ħZ���+O#�zP�2M,!��Y�F�D6�53���6����Xn���b*��#�N�~�ܺl����`�:����֟���w��	�	+9���t���`P�3�Gfu�9.1CƵ�!P�A����x8q�0�!x������\��A�U�	��H�$��L�c��J�6�D��4�M�r�I�~�N����h��0�͔���C��W���]�%CpMz����p�/����\�d��ш��k����l~�|��,'��fF.<Be�=OX�y:�E�º#���F	�'�Ƽ��xGT)�_����b�?'���=��ϻ�3����m�4��RH�P�I`�t>��LOӱ��a�+����]Mv=�-O���,}>�,@}NV�����rǈ��k�ڐC�aF��O½}�w�"��n|���|>D��C ���vP�3���&�hu-����F���{� �]���Im8U^�"�[�XHQ�(�aF�ӈ�S� l��weU��럎j��v~"�&ϱ���eY�*+7y]�ܞ�r_�/=��>jj�ܳ������Pj�F��lG+Ʉ�i��Ǩ�-C�0)�_�W-9���v6g�T�ߓ܈M�+��	Cz�w.Z��e���ҨБB���>"�V�#�������2;��U.YH��O_�xX-�`]q��]�b|��]F9q�?+Q�.�UN0_�K`����-���۽���W��<h�	�]s�����g;/f��w�O������,���~=}Pu!B�N�����\���׎E��Q�O�t��$�N�j*"VГ�Y�����7$��O.��{��z~��<[���=��@�V� B�
ρ�u��a����
=g���$�I�9W?��li�
����<��k3��S�9�+懳"� ؊���+:66l�"�u 0��'Q�U�v��Ѡ��҅oJQ��������w.�J�y/���e	�Q��W�'@���cf�夗�#ƿ1��F� �k�p:�"����Lܽ���>�|)!88��?��1�z=����b$�������_͔�� p�+|�v�Y"�S���;z�Α��zI+�'���`WE�Ǟ�M���<˲�u�����8BL��&$9W��wa�rKmF!=9%���(�߳4��l�|]5��M����X�Ti|�^/_$�z�ܘ�:S$h�t�hwV\�,��ȕ=���`�H!8K\[d.��_�Ʀ�=h�kb'�}Z���.�#b��=c��(�a����X�(���/m&7���U����)oߦf�ɝ���8p'
��E!��iz��7ꮙ�R!����숩��f�����F6�N�?Eh^�luBAݶ�`D����|��(1�U��+�'�R����C;1��x�A�M�?������籾c']�Y=zT���ܤ0@uëS��~#��%���.��E%����[�4����T�7�0h)�T6ҧ5��OA\���4&��
��}F ��-�*�'�DIE�P30>��0�t���~/֖������`�N��1\ND�1��)����*�{�g Y�W.�KW����c%��bxA��-�_bd̹Z-�����)�7�t$����# ���"����^�iQ�,4k�OL�6W�O�&.�nL��W/cgý��s>�f���ӻ��!���u=�K��iϚz�(iC�f$j?�mOr���ؚA��[%**���.�7_���YQ�R����.2�OM���|ϝ��Rǰ��_��;K�gY�X&T߆>4B�-��[R{��Ń�F�w�gZ@��"	5A� B��<}��`��8�	Z i�f5A�{��Z���	v,Hey����aŔC̱(�����Ne�W�u��:�-�{�V�5)�.[]5wy�Z�+��3��q������奺���|��>�ܹd�=>z!"�j���A�3��,�ڐ||:!�q�$��
5^�(x�6�a�9&-n�F�1ׁ��������I�(Z�^�1��@S�H㪸�ī�ϱ\�m� �q�]���:��C}p��)���L5�4�������������l��[�ڳ{-�|=�R�D[��goĀr��2=�e�*6�z��̺}GD�vh�d�"q��s�&��2�.�K��ΓW�'���A�����j�ⶪ��J�_�fCh_�Uo='��Qƭ�?X	.[ᵿ 3�=�J��x?� {a��1�7�J^@֞;C�,���oIH��,�BU+4n[��@z��ǈ�y'%^ϳ�c^������0c����e:�En�M�lߴ��1�pX)�=�h���|�On�>�:l��/�<��W�"V���m)�_57-)pj ����q%���(`lP-�Z䑽����+^ڇ�3P8�����A�[���/�
�!�(T�;����w,r1�g��q�v����^#�����T[g��\x�	@��nN���:O�t��1����8n�(xÙ���n��{lR3� 3�����qcZ�SFr��x\P�����`kH$�Lc� .�= T�aߖ�^2�X�VtK�s�9��c�A�f��J�ݶ�cۙ��4Q����`�vy�.>I�H���m�K�r�r��%Ȼ�;���DB\ĸw���1 GɅI�zh~F:�,1��e����Rp�Aw�?�B�4� �ި�[�˱HQ=�m���d��5��B��uLSpVm*��P��T�D����Xʢ
���KOI�%�*��o�u�g6��2Lݘ�o��;��g(ɢ����WT�/��H)f����p��ӞJ!; Ѡ��8ߞi�]{��m\I���*�C~�5���6��O2X`U/l�9�HdU��%�xڴ�ᕫ4_߂U������nI�2NF����:�"X��ۆ�pfz%�L�0u4�q)F��3�"XK��܌y�j�h�x �Y)z�\"ju�}�\~"^@�T��
~�?B�h6f`�#��SpV��)�:؝fգ�<�����BG)2������ �0#g����1V����^����U�<Zq��O#7�]s�IK�ӛI9��yW^d�������7#��h���NnMT�z
�_zN��B�Qߔ�M��ܡ�%���)�+��
F�r�(0�z�J� |���}���iT8��e
���N#��[��.i���E� �B-g9 �U����)	��H�v6U�K�B�<�_�m�BCQ���[	�,���1bؠߎJ~apPҫ���Q�&�J�9�%/��2�d��a�ɫ��:�	�|��yK�ME�V�����|J�M�����ІI�JT$�5��A���-F2�aaiE�֭���g��&)k,Yw������ϔ��$�i
q�ಚ��\�x�͛�Y<��&F(��üTk�>nf:
X~sp�5�ia#&�^�����~b�d	�pWaC=\J��@c4'%~vU+���O�J�M9�Y��m,Wq����l��w���
�sW㱖]T:(mqL�ш�R"59T�47�����+:��5����ܞv����/B��0Q��j��6�[��� �l���O��G�k�⯨�r���@�����<r&��;-
���]l��H�du��&X�������>=�_���{�V��s؝i�&����N(� m�����zF1�@��'�VI�2�ɡ	PJc���<*�ζ����?E�N*��є_��yӿ9����{�.a�n�U��0=7�\u��ͱC	]��W�h[-��?:���ڀd�*P(]����C���$i�i�`��v2���\�L��F��bb���c��KK��+%��b7�L�iN��F��)f��G��r��M��ǀ��V�����\&�	w=��ɩ|��c��,��K���&�� � �%��s6���ZX��W)b?~M.&N�R�tP�L_��$�Yd3��yјέ�vLᗣ>����p	�
���Pf�q��{T��C3�t�|G]���Ԧ����Gq'�y%�� �f:@e%���<��3��۝�x�D7�M�cX8�,�M��q+�{ـ5�m���<�,O7��L���瞢G��E{+�d���Y/Vjٌɭ}�S��}D��4���AP� �Y�d�n�����"#>Z�n�\t��7Pc猏YQ1���B����g�P����
ڲ{]���F^�B���#w�ي�h���?0b�nt�6}ߔ��,�2�%i�ᾂ�Xvi�$��ϠCv��B/�Lxe�Y��o8�J�!�s����.|u���|��7�;.��r�PcLSP)r��
�'�e�0�}@܊P-��'�"
�o�"s�f�����Ժ,��\۞qj?��/g�����g�YsX�L��g9�+ ��/t��э�[��|�?�Ζ�zK�t�����9݊Ҫ�Mћ3[�[B.f�UL�Y@���-�+o�N"=a�^��qqd�F�矰[<��w�T�)N�/B��	�:�xOԎ�w�~���B�r�qĴOǢ�W����O8�p�l�.��[.����b�V0������8�a��0��j���1���rdqGS��ۀ���U��cmޟ���11�ue�d�c�>-0�y9�2����Z�~䣾'�����
���Iږ�Qr'$ʒ�������9��,A�U��n�T��k��X̡%'5^�POb��H��6h���Ư�c%!� "�u�T� �^�G�2[<^�`�kQ�z�����qH��OV�����4\�C�LO߾9���M�%A�m����s�x��@�KK�������Q�'������s!���`�X���Oޓqb�r0R�/���$}�U5A�8�V��L+ �6��77�Y�k�����=�b�+��Z�]��a���+Q7Zqʰ�9n;w�踦�*�˓�5�<^�w��=����S7	�(���v��Ý���zٱ�(���\�n�����+.".*+v$�2�6"u��ҍ�޵��W,�5Bzu:5�0c*Q%�I��]��{�XOz�������;���vt}P���w�~�C@�Y���ݡ�*[�b�b=ω8I�3F����M�?(q}��dQ��>�l{���fm2+�D?`��ֲ7D6[,������r@���I��$��}�,b��E�H���{�Z���%x��iA�Λ2��vt	n����mMIU2U��<ojhҝ֮�x��� ��;��԰��g{�)���1��a=2��P�P��p̨=Mݞ�R@)�|��?4o���/nW�U��R�~�C��s�g��MZ���>PDԁ�:�V!���E<� �Ld��\�Ig���2�Z̓�TC���]6�Tm�!�A���-w����r��U"ܞ�"�<���?d�Y>K췏h�+r��ycLR@��zzA%�ҢE��P��s�So�=ąZ��ˋ���/̪��J(�+m���un��thO@Q��Lg�A��<~�l��c��
�z�%�ӕ��C *d3?�,�Z���C8�\T���K�F+v+����@/��=��1[	Tg����Q����+�#�O�q`�q3����q �!>�-��d5�<�=Z��]r�6 �f�i4�=]�G���A�2�#�*�d���ժ����U2��6[�c�ơ�TI	�m�l.�BVi�Q����,�2
�����ֱ0�b�f/,$36�e��I���V�N)�y.C��Q��ӵ
���/�>U����y�M��a$|�����ks�4�T�uI������;�#�8[����	�|�'�/<�7�0�k�����v}��=� '�:_5-`ՆuN�ڊ��)�l��K\�R?p � �z1�5Zp��EZ����H�ȹb�t��F ��E�zc��Y+�� �I�.�nJ2x��Z�C>����{�����nJ��+vZ���&�I]jؼO(:�l�E��gM'z�c?	]+rX�|�fӵT��	� �B�5 l��X�|��{�d�aZ
�+�+j�����u�nf{���>�$0��]?r����6������(���͸Q&T�:2Mj
x��q�zʢ�??wO��
��T�Ё=�x������B�p5�F���k�<"�� �j:̷�KB��wZ�S͖�/��f$��Jr_�'����G�ǛH)����P@�фxd-��;���v�XH���߯�lR�	�"�C�x܉h��H�X��oϔcj���i�j:۪�N@C�.T
�������+��*����٤�8Kޜ1��j��^!j���m��h�~_������Sd��h��.����b�P�.4���g�#��_�V�>���qv������	�*\�5�$Pn�f�ۭ��i�[_�Ce��G�����W+t,��w����Ϡ�6�U���TR!$�����!���z����D^o�!�!�a;�pW���>�T�.��q:�cr��"����l�3�HCB�dkgX�7g�1\�pa�0�wu�p?e�`c��c�a����z�0�`=��?���QA 6��U�O,5y�N��IcJ��(��A�6�>�D؜s��dω�c�u͘�"�4P�J+u��_�bc�5*D�Wa���!7:/.B&�� q1K)�?jh���8X�:t<O~N;n�@�3�CSȚ>pĊ%�*|nDHݬq�$]tnO]\�1�!����	6)�����,�*Spn�
q�[A�ajQ�]`�w���3�o�u��;�.��'����n�*N�}z���'��
W2�����N�`ީ��=��&ޚ4x��e���|�T�^���n�7����ILܮ~v �zP/�oc<� &'�h�}M�q�7G~n��%!hb-�򷘯&\j��D/����;1ew>S Z0]$}%װ|b�3;����8q?!.�tZ�p�zk�w�?�a���D��=j7� Vr�	�E����XY����px6CB�J*�p_"��0�.�i5�̃J{!�0�<���t��aN[�7�'�(��ceaѭ��VA]�����	,��T�B�/N؊X�xٕ�she~��lH�\�%���e����o�v7�s}�Ц�M�5f�O�d>#H�3�$K�_wVd�[�Xw�����P�qm��Z�ޟ��w�vBH���M Ct%�� ��̓�rd
�m&ـa[�B ���qu���	�����[��6M�)���[�."�м�w�a�
J���h��'k�따I�����ʘ� �q���Bo�b��({̶y�j/4�-6�>5̫Ɗx>�t��n���S�4>
yp���@��[C/s6�9.뽉�Ɲ��TT��~W�D�=��܁)�-L�z��2��і�qd��d��hѯ`���Q�����le;y	�&ͅ��%�Og�?���z��xK�sF�|��if!��t˝I��}���>�yC�At�gPRP�����E�ȪL�9��'{��,�M�y�}gPI/��O(���8j�,hj�����܅��A�r/lc!l�XFR��n�)�-��9D��gi�.�f^oD��7AZd������oδ;��U�����k�%�ҷ�M����&����@7B�]]�(��|�d���;�@!����:�k&��߭5��L.���?�8�W�M��	��A/D�Pxc�$+�ӯ����W~ۂ��]��x#H"ˋ�<ٰ��X�\�z��K?O8P�g�k�P�`q��n9��C&GzSmK\=�1���_s�X2|v��}��r��?0� ���u�19k�H�۟r�ٸ���y[��R�+J``��W�\�j�~PKC�m+�hkLK<��˴�����C'��㼒�D�����
���$�#>붳:�r���ƀ�f�,{��E�����\�z<���t��g�i�~._�\w�
��ȳ}�q�1~[f����H�.1+`5�M�>�8ր�`l"T(�������do�e�A��Ic��D�bu���z*�Q� 3x*쫡�p���c��sJ�������YS)Mp׻�C�/V��W���7H�^)_
�
�,`��
~7��i�#c+�W׿��b_o�P�������[ܒ�c�-fT�Y�E&@G�0�� �]ρn��'m�E�w�?[�W腉�`m�h���"�65#��ˏ����ߪ�6��C��A�8�a��/2��_ӪڗA������vN4,�q��`��,��n실��=����fv@���>ʇ�?�zc8�Z�gF��0p���t[�gk��q���ϥ�����ɕ��5�*�� ��o��⓻�ϐ~�����g�ܥ���C7��)W!��L���� @�s�d��a�V�n4�r�&������� ���M�Y_�$
j��L�j�Ւ�Y1Kpz�l�H�WO��cor��4_U%Y.2��N�M dpn��瑋��6Q�C"���ɔ�@{@���"[븠���^:qĽd��?�5��8ؖ��4}�L�����+̸d�r7�~<�3�oCjK#w��p�8�Ŝ�ٴ-20�^��NGPWV=�<�M�ڡ�Ob�b�|~-��ȴ��:sT�k��)#]���)�؂�K�):Y�Z�-��]^�Yy͈o�iP�h{��6�ڦ��C���M�v�6g�<�Rh����!�) ��?o��mB�n�F�7�c��R ���Qf\� ˽G��w�����b���s�[��)pM��sr������Ƭ!k�ql�q[����Tf��6u�	��T��+ӽ�"�ș-���#���BF�O���#����i6�]|���������{��{��4�U��i�!'7F��^���a�^���NW2�π�:q��36��ė�UR�}�ܶ�	��(��O�N5���Fгðil�TGv�ڧ}���,l�Rb� o��8,S=a��W��x�4����Ex�fs�2I�ImH���q�� o���Ħ���^�IS��f�%2��^Vޞx8a/p��d9+��@'��/o�5_��e"�U�S��9�-v�o�3�y��q|Q3�8f�~m����]��5�!L������{ls9��ɌB�έ��Mp��Z��L��1(���擡V���4���B�\�	|Y=Hi[i��*�k��RC��2"�(�M���e��y1���� Y��+��C�:@'ۈ1t�ط��at9�$�f�S�t�C��
ʍ��C3.M�����6���(ׂT˶�iMc|%� �����(-g���i1�d���G_��B,2wVD�:Z�x�b%J=pT��=ڭU�1h�`K%�"��|=�j��N�YX��?B���9�x�=��v�-5���WyJ�q%��S���� ~8H�Ɖr��9�F���5�6i�����0>=C6��99x~��!n���f'w�RNbܳ?�]4�S�X.s~{3�t��6j�8ޖ�Cm3)�f�8I�鎆3��h�)��c0�{�
S1����Ql^[e�c���U
�z.���g���F��b0ӿ\�-�H�D�[�ѥ
���>���%�Q�C��k�cN�{�ӟ�@�%��Sb��}+�9�a�ƽmQ{��0���HQ:N�h��R5{��$^̰���g�*��6����,���Ky��q���j�G$�X����ny��9��
[�UI9~��\H���!�M�6�Ҥ2��"yn��lE�vb�ȿz��Vb����Ev�]>�ŕ� d�+2AG����!�R����N�ɼL�'ݢ1PA2�
Ƥ�k��}�	��m�aF�ˎ+B���7a��|�~CH�)�X�Ύ�f���ѴV�Y��I}}.��ks�/��D���ٸ���o3���Ҁ�,)@�,���3��O���%��PU����9S�T��v��P��E�#��2�P�>�O�\0�8�o�Q���-���q��=T�`�=�����z�3�W��CiR� j�:��$����U%ځ���3�d(�A}7�%��vM�(i7
i+B��$i�Ӆ�t�a��Kd��C�� M��P���S�E�����&H�>w��t���%�����F�Q���M̃B���L��9�����^rۜ������ܩnMYkHq����w��_zX�%Z�wQݺ���C��N�'�N�ԋ-V�9��L����{�\�<N.�JG��K�q��.�����VjR�^ $-��ᮋ�Z��M�>�����܋�	Mѳ[~�������@��$���h$����/��]�V�;p1������}ޮ�Be�N���0[���C��6/�'�w�,K�%�xBŬ�0 :������1j���U �� qspD��Z��U�0u����C�����Z3��y��v.^3CjD�:@����J��6�)��+����#9�!�v�����.�*���8�����-�¼p���k}!,{֏�Z��Q"�A���XR�^mf2q���Y�uW�"�ܯ|]�l�̪�D^��ٵ�UI���ص�zKm�c.���V�+P��υaw��_l�r���C��������~7�,�l���~$���c�@�S�%�	͒�Cm��ji3�S���|��t������~�5������f5�l���RZ �����am�����U`��W	,\�{�u4����D��G/�z��JK�H���&ۛ�r���ڔ��q�P��4�cG�ڽ���3���Y.�s���}{#u"�h5	;)��v��ˁ�Ԥ��!�u���Yh�F�K��46ɯa0�}�>��a�NQ�K�W��G�_��3���O��1�4�GR`qQBt&��>�iy��&�v晦��`S��xO�_d��2^H�?�Ϋ�e&�P��e�c��������Ea�^�e�t��#�Wݹ�
�-�YdI����.��L���(29Y\@l�*��V1�($��v߳������X�Br!0v%�i�@%`}�Δ�����
��Xj�,���-W�u�/G(���7�mtɸx@�d�?�(���������I%���U\\W�u���c�_�p̟U�/���,��ۇ������RNT
��h���=�f������p��9I�3��i��o���U��$z�"�uy�s�~#�k2�Oxl�4j��~�1�\��x��BW��� �ǹMp8=U�5��^�#���&@o���;�`\F|��[H?+�Bφ�&�.��)p���HK��<#|�����s��+a;������� ����H�8��]�{��gNvu�$�=�U�:����1R�l|-.P|�+�!r+|��~��V���h���Wo�nWw����6?2�{`���E��Tcވ?S�Pi|�R��P@y�E1�=�yud{�u��%L7,��y�Hv���#!���w리��bWI�E}��c�-��� �B��\�W �6��Ĳ�*˜H8rsL��N�����|�N�׆��C>�%�Ii�nÂ"خ�E#0>gIE>.�N8r�n�k�+�n٘=
Y�:�egZ��k�D^Q-f�wZ[?�EQ�������w �~Wy�~���p$����ѯ�
�[A�D�W4�p��������,F��G;��oG9��G����d���fJ�=�RFZ�x�wNVhiBg��j߻gD�Q����	����z�����f��j��/Z�#�Y	����c�V��3U�3Ǧ��fZ��h�t+�i��L�'���k"DcHϠ��*��)��Qla��3����&��E?�����j4:xj�����3k������C�t5�i��'��E_�%��X(/�T�Z�h�q��Ĝ� \�q�X�w�.cZ�~�lO= �k����G��P^�sĪD$���ނ@wI�'��D�1���;M>���Д�`
D�Р@h2���]9�;��V��ꌰE��'����f���ij �Э�Y����Ic�5��L	z?0��Ceɵ������3�5BR֛`m�a弅����X���ed	a�4��!�]]7z\r���I��Յde��5�p>�1a�n�EI	�2i#s}>W]�!8�gh1�j�o�f.�Wz�����*�$���!���1�j���Y��EQdv���nǠ׸	�"�ΐ��qK�\>�^di� �����B~���p;���x:_�<��/c,v�8�A�ӊA 0.@����+�Iu�u�U��@)@�EW�n�]�ٔ;��"�^������/�L4̹6�ċ�Q�4�Y%��
�6�G5��O5Cw���ɠOޮ ��
�D�C-E>-6�?`P�?n�F' ��R�ge�Y�^|��#����J��*{o�@�Q���y��2��[3h|h'���=j����Ǵ��RT��H����,/r������ L��vg;�$칽Ev�`��<m,	����Zʹ�6��jڟ�-����q��caJ'�Y��mݿS�	Z�N�"��`���f�^n�`V�ea~xW\@.L�&�E�����O�Ȭ�\ޭ����}�b��T��&�e��G8��F��F7'ӛ.�4�.f��r��T��W��G�`�&����,��L�ˤqv���;���Ve�u^��Ʀ��A��M��Z�^�K+�]k		.	��eபuF��hM/Gc�֒zL����	���GlPU}��ʍ�t$$o�!�ߢ�7	j^��T`�0O��-��}0"��mG�O
_�=Տ�'���Ao�-"n��*�FT�;���K���L���%����_^�B���$�M3v[��;���"'^�;᪆�E=\�F<�@i�	�s�Q���v�_�ײZ;3���U��<Ɍ,���]/����N��<`�����6��d�.�o�h�	w���̊C0f!%JFkw@S��᫞#Q� E��>]�bI���0c����,>Z��C;�-�g��|�*1}o�H�I(	���J��^.�C �V��Hx X���x)X�=����
�O&Y�q]�6�!}��[�g&���)��}l��\-E&��������3��U�Qh֛�+�|u�p"���>������^��Ql��-�^�g:�U����ۃ��z�"�a�<�H6�!�چ}�=+$��V[�P_ۼ����� ����� zv�s_B�D|+K>�.��G*�jR��^�޹�eB~�ǒY��a�Ϗ�V� I�͑��m
e���+UK��]�y���Vx؎������