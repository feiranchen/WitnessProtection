��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g�%��'���s�V�1�	����'��.9Ϧ�R�N�������2X�F��1Ui[*��L`���~/߄� �b���
eKŪE����,w��� �̆F��I�@�x�nƖ�I�Y�,�ȉ���}��F��OsP%v��x� ���V7��?K���S��U�����vO!D��$v,� o�f>��� b�f!���n�Z�{��I�9 ^f�ǒ��y� �n�eA�������Ʃ��k���HD����d��p���~�HbY�M[�@1���}:pm1L�Å�⪸U� �#��b^ur��sB��q�̙�:mZ$�7q��yR�������5�#�k&�ل�Ĉ�����M�]���}�s�p/�w8��XGd׵S(���(���%yx��0��RƳ硓�-ƪi�(efq�����ǿ�c6xm��b8]��p\����S��v�����Jb����3��_�l��9����eB��A޽o6���Ԙn��N�?��j�^�rJf+l�%�bH���5��)��`X����Y���j���e>~��b��:r"L+��ߔNV�{���5�}l̯���;� �����+���&�f�!��>���3�rjO������b����}z���W�`��\e�	�2��;�v�]�C�����9,�h.�.	�OV�ĖD9��8#]�겢>�^
7*1�^�+dt����g{��8�*^?Í�9�9V�FP�*�B���Q�[�������z��勣�S�:��[}��]�|��s>GqX�z����-`�X�	�Z���g�yX}�;�����;�\H&�J� 9f(��
��]FZfCY��4ba
�k��(�3M��e�N��N��F
Gk����2�A��]W܌5���e$��,џrApw���3�`���������X�i�<��3�y�U~l�)���x[ԣ�M��2��RA��i������3�:�{�>]ʹQ��H>���s�Y���d�6*Im�/(G�u_Kr�@�ك��¬��}8��5o����,��� �5�ځ�bU�~�Q�DuUQȄ����b�Q��\ζ�bB��-�[�I�S����>~(�Ú��k�����L�sV�_5]�l�-шZ~T�ߤ�m�2�Ґ�F"a��H���`5�V��
�90�D�'+CJ�� #���<��MV8a�Q��e�*]��N��I�?����P�#�P�f˸��O�A���(ր�q]ѽ]w.=�����~�HD�&�����~D6-T�?)����[�{8���#��TX}����h4R�*q�N 1�M�]&���Ev_CR���5��M%�z�	D�
���r(ѱ�X��Xn�����)�P�:�����ۻ	�˵���OL
7/h����ԗ��'x-�	a�I��rs�Jz���OI�����ʁ}�zD����{�As���~�}gXԄ_az��*�1(~��P���˷R�FU*T��[��w6�C�a��;;�{�;o��t��ᐶt�m���'���G�wt�H��rU{�%��Z�t��v����83䖥a��1� P�
B�0ȑ��z�27q�pn��"���>�_/��f��YG
��������|.��!�`�h��H��Z� T�(�0	[!�����_���Œ�K�������_�c�a�-��{��aSr<7������x�]az���z	��@#�Ɵ'_�X4�g2a.��'��ɿ^ ���Ɂx�� ������_�U5��A>\��upM�������A��剒)�� ��*�s���JQ���s�9u�����e�|>�H#p�V8�nE �PX~'��K-�������KX�L�c�E���v��F��B_8w��}�ɫm�"�w�Y�(*/��B����T8��`k���`�gջP��k`�NI�y������aQ� h��64J`�R,���6��(�ĭK��.m�� �N�q8V�ʗj����#��h���H�-���pg�������n�2��Suc�x����R~
���ç2L�:�x�nSh��q�5�헗"/RT&�ʕ�����G
#�1��&���e�u�h��$��޵�5�k�l�V=ޖi��\����m�K��.emB"#9QӮcD��m��O���p�<�*96
f�e�;-u#!����-7��������7�<W(�#Hv�`������5�Ɍ��Slo��ڨL��~5�Z��"�H�5�9N�.lH����[��O���y��t�|v���|�ި��Q��z`�_x<�&�al�!�d�'�z�	4�utw�'�Q7v}��e?��>&)�Z�V�������g��l.=8��-e��]�����X��:����ah�K��\0f���!�� ������`�&ebDǗ��y@� 8�OM?�c������m�|�u,ĭW�X�D�zs@# ���?��� ױ�y9Y����8s'���
Y
[�E��*�7��)��س+���q�@LvT��E���e�z��1KZj���S��ېC��Q���3�'�fu��Lb��A�n�s��� �m�6|	�V~c�w�8k�&�2D��v�m&�a(+��;::8�Z#^W�F3�� 	-8����n]�����;*=ʭUM>��� �/�>H�݄��m��J���%n%���i��W)�	Z
�&�����y;LE�<� D���Ҵ�xP�w?5i����-h�N[� 6+:�����9�DX4ʜB���6:�����c��ԛͳ���2�wC|Γ�i|�&*���f�4k�~c6�1E��K3��BԀ���eV�>�L�7��Z�RzKo.�G����:&k{B�Ϻ��H8�"|o@��۫�:d𜧂��2� �K\�E�M����"�:�"�%u�+��;�>����r��5����鍜˼���%Oh ȉƝ��FY��遣���z�]Z3W9�'������N��H�F�͖�cM-����F�'��������g�gC��'���a)�������2\K��@(g��T�=�.��˲�D�$���'w�΄1�mȐ_>�I�p��������i7ʒR�����r�T�#�(a.3r���+2Tq+�Թ�}O����y�Tz��:I2zQ�p,l;�⯳�ZЦ��<�;����@ؠ.AV�V�oH�}�5��)��&i�-J�wt]�D,�ɵW�A��OX�c�n���C�{)�3�y�����]��0���g����2�x�@��H��X�ǯC�s��(���<(�}D�C(��z8�p��d ��U�����K�#gU�F/}u;��	�9��-'7��>�I����3��W��0J�.&�� L\�{ŝo�|��̇J�&���NHX^ā�Oo\��{�4$�_��=tm���l��W8C�?���/s
Y	����_&�������o`AP��~w��b}�0|N���}�Iى@�� � CHX
�>oI�����K��)� Vu]�>����e�\�*1�M��f���'HsKϥjF��݇�ŏ����V
ʙ�����'�� �ux �l93|�䑢��z�[+Qq�s�%�gJ^���DNR���ʫ)���o�7v�$g�����}��y�z��Өw����� ��oeE�@��}�xPJ���.1����2!$8���׀$Nx���se�ĸ
SJy�o�2L)�x1�4��k��Q<��)9�A\�VDezR�,�y�d�#�8,T�3��c���i�E��2VzhNq� �/w9��94p�:�z���*�
Y*Q�66u,�._W4M��g��0Wމ�����Sj�@r>�a���a}���q�d���-����Os�Pm�o��N���n����
"M���%��-DF����^�o��=4��Ǧt'���N=�!�m�87����眂`�������X�4:��-�8*F����Ã%bo|�d��
�m��Y�U��<UL~UW�}{B<��,��t�K�J�|Ώ�iENP7��~[�z�t8_������8� �y�o+k��v����MCr�-���X�!����3cd	��,����iݴůX��Įh���	&����R�1�}m���l��BXN�ʚfUvDd�4v�Qm�'�������6�ڡ�ذp�����e�A|y��L:�������mS`G2[z�NQ��㡏��ˮ����ڈ�Hy�XW�E�O��v�t�`��xB�v�"uف�x��Ēe�rw�j��+�m��+8���d�����%��R9��R@��/'��y���L;�
j��@���.��A�����ݐoz$��&�,Z��F�~"��A�c�X�,�&�$R[�y�<NϾ�]=��Q�#���8v��~���]^�m�90}\:`r��D�Mϥ�v�~3KGX��u_��4d���>��W�I	�"ܤN��oLD����(��dfe�ֲ]"~������e��w����Q��� �F����\x(�l��,���V�i�_��D���p�`�ݶ�e�ٲLy�y�	>e*����˂�@�б��#n�_B+;�5�1�VY�&���XFqk�� u/���c`[hZ�<^�T<+V�K[�'��[Z-~��Q6;���r�E���F-&F�тp/������H�(4X�	Ws�T�%��2����,�A{��p�Դ�� N�RD햂��
�r�Ȫ�ü��.x��]�f�{��X4|+�3��Zd����
�A��Y�����g�x8�%:^4��� O��7�$�a��q�@*[aU)�����B-�O*��7R*T޳x{��U�S��~�Uv8aʄ��~uԋ9آ �Bfe���g�F����<�?�|FѪ@O��o�;��(�Y��G�`��B���M������t��\h�X�8b�A?�(�s'�T�����]r9%�L��K����v��ð�I��V+jҐݺ�Y�.S}��D��P��)����h���u.�	�|I9
!C��J�I���Q�)�#(��ZJ���>���,�w���F�����*�� WdN�E����n'�YѪ4M��$��dϪDn���^�=�����O	���˘wBnme��-/@TV���)�~�ZF,��8��
!��Xg@R8r���BYk��շ$��V������69�� ^y��%Z�(ȳk�q˿)�z���ɺQ����B�C��a��6Z���F��©�A�p�HD�2`�q����c:#*�O��dxṵ�O���K�Sn(����L�@�6?FMS|@�L�ToH'�0����I��oT.���	�Ta�7}��f/ߑu"h�>���2-"�O����Bs��]h-bb��ތ>�D˷x�"ԒU�Vs��M<�T5��$�9쐠=���� �?���M��юƌ}gn�vVT2���b����u��>}��D��苚���GA������{�<����j�
,ì�Ҋ@��Ϲ���@&�}�����D�����IQ��ݮ�s��s�ш'�
��!�})�me� [ɫ��ұ+\�j�Q��i1o��t�E� ��4�+N��6�t�=��t�s����\���\Qw�>$�@�ڰ�C�}�)��E`�����I����6�I2aYM�6�O��ˉW �`h"�U��V�t,۟��u��Sf�-i�9�����N˟\����	��w���QBO=��+�2�w�Wl���{��/٫lQ�������Y� 8����+�����r�;A2��<��ɶ✆�.����UM��U�0e��LKȉZ��a{�Y�I��G�	O�Q�9���f{Nz�}aOo���U��:1J@�<@�g֍w�4,A�"������g��$e��I�c����{�\��_I�کq��sb�`XQɿ0�$���L�j��l�>�oGJ�e�H�:yJ}ukQ��iMq�����y��VM2 iOAZٜ��hm,Y�g-�h\����?/�f����䦜�p^��P��j;O)8��R�"P[���4����g�������t�ߛgtȑ�E���aT�߉�y��p�`[=��1v�'����~�x[�w�#��H1��G�?�᲻�3� D�9��NAE.Pkb� ��#ζ���fG�7H�rgL���*`�7��q4z�UC�Vbm���Pw9����M�.���ݸ̂H!&����sI��77�S!�!�T������-��ٖ0�ZjB_\M5��W�yo��,�F&s���_�������X/|��;7l�̯N��1Y����ia��L>K� !m�#�o���=��|�7�8q�-ָ�]��2ɣ9�g�/��}?���G�ZV�+~8�Ӕ܉��C�wm)��T��ۍ5-�&�������6U?BK�����
R᱿A[�FY�� ��@�	����V�d\o�����4 _�!�B�,ǖT�[r�G3h��ҫ�����AmJ�'<`x�:�B�ދ\��]�m������>��炖	0�*�S����OKV�Qʫ���!4�I��EdG�l�Ě�3�ii�|�C�򮣫�M��<��� `fKc���ԕ$�X{T�u0�,�c��� ;�Þg��m)�)�vC��b��9GZy��M��Ga8�
���7gd�����\��
-]�����/q5�f�����v]W��#��C�Q��-Ƶѳ�\?}a��+��Y�i<��-<���
'n��ٱf�נO����oן"d���UJ��5��r,]�t!�f߯<�Dl�:d�Y'��7d�F��lkB8��g��d��<��Y������.��S6���UY٨�H��w����FU�U8/�`�����0:�L�g-�+��ۊJ��IM�2�x�+<��c�Z{n�&D���bw�A;A��o��8̈`2jw�2%7�d��O ���J��r�h��@�D��M���0�/|"��?cU�򵴗f�N���.�7�V��z�d,v`����1�,#���fs�蠻�K:�S:Y���b}�gR7s����3�3l����9��	��a_��=�7�ِ�%6	�>-}J����f���Ȏ@1қ���y�#��ƶ��~��}�蠻i�H��k5,�� �5��K$*�J��`j ����UG��]|I�Zɓ ������w�7�#©D@�GMs�*	ޢb�EV�̈́(��@�R^�h���҄�*�u�G95)���D� ��r�������}���8�$�zT��཈�o��x�0Պ�U���41���C6����8���n�0�)�����s�)CDs�f7^S�d��h>����ƴě�%��]2WW!�����5�ʢ=����<!�>L���� ���'4X*&MU=�S3�,�ʶ�=�� ��e��]���2���=�kc�z�HF�����h�V�U���$�@YCp��;�Bp��j��O^	L��C�Z��!{J,ғ>�F*>Gi�[`/SP�F�Q�M�j玕�-���zZ7��A�JN��G�3�|�H�Q}�:�_�F�c_v�d�F@R���Y�6]�n1�ـI�ea	$�8�5��MTQ/��~+%�iK`b�,��U��=��YE�� �k�s&�s����b�u�Z�pϗb�H�ԯT��e+ͦ�|�Z�:��%M�s
�ɘ���GJ'pA��#tPo���R����5,0�RY�0.?ꦼ�0,]ˣ�t��J�Yh��I�S?:u�	S�a2��g.��1`���{�9A�䟪g� Y�}݈�� �
Y�"����錎�w�i�PJ��� ���"�b/:� �7�����e��W��h��=��0�?�]h��(
S|v��׍��8x�e%�S:�&3���J�����KM)پg��/�;w�26���w��U�k)f�cO,]�c�������xX��4����Z��>���]��	��[Z�;n_6Wi��~ ����Ү�tj����xRqAwfWp�k-P�P�*u� �K�o�(�]@5����؅A"��D��vl|]�:r鳎]֗�������Z)#X�.io�����4�m�63R������Ŧ	�ƲK���_A�|U�˩K�A4H��R�B->�4���]`�T
rLȽ»�8��|]����������ח{��|�e*�̬EYC���a+�2X���,�U�vӂGˇ�࡚[@9�̧������l|E���٩eX0<�J�@��j��kJn+�{�!���Q�#SHB�/v*4��3����\>m%9ۇ�װ��*�5�f��Nؿv����w9�n�5�wv!,��m>����9&8��_B�@c�@A7�.�Am����F�ߤ!:�xjz��U��ܣ��R����a�R ,��/��e�����Ca!:o��O�H��-W�[S��g��z�����;�������Z�3�gZu3�Ôb�U�W�����J&���`�*y�(���2vt��>��|�,�R�fQ���~e�
�j��	�L�ܢ���3s3�Y�F�6�Q���8*����i���҃e�h�$�Ox���ս�u�~��o���Ѣ?9�WD���2�8�}���Y{p�a��LF3j���:�!�R��w�/��S��9�( Å����g!w"=�X��
(�����ץ�r���Q�`�J����9�˺S�q9J.���$��`ɜ�B&+O
�1��4�p�(����0�AM(�<��%�xh���06������/Z{#��������=F��Џ�=��R� ���ΧB�l�����H��/���uBuD�Nh``؈5�>b�9�',�HmEwfa�؍�(z���I��� ��5N$Wf�U^ʌdOv���DvKt�c[��^�� �s�u_�z���B��,����j`������΅H�ӊ�hoc�������8��\�y���	H5k�T��iN��? ������&y��c׺��L�  �_�u��˯��!�v{UOv�%�m��ȭ=45DsIr^<�f�M���Z�Yn�S�MWH�^�(�C��f68o�c���2��&8���1�>������Wg�s�kx/w��^H ��c�����ZI��M>̥V�.!;����6��K��wV�Ť���$�Qq�G������/���eqPf}���#����������춈�z6:�����_#^~��{��|�w�ݭIE�я��::��X��E�@�/E�޼��u?g��@�ca���D"n��<J���#24I���[�z,"�T�W�Ӯ��]�ʰl!%.j�O}�s6������w'^��w�����