��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jå���s����ք��4��MX���̓&Po�.���iI���-����q�R��&��Ԋ�,����m�au���p� G���j���P�����@;	�a�l�N]�Z�:�!���Ƙ�`�R8�;kC��p*x�l~/8պ��f�i}����(�|gC�(�������oĹP}C��� �ZF�����|S��M�	~�7Ԫ����twg��?�q�D��Ք�*\�^��o:��B&�K�!��2�C~�z i҆����&C?O�J2^;�Ͱ>r��$H+�ذʽ�̟G�ݔ?g���J�Qz���#wBI��ͷ��`�z}�����#�b|�$»������zF���	���)�/������}{����eL��d�L� 0
�ժr*��eI[-�|�x)����Y���dP�hQ�����y�(�[ȁ4A�o�g;��*����t���'Idga�!����W7K#:u��9�&�|��0��V$��p����I���^��,���#�<ң�DVӬ��o��<���xdM��VMr�fOK�=� �8XП(#y6��y�����/ǎn��n�~�>Dn�+�?K�WG*��Ȝ���MŻ��T������{n��S����Y��(�ܱ6lJ�VؒS^aE�5 (�;���H�b�VS�q��K��R��8��
D�!0$��{�86w���G����z��=����
u�0�d2%=5���
��)T���$��c,��˔��L�`���Ё�[_O�>��2"%li?�JR1��3�[�$S̟@Js'ʰ� �D��g��\��M ]W���%!�.w�r��!z�.K�;�Mz����l��x8�I7��6�A�N�f����gq��О��Ki�~�B�_G�r^������)3qr�M�I�'�@%aO����ǲE�g=
<��,c�*�OX7�����8�y�`�����COR�G���bĜ!2x��
V#	u�rT�ҡ���鼶�ƻ��k��.
x,7���q#��M%����guԖMs�����(2n�a�S�*�z�"����I���X�ւ���JD�_]-Y[�`0����y���>h!�A�� ��>����xZt6f�@��_ة��d{��O=k!->�!��+�i��q�a#w�乔�m��?��gVd��eݐ(Y��9�H��cGf�����<�S4�v�c�a�\�c?�]�ͯ�eɌ`_3	��#I�H�$^M�N;ꗟ�0����Y�"�J��T)�߽a�Ɲ�`8,Y]t�"�Mp��~�>ڄj�����S+�r���l���N.�v�U�'��8&�7�z�&�f���ZtDF�qDO�����.ɩи���k�Z:������`4,+.f2/��~�j��8@�H�v^�r4T�P;���u���ŝ4����3�U�Ђkh&(A�W<�":4H�[��.�BQW�[�C	�Ð"<��˅µO�W^{*�{,B.-�:���n��
k����ʞw9���l�6�\C������x��Gh�3;e�N���x�I�Qq��~^�'ȇ�[bMRd8��2߆�϶�����5o*E���8�*��/=d�F3�)��J�zF1��k��\�&��p��s-���k�gBx����	��C�->D�H�	,j!�缝�8%�f2�|;1�Z�c@�s����F�5����edh5%}����6�2䉲~S<W�"�zI�Y���㯭@v.R(�X��h-5ðX���c=���c+���Asd�V�F��y��S|bޫ/t@�ܦ��u�ó�aT����V�|���frkC-��!���}Šp0R���\@��
ߊO�3[5D9m�Zup ����\� �Uf�%�Or�+5)=kIH��tD3�d��ꐵ���⍕�S�{��r+q�*G3��_����ںY>�8��:��3N����\ⱘ	�t]"?�M���ʈ���LiA���A��+���JGF����;���-�C�>��l
D�r8.V-;2���;$����#1��K�)� 6�=���4v�e1q\��n��R�M��ri l7k��LT�+��d�9[�����,�qȽ��C����Sz��ݲ�8`��������j \��<`>�������v$wZU�d�7~o�g��9�G/��IT�	є�v�'p9L %s�s����7χ]� <H>�S�s
��n�z��Z��u
����?T)/l�Tݽ���:����ا#��K��0�����S����W����i��<�)F
��hi�뤧��������*E_��(�1��L)$�	�r�K38	}r"q���<�A!%*w�� j����Ω����O�A�߅��8F���d�(�m�N���f��p��ɕ�C<�/S�W��xR�7��ןf��- ��4y�|yG����N7v<%5sj`���نt��w;��V�򈳁�K,�p������7ҁ�Y��so]Kh���?p��<����]S�\X�D��J���=KI��?97{mĭI�86f��0�O���KQ��F��~�~Ⱦ�cުg8t�?�'�	��U�'Ed��n�}���X���/:��	�_K\$:��3�4���CE����}�)�������g���9Sf�W���
��|�_ٴ8��|U��~������y7��Y����O�bJh�+�v�<K1T�ޮe�16��x�$o3ګ��)�98�=�50�pU����`ݶ�ɦ걋)w,�Y�\H�c&.AL8�����`պ�ia\�g����/��SF�j�8���s�$
V�$�|��Tp������$����z�P#-��U�U�ʖ,y���3�.ĸ��u_ j\zAY���7Ȯr�MZ-��lSF+R��SJ+܁%��p��|����^����O��.�FZ�]�e6M@���.C�G�y'H���g�z�t���'�߶�&��|�ᤤ�ꎧ��{"L��^�z��=��+���Z��Ŀ�j���I�d&��WӐc?�Π��
|3ۀ��r��	mk�um�`v���}�|
�au��N����eљ�vgݝV�{e��B�}S2�.�ma�L����	Ks,��!r!R�=� �poU�lW)�]�˿�NA�e��0�����T�ԃA ��D���%��VibF��-1x(U+-b�����o���r��������� YhV���h
w�K�Ѡ�@��g�=zgu%�%��e�U߂Y������"��Q��h9*RрR8��3�G����k!�7%}ѣ]��q��hg�T��"�}��iԭc���^� T�k=�w4x��`���9 Xa$	g�c���9����ƚ+����� Ӟc�F00g�����Z�8�E��7���)\{?����9�"c>杖Q�%�'�ؘwh:��^�D-����ʏ	R�ʘ��ɢ�����8��^��(�s�l걄��
8H2k.�BT�0��~J�A��ru�S���N��s(��:Cgfg{{W�Z`��o��t��7mh �֥Td���P_�I���P��D� ��-D��oh�hE�s-�ʧ�%��ze��td���5�2k㕆����ɷ�#��Wp����M]�=�4?:��9q7�#�q���7�'��K�s�6r!ۗC!o�DFԨZ�<�0���Wdٟ1,�D�X��8
����[C��6E����ѓ0O�ϻ�Z���+ 9�_�����H_%ŝ�a�sr)M�h�.!��d�bn�h�X̾��CQJ�+��r�b��G�ģF	&f�T����@`8� ��Na���~.�N;�k�9+"��9���
Q�~�[�N'�^"-�k��r	0�.뎝���i�q�0�;eF�ȠrT�t�,�= ��^M�X�N+]�=H�N}-j���)tf�u0�j��qjS���3Q�Y��$�.�|@GP�5S������Ÿ�=�E|���Uѭ���zU)^˿ml�>ԙͺzqT���(i�^�A�r��m�ޒ��9���
�G���xﰌ������II���LI�9��ő�lCdL	)w���u�ʜ�^>�}�S��	�_��c��G �u̝�� ��=��78B�f���x�|� &�P��<�H|� h�F�,w�7�Z��(��¦��(���C�JԳ�^���5�k���C�&Nr��Y7���|�@!<L����R�a�zr�R��p{_���
�Gx|�:;��ޮ�>L��fS�.���"M� �0&I���������u���J|�
��I�-;s��Y�M����0%���Za������N��b]���D�o�����evĺ�w����l"ؗ�a�x��T@��0���9��NK�yTS��O&��3��*R7�I�w���^f��b��B��E��u�F���8���m[z���o�)62@�MŌ�cv��f�Э^\)Fӕw��������?[trO ���\W'�'���
Zn* L/$�`�Z��M���8X���-��,�)����[(�M8�.a���Y8n��1���H �M�E#Q���ޥ��i�+�w���;��6�M�LoyT��G�~2׊�����2�Q�~b��l��C/��;�->��E�^6�NA;֞�6���쪬t�$0��*�E�Z� �\�a4��׈���o�"�eҴ�ߪ�H ��$��dI;�^������
p`�SƏ �^�u
�jK��(�Ļ��m)s����ԧ�-�	>�H��ЧX�3qXq��qA��ɯ�X��]�M��Oytḱ�!ҩ�oCԊ�T�A�V��]��iߘF� 8#Y��N[�~��̭NN�o�1��S�[�hYD��0�,�-Ѿ<���1\���ܔkA/?���.�雉������.��I	�Ax�VK(;ƥ}6��;R��a�6R�F�������K��o�i�ln�� h�6��8g>���T��Xu�����uױ {
�t�eF����WI�k�wضpZ̩PC��m5�g1��������k§�S��?W�Ӎ���L4���0iG'��j�y
�jz������P���6�2��%?1�2�:��ke��x/[�p�2<�C���T?�K`h8�n��~�����{H�H�_�d�������
����w�"S,�,d���:E�j��BEm1������ac�����Gی�� c���/�_���٢���3�*(�k�+(%��DkKj/�q~3h�b�@��$��AKYA!���q5
%�i�	�G������/�3"��/���nz�R;PF�a��<.���wڦ��~L��)� ��E�iy���\L�����[�zX�6�kP��v��9���n�z��ά��,��թ��	�o٘��7�./h�}{8�m
�۾Y�Z�]Х*����p	|�U��"]Mk�s�c��
5U2'�=|�a�5����4p)1싖�}�J�T^߉�R�
R���}�3|t��oi�Ȝ�%r�[�$Y+�5�/E��AR�BQ�|���W��W{,�]�{0����m��%���a|���DEYB�?6�~y�4������W�rI|u\�!�X�D8V� �`k�XL���6�nB��颤��-�\��/�����`�b����R7�u��U`�qѾ70
�f�������_�5POs���XX�����N����Ι�௤��� ��U�Ͳ�E��B&�ْVGN뮜4V�	b)躪�������㻷�[�'::"��x��S�����c�gM���=Y�mK���]		}��T�av�+q7�tb��?`��v�5�X��
��(��Ԭ�]�����RtQ	v�M��d�"�c߂��cH_|����*�!���`4&ϐ
���&��|F%v���~�.1�o�r@Qj�%��J�4�<E�M�6��Q2��7M�7m���Y�h�>����=����yuL���2b�SH�M_���ރZ'*����� ��DvrI�̘����gG���ϧ͗%��W����顧2����ѱ,E ؖ&�1Sm���RC�(~ItCtf2�_wJ��}{�
b�ۨ���:��u��	c��K�?j��1�^G�	�p�V�b�VЪO��#c��������rbF����MS��Ny���y+������RP�PP�eX��>G�Q_R�M�M��w��N�
I��>��[ b+3�U%&�a���(�����k���Gu��ܯ J���A�<�M�L6+0�>8��K���C^����Wicn$��)Jo�C��E����O��֙�gZed�CE�ɹ�%y3:0J�oʕP���gS�',�!>��DE������gg\�|ڏPh�	ķT1r��l��*��L_,��	��~Ȇ��8�ҵ�i�R K��w3�j?��FE�^k�cԑ@i��ά�(<b��"5G�@|i�_�����b�����פSVG��q�tB�9��5(�%> J�a�׆ƨw�qy\!ǈZs�t�?� �q8�~�/��&5F�@{�t��)}O�O���j4,��C��˒�d5����@|�J2ĺ ��7DH�`gt�Sqt��ф�9Ou;�COdpqtc5@\�Tx�q���Ζd�B�3������[����n��\�i�>'�RS���847���h�}p����7�$.t�̉�0��(��^�t��ee)���>�L,s
�� �<Ԛ]M�+��
���S�@O�5L���T<�J?�#�#�g��]�Z'b�A+|b� c�c�!��T��*��7�7ꮿ��k"��-5ᾣ�.��J�#���)�)iݐ��U.>kZBŉ0�^
�	�r�W9���j0\2�zEL��(���ӺI� Q��/(s%m�ml��]tr�bNQ~�|F�����Ö�͈�pM`+�ב���/P6ˁ��w���1po������*�N�Q�?��j#����}=��w��>r1i/R����[jD�K�XL��@|���A������a�c��aB���D_�I�*��0hTѬȝ��3�izA�W(r�[�2L�_�B?�DyO��p,#��:����$��XAJI�lh��/��ut���hRWPѪ�����6��ᮤl�9x�ӫص�أN8��`xc��Z5��������aC2C�܏B�ˉ'��l{��<Ӊ�<�_�{��ʿ�L��(��}�T��@�*���i�j� q_��@Q;/J6��g�j�2��V:�U�����lc���ѲN=b��ԉ�#'��'Q�b��i��4�k��D(ɦr�qq�u����{�G�#`�.�O1���C�ϑ�����"�Ү��B��3#�8��҃v�&c%$��#9%d� #]=s��2��v��^pdX�
B�E�,�1k��ʰ�XǪ�jg�`����@O�������F\aJ9�
+1���PU��W����R���0>���T/H9�!�+t���=6:�ch�X�ܯ�X�·���0g��A+�<��W7��uVxT���azn���U��̪�J�\?x�&�c�Ä�[_'��߫� ����cB�:ͳ��?���p돥Ez��*��9����Lc��]������8x��M<Zs���J��Έ����J(� ���*|�6�\�Y�P����&m���Ȥ��c�0�.���M���T���[�����͔�?��Z��}���e�S���&�H�ø��Q/4^6��n1d�o��[�O�:�2��wRh"M���~�j�������ZZ�iѫ�s���EH�L.ς'��b� Gf��[��Tm�TШ�Z,��%�m�:Z>O��C�)�V+U_��?
kix��%D6f��W��	R#�3rЅEX�EżqQݽTfp�7�M���L�0�:��3%�k��=�y�<5�1Z��9Og$7�d(�c5�(<h����5��S�}���t�Js�>���~��m��E��O�s�����jl�G�B.N�]O!����p�&��
����'4)�T��z�)�������G�'r�����g����"�	Mw~��쟆7�3��Ӣ�n��vr`�5r
�wp�8"W�=��^��'�mg,0��j�w��Z<O��Ç�E0���r-ʦ�
:X�W{B�0f��	t�?`�Z�?N	��L�J�~����7WM��J!���$)j��� �!�6I�szo{�c�1�GX�����BC��c�V�Wb�lW @i@M:p�F�	X�:=��Ig�Ӗ=T}AT.�����"K5v�
S�[(�2x�kp��W���:��	�����:JM<��&�}�^s������-:�J�7�G��3��1v���3κ�5$ �ɚ#p6w2ڹ5�)Jƥb=�m��~|�
�|FN��윐�͋��d��:q���O"a�+֬"�K<]:�Oa�?��|h��O��	ѷ�ԡ6q� ��%��L:N)ܓl-_C�z�N�������	P��B�=�աw,puU��2�Z�b����U���@8I�K#����~G/,�{�(�(�w/�"/�p��'�F�7l��MJ6|�6�g���N0��W����f�#�W8�<aׅ^�7�$�S�Z|�����n�������!�~�'�jE�L�}���3Fh$2����%�O {�8U#~�Ku��A����˻��?	Q�:p����}_N7[���9�uQ��!\���'����.x��,[Pkw��������TAe�����zС3�|�!d� ��
g���������ӹl �z�ބ3)�V��j����O�S檼�>���%_ߘب6�j�8��7�8�>Ȣ#׹���ϗ�k���ny��H��;�)1�8���N!
��T��č��k�w��Q��]�xh�x~��
����M����?~��G:�二����F�Z,P'�p9¾6	��u������`�xG�T��`:����'G�c�������x�*5��+�������k��3��{ 
Ԫ%�+޸����	�!t��ֺc��8g^XF,�%HOD�g�}i����3�˚��(iJ��M�?Zܟ�J�I	4�,���F��l�����(���2[��3��?��ȸ�5~B�Ф�<�
(��i#*��o<���xBj�{��=]�c`�������;$� EÑJt��Ǘ��V%�K���v���N�t?i*��Y�� -��2Ѧ��K5{Z4�JǺ�쿦����Y�������=ٹ�Dh�T���-���g�Jc*�X�V�@����K�foB�q�'�.Ӈ�G��Az;d95��,�uΎ��)� ���t�㇠=�"x޵$�3|�[U�'�Ն��k������c+��L���p����t�c�T-H�K�����\�"�/G��.l:�8��K�vHL��-ޤҫ�Fi�,)�*��[7J�W�IDX���w��OJ�����=�I���$u��W�AX>8������݃wl�A�f�!���?��n"��jW}=�'�#�E���W����H�wN���y�V��`��3��(
��jh_7]�.�cE�E	���+��9�D>�$��W g6�9�����+�,�+��ۆ���P�!�P��o�8�''�-���!{5'@�ݜ�ډ5����2@��uj�_Y��r<�<#| �s  {,?��J��"��*����U�R�W�rEc�L�y�ѐ^\�-8�R�um߁���p'�Q��V���0|,�_=�����5�$�O���W�ͼ�����Ik\Ŀ}A-�61��|�֞�����*��:隈�ǀ�YE��s|���{�3�r>�nQ�K9��
?>��(� p�����#��]���;��f�w���"Z2�|n��4�H�A2�U�eO~���ۀD1@���I_�༳On}��F='�JB���?_�@�=�+T>�bv.7Σ���\G�&��DN�A���9���H	��e�.�>�gca�� �N�r'�X7�Y�,���8�En f�"�����S �
Ў�������ݲ��sQ	tG���u�ފ�H�9"����.���h�a}V�@@���q�g
�4�����C�����@1�B�	=��/��#���R���f�U(�����P�E�V H�W�	�ס��3L�T���Ӌ���2�p�J��N+��V�-UZ ����و�����ӾJ:�J���=���o�fU4Ն���̺��j�vMؖ*�����w5I��UXl�Lv�j>���\	H'+ch ����Z�B]��y$uA�˶�\,G��x[=�.���]@�*i��L���T�uy���W�ۥsZŪ����s}'�A�		��s	4<��T5 ��ڵ
1��_�<r�	�L���]��5˰<�������BЊS�*������
�*V���~.�`����]���9���˧��_��nꃽM����m�#�OHO}OnT�;C.�A�>y�c�z�"J�^aa�$Jn��M+��s�M�P��	�`�r�?�7.f�ϻR�)��U]�%��:�p�#�1�50�����7��'~�?�\i�T�g�r��������m�i��NLȅ��-�Uq���
?�[g�!����"1��'��&V�B8E`I>Z0�c���u�>�؈���;����R�e(�-�O��W3�M�$%{��Z|��z,��P@V;&�y�U��,��Y9zX�-�ò��.}:w�������;�K7��Ъ=@R��JC&>'j��e���!�1����W h�>��QA�����(�"����2o�[v�U�i�&G!I/.HFt�}��ᗷ��m�+a��Ri��pNza��J�R������,c+�����a��]t��2��e��0^LF����AtLG���!���n���PA�+� �b�,���#���,�w��S�4H\����S�s`��߂=bF=G�f��9g�J�d������7 �c�C4�s�4�ȳL�ӈMڨ,l��茾�g��'g<j�iȍ�r�41M�NotҼA��Gqd���	��
�υ\ֵ@KZ.����6�����F� U)�����%�k�I�Ρ�;S���w���p��j�Y�.�����J ��}��'^[��X(�a�I��z3�B?B�u�h�hU!���mgg�]���N;��}⛣��4�h�ѥ$G�I��J������>3�d��Ei|�t����,��!�Z�q^�h��zS`����k� �Vr�F��f4����/n2_ ���(SMH�b�Z9'�j��N��om�?4?P�79�w	!�^��V�;p�f���e�.|@��ʒ���l�_�E,����&8M���}w�����u�w�R��TJN�!�Z���{h�0G#�]���#uZ71�7��2C�����@ ��u����o�6��ІP9e���MD~زW��[{F7��+���~��������_u@��.�Dpawμ�p�[;#r�m5��9I�z��%�^ۋt0A���˶�w!L�*94g33��K����~`,p�@�l{#���n�`%o�!T{�\���Z��5��<�3�����1�Aho�ڦ�Z��}�Q�t>�Ý�m����O��5�"'�}B����,ک��`;${�t W�CAEJ{X���6&�p&4�����Ij��L��M]WJx����ܐ��Q]�T�h�v9�XI]�̂eJ��T�&���6��S��3ee��98r2,]�-�.
}�I�zꚰI�Bb_z";y{�e�Z�yX���;�}�G���X�K ����FP�w����T
����I�$�/�(j�0��Ϝ�@�3"�U�u�Y;W�#n�ż$d�����}c��s�f�]x�ф�E������V/����^j��'�ο��Ѩi�Α�|�">��Y�$_���� �v����a����K��*��-r<���p���'`VxX:��D8f�T�/��W[]���I�[٬!ҝ~����h��v�wJ�x�>��wEM�Y���eO���D��F@���	>/���6CBGr��6����!е9���fѱۺŋ�L:#QM����lT��; >��X���0ujN�����	b�9�M�����˧_l�|�. �#����k>TL���b��\̠��z�`���z^���J<MN3}���D?o7� =�jc��N�yt����MCo)��b��&?/tF�?y)Lk�NP���^��r���z��x �4�V��"g�e��GNS����$Q�y�.u�?�`BK�I�d�"�� <�dR�Oo���\ފn4�0��#�t1���?Un��3��+��ƅB(_0&�o��{�`W�t�FR����_ ��QZmB�9��Lt����@*a��u"#�Š��$Kq˭#���Z��W���z�^8#��s��)���&� ���ظI��Hs�޴�������d�{I <��Ǟ#p�&*��;�4	t|؅��s��ʐ�}���_ϗ���$�5����y%�1ѯVwZ�o|��BhZ���~�k�Y�נCr��]+4�\�t���-�z�#T!�"�ܠ:S�N�\�H��B,����.���P�?4]���1��Ob�ʺ���<d�{�������9b��K/�B��pW�y]�k}ɿ��j}�2��G;��we]�~��p\͇r�FoN�ۀ����,����P:�.��W�[��U`�)�v�a׳�w������Yܠm���IN���xYz�Ʉ�dUF#R�bC�0�ر�qQ��O\H��A��.�)���	�9��;�O�	m(Z�J,XA����2r`ta��m|�iN~�&��՚��]'��tBڛi��/����B�6��b����V}s�G9X�tb�Y��Ǝ]�� �U����Q���17CgȪ����j���`�� ��=�mѧ�gi�3g'�`����Lǵ�S����*C�F�Y+��5��
:��
����
+��[9�Bm����=��U��U�ڔ�s�0�K��WXw��%��M&Azֺ�����L�&lo�!q���#ѽ�W6�(��*	����YTS.y��j���6�e��wm��� �B~LS�� i����x�����x��!I4K�~7,I�x �g��5�&^uĭ�V�t֟/�ִ��!�>>�B8<Q�������ZP�P)���"q�?��x��5R�0+(+֯�/ҩ�b�5�]�b�,�bL|�M�A(��rx��bl�������*~�>��)��[˦]�t���ٜ�i��-��)�6 �U,y�c�t��w�->V��x�I�&��6Ôe��b�F7�10>9����5\��+�+h�d���3�׌��HEHk���3.:�1f�,��Y�I{
�y��=��9�$���]�E���X݋�2^���`�e���؂�~�K�b!���k���Q0��L�{5Ľ� m�Իv'�OJ�gU���>KE��Db��
��� e0�X��gPdf�*; �l'w9��i�C�Ç2�u���L\�ZA���!C'����e~���i�R�{�z��݄���/ki�����S��~> `��q�ME�ː�1 5�8��Vbx�JI.���Le�\����:�����8}3�־:��J�m�Zl4J[*�����0:�x�]�&�x�n�K�*�!�s%ZH�ɨ�ridm�
Gg��=g�*��0���pB�$�:�`����p�1Tfz�T�mE5�2��q����/�vJ�)%d����3e�#e�\1wM����B��Wv�H�4T�Bh�(����II��!cG&�9y:atA�C:��w�6~a0���\���,�T�ơG==0������l
ciS2�~ǌ1�^�Lb�K��؍��g0#�E�T����Va��{霒���g��P�+��S6��{o�������>���̧��q	>K`��bsv)�fV��(��4�f��DQ����~(��)zp�v�����Ȥ-sG���ο��r�Jç�
�}F�~:��� ���~ON֑n8�
�M�'E������P$��J�2�)O��%*��u��$nJơM�j��+ʽ�%�k�N}H����
�!���=s��}��J�i�	'�u�;'a�2ܱy5$����cK��h�鼃ʵ�KR����;�#���e� ��q��ֽC,w�ɢ$�϶8������C��\i2Qf�\�rD���}s6I����4B1��p' ���co$����`��|��TIt����O���(��
ٙP?
I\��]~�����;|�62-	t�z	h��R(���4���7����ܐ������j�j`�]�7�H�����1�s-�����g�j��-���)Qѭ�.:��		�|B)�<R_y�O/����g��J�S��"�������]�m�8n�HB�t:�A��Y�O���ؑ�4�#��N ;�y���T���U;����X�
���&B��F�.��ҹ=�}��R�=@���Y���GjSA�Sƪmv�:8SD�B�8= ݦ�iE
���������RT��� ��~Ѵ14�a:���vV#�C&�S��Faon�4�Z�bvo�o�,��J��+�8��.���O��2ӯ���){�\$l�PO�s"�-�	��%?}����p��A��D��1�((h�jA�����55�����rGbJ#�Zn?(��ʛo�.���$i�e��y���@�T����W����!y�&�.@�������,aZkR��d�1GH�>�0��}�]�I�QÁ4��/"���ȟ@-��R`�s�̴l�Tn�g�j\�צC�@����F�U~�c>���pO!���oV*�Zjv�ӗ��5=$�x���	����=?\�0CnM�d@6cZ+�wR[cUr�E5���ۇ�2�u��J[Bx;��F9O�H �"����
��J#�,���JqȲ%h�|c��$,�Fj��q��?�HKŅ�>�,�_�*ʳ��.��t��?Y�ӭ&Bo�y��f^�1DY-��1�N�'�E|�}PЁ��T@+�v�^��m�<�;���sz~�5��IY�c��\��T�H��_?M"�s ���k�,��<7����a+�����z�G���V��P���7��W9�yi�bUɛ��8�ò��-w�l�����8��%���P�UG��j��R�D��W�,z]��Ӆ���߂�����d�Zw�}n�rS9t[��Hzk����K0��}��7��n�;���&rtQ�ms�6�E���9t�s�KyϯÊ�1[���c��`c}�{s�.ѵQ܂�}��"����|\�0��̆�C4�ͤ0	$�t�GEз;"���s��E�3j��$v�.-�p�.�����F%�6��4��(A���g'3���r�����HpL^��I\8$M.̶�Ee�HϕHPRp�������g�_3nXX���o0�F3��i)��H��[RA�V�"R㶊V��p8�m���Q>�iG�>9p�"�!�j��|ի�s����ˣ�ZO���m܀�C�� \�NTWeV��5`�B����+�����W���0>9�Y��J��͜e��㎠����T��$�,%�ћ��u��Zi��]�=�J�M��8���~˥�?!S%/���8��(M�"W��K�ɺy�N�R�&�y.5�?�<�2�{d���n>v���8�-�HZ�^�gu��do���Z�ِЮw��z�
�G��ͥ�\VC},�M�U�e%���6 �|ͩ�C[��tP�'��ɫ�&t{X��E���e%�;��i_t�f�o�P��+�r,,p�b�� )B�_�9��,�pF�ko�m���o�=:��'�(fLK{Fq<`�EXtYRZ��C�S���Mz_�el� �y��=�WU�_�����6��g��E��p���F��02�]0�d�i4����|�HE�Z�J�t Vԓ��Ii�ـA$t�*r���Xxi�p4�NA�W�^z�������<�?�_W�\����(sx,_S��/����4X7 �a#@�`�cZ}4��`������En/��ǐ�d�R�#��\�M{�W����2[�����!|p�Ӕ8�����ղ@��o+!Tf^6��8
�
���6���	:L/ڰ�E7�>�D}��Y=��ܲ�nt�y�����\����NPV�|F�=�7�p��)q����Й�y�ڃY����ZK��ҁ֘�v��H�A�W._K�m��M��{��.�.&|�����h�� h��
:ɥ��I��n�) x�AI�V��?�>W��Q�B3�9T���s�a*:�A����b�'��|�'��� 2+e�^�~֛�t���<�2ev��/O�x�,��P�T\T��]*���9S �1�cn�$�r����I�1��~��r�yy���l����w�`��mܥ�/�5�7�k�DW�]*g�E/�v�0@�B�a��9
��f�*f�@�ˢ'�E�9��3i8���Ǹ�F�SՕ�\� {��`B���N�|�a2�����/L�`.��$&��0k�_���WwVw
���\��z�jܟ���=��M��T��-G a)ۉ.Y����N�������UC����gT/���Z��L���I�c&��a�1�0=��Vd�C4j?�GdFD��)ٶY��G���53酸$jo^�0i��Q���܈r�ud����k�-:b�G�E�ˤd�����u�@���f����!���uFĢ�s_�ӓq��_�:���vt�\�f��V�&en�;!F�z.��e"5�K+@Uy�	�fy�&S�����dB,�8/L5��!�Uɀr�����'����q���g���;�-�i�Ó8�R0R��;"�]�u �hN�JU�i9\#��a(H�L�|�21b���\)	�K+v���#M!}���V�L��A�'���(�+�g}Ü'��.v��X�H�7��S�HW֩�O��V����ٝM����ӌ�5[_;
��hc�qN�����b=5j�]�e�E*2�L}b���	���x��q�ym?�����IU$�T�y�1b�Gw�ë� ޿i?bxP����ڂO	~F��t���
���6��znr&u�
����k��H�ҋ���A��'�7�4��ڛ���/���sI���S��h_��O�O�`L���&�AϺ�9���w`ÊT���m)Oxu����!{�$����j�:v�����CDx��c����
��x�uUN4�On��N�Դ�췃#�g�]�Z=��\[�Ĳ�r�X`Sf�y.THnh9����i'���E�<��0�&'����Vّ�^f��}���]�O�9w@��Sc(�M� ��v�\� ��E+�gj`s���B�Cp�7TϱPY�{���#Dpn�N��[�n��JTMWCPr�&lH֤a�6�Ĵ�D�:��ƞ`#�N6Q���^h30���_I��q���J��uI���O�}����9���TiZ�	?��2ޮ��0 � �!�pCi�H2=H��V	g��Wo��n�����0��Y�*CܝWt���h�Id�~@O�Y\�t��c��BhPP��l��O��U�����ٕ!�"��˟KR����\�s����m����m��}��&�_�>U �n�����w�����؁�.w�-�dvFa��:�*u���H[�
9�� J.}ۿtb���$D�D�J�~r���('s�壵�ꟍ�y��tXN/�+�a�GB@�)��{q~gX��ٖ=(�'�oS޷�<1"S���,(?ʐ�d�Y�ʙ�0����u*A`y�y�M�!�f�ӧ���ƺ�L׿�S�n����tL�&h]�\��K�W�
�J���yQ��7+ijk�	�ւ|��5ꊈ��IE�>_�R�h��m&p*eG�s�P`R�����Ù΄M���!˩�������1�K��Ή�K�H��H��5��I�7�hfsճ���.��V-�mO��a��G���2DX����?E CB�V3Dyu��m���R҂�[��G��?�/��֗�������˖\<5�~�r�H����ON��]����2�N���݄��	��g!vd��h`mUNz��8��Y��D��U��G���� k�G`O(��"�3�Cis��(�1syJ����d��[���o��|�Ze�f��k� ���^���bVz�Q�Y��֜�P�?�Ҋ��N��H�4���|j�䈸�:�d�`r�؞� -��A4V��� Y�T̔�SL ��'v|�s���!G����%�&`�[�KD��Bs�EH�c�^�To�rX����٫������E_U�����z�"?R�4�~���*�oX��5�Y�"<C��f+6X)�0�"��P�*�|ǒ�U��N�q�u�����ȲPޫL��d��;�^qp�|˹&��x�{S_-���jPW�[�P�oH���QOou>�*Q�]+d�A�4��6��A��FG�C��P�,���ꔉ�z��x�_!��ŴLXF�:���6���ty������Ęhw����Z#�B�1Fؖ�$����9�ؑ����U�����x�&��p��!�{w_
��5�|�{}"�	^��t��|j'a�Qv2��&�gIM	�ѻ���yAy�)Q�jMZn��D��- "���&6��q!�_׏��̥8�Ha��^�����^,Y#qp�*��X�z�ve厓@���Kr�5�7 l~��o̤�)vn�z\iK���+zb��F|Y w^��2�|~�¹��}���e�'K!V�Y��8�	����dy�������T/1-�o#���"�.��?8v��bF�h����[R`'&½�ӟ�-��3;�Քw �����f��*��D��qa�Z�"/�H��ә��ء各���2Z����H�k���r^6U���x��"�>�Vy$���<h���\��1�𫶎�1��%9�O �`�Nx#:�h7b���~@����a'é��@��19����zm�NSЮ��~���J8F�9�0m�IK5�FH��E�	�#f��
�9���ٮqMq�.I�����Re�ݹ��`�l���adz�º���WWϷ��h\0��f�Fz\�n����>!����L����K�(��w+��R��V6������^�h�Lw��'�i~D'�����reѭz��Af�Qv�9;�tR�E��������fX��Z��S̷ȍi�aN���S�W�?�^��4�,4~�4��wEtd�w�6��OWf5�Dr�q��Li! s���"��[A��.3��B���_��K�/�N\��Z�Y�ZK�~܇+"���q�6T�����,o��5��Z�}V,�`C�����$�a��i/wl>���18R�����?��m�E�:0J4���&��\&�EE���z�)z�#z�[O�^.���h�|ш�_�[�yJf)��]?@$!Â;CB��ǥ5�m:T��x�?��@8*>�2������O��\���C��,��(��/I�n��#>�I�q"],��GДWd�k���S��g�ĉ<
@猅ܐ�f�� 1�g}�I��y��>��tR��X�qF��@���dn�c��t.��^f�8ŊX�����t�/�]b�tw%���6�Ta�#�z��U�}bb�EVeq�j��A��kB��~��p����;��5xc���-^�i��G�.�܍��{p����E��+��E8�"z$l�H�2]]m��p*���m<�ӆL��+܁'�U-ʺ�l�Qk�^b�Lh�U��^��m�$��6���
��wM�x�xp��?��D93Ive�����5ods�b:՞��K��s�B�Rߓ��5ʇ n:x�+��ۮ�R�֏��Dk>����tʽ ������e�ȪD,*\��N�ʲ����7#ūL~YH�ܯ!m7Vu_� �$��.Y(�;*Fqer=m/��y;{�K�
Xw��/�ݺwk�'�7Q�����"��ﺤ#�r�F�
˝�C�P�\1|'l��m�!t"�����Q*mh��cZE��%_�k
���a�p�����V�h�Y��T��R������f�<�tryP���i���u���m�5��0z�"����(A��K�ӄ���-	#+�/78��y
k�ԬǷ��e�{m���6����q�o<�J0ǐ��HO�䧘��rG��c��^������K��K�Lb�������|�8R�Z�o�A��%^c�Yvuw��j a��4 ��Ye2�*��@]Q���;��x�-�:M���U (�6B+�c�)�YӒr�p�;&F;s���Հkk`��������j�Xr�J�e�L����a	0A�\��}�>ȿ��\�R{��2f�l���`O��ۜ�}�b�(��oA���4]��š�r���El�Q%���1����
Q	|s����U%�jK�Ul�`�GS6�9&#�[9��S���j�C�li.�A�������B��<�� zb�EQ�ٗŊ2ΰ�݄т�����U����B��.��c�WU�I"�~���SA!��� 1#�[�U9̳��M"��\�U�V�"s�U�����5�\���EW2R2K^�o�&��2.7�(��$=��#i�����*��c>@Yq�L��&��k�,^Μ���J�.�4Q@	C��ǰ� `Ѝ��UG3q��7�.dJ���@9�R4��.4:~!P�5���V��#���0�	���,u����M��sX��:+�C�:{J�bjA�  e�b�@���Ѓ6�s����ǚ����t-I�V���s_��O\ka��lA��r,��Uo�yz!"��X��.0�����jv���� �����'���2�
�^�^��F{�H�����<e*�[q��Hƥc�X����bq���:��u��[����j;�[��/g<?��
�OZX�E�BـF|U���i��MNo��pv7�3�"�>�|�x�DL��#�Z=^'��kc�k��I�Μ���Pb"�%�:���Gע=O�v*Z��E��ѥ�6rJ;ZC��^��(�
i�8^p�;�E�)̐>�,���_��4V�yB齵KT���J}�y���U��e(�(Up\�F$@ڻ���$jD�>
u{�w�n��^�zkś`�s3yv�b���)a�~���8��Z��bh{���6	��C��c�V)H��1	�f"`����~^J?��~�GA�����nT�S�q/~�y�{�@c�v���]���Z�W�t�����Xy�z�\�T��6q�Ȳ�~�сw�F��	b��龔�?��(�oy�^�װTzݰj�
Tc6�P�~�w���� gb �w��[~��O~�~���� w�	8����{p0[���ق5>�������`�46�ͭ��5̷�� `9h�.���ۙ$��{ �jZ~��¾K�����OLeܬ������W�i���}��w���+��]�_��Dss�A�,��^@Xx\�|\�o$BmC�@4������{�τv<!���2�w�L��~6���Zd�^Z_����[������gϫ��п@X��`���PT��=�6L�om_OS8��l�WMb[҇�2�������H���h��$�Xx슾��c
 Ohi���+��Y%��o�e�^>B�D|6�2m�� ��Y1�H[*t�j�zѥ�=0�v���(?Fc��Ԧ��g�Ʃ����[J��#�y�~I# q�TVum�J;\3tCf��*�%\L�s�F���NE�7�m�0������@��db�[��~�g��m�e�Ʃ�R �vn��J5'Z�YA~��,'!#z:�)ƞ��Y��~��y)�r��(��q�}8�,�ձ�OI�yqz���9<�ᗀ���%�<q�K��a��$����g~�	?'M�&�(���$���.��^�Ǫ���AJ�(x>v��0=\�O������	Ed�>K�6\��u?(X���׈.�=�,?����n} R�h�3�<����D��� �M�͔�^"s���O�p�~4����&JS�h�x�~*�?hmb�M�Y�ݧ�I0=�ˑO��{�o���*o\s����-Nxq՚���LL#	�O���Br� �3�z�*|�ɒU1WeQ��SSG���!��`p��}P���p�2�V����"��$�)�9B�E��E���z�5IM���n��VݑN��G�y3�Pz��|_�����Q�K�j�eRq?)єí�V�E��<��u�⅏{��d	�O`{�0���J��Z5�	|��J�T��ǔ�Go���(�V*,�����h.���}��:��K]�Ki�v[���s���a��x|<Ȳ�X�^Q�({6.7�����rS�m jdȖR���X,��]����������8�ey'VP)Q�V��L�;��<�o~���U���y���LX�E����a ��r�0aa =��p�we���a�-��g��P���d\��:T�f]e��{���]�塓�Y�ڳ��Z:��e��)y.�F��!� u�.ĿQ'x4�VO�N��@�����h�G>�h#�$�Y���$u�Ƽ��[��3��p�۸[��L��7�rߴ�M!͡�)۟Qv��	���4�«�I$���Qe�T\�@��`����&���	%鼪��D��f����u�� �b�j�
6���
PU�?�v�JT|����ö���5:��E]��0#������.:pk�k�l:c����g�*f\a��A�s�c�;�~Js�O�_��s�	�����;�� Ed�J⫝̸u����?�N���ek���=lµH^�~&f*&?�e�6�ԡ���Q6�3:A����@�Mژy��J�-eP���w��=O��$5�۲�42�������@+�b�ٴy5�Ӊ5��@QSv���^����֤M*��kMn��[QCJR�~���|�]�������6-u�&;���Ӣ܊6�V��p4���,/������8�+Q�Wă �mo4'����i�Ok�W$�7��-yb�����0�t���d��|���x�E��I'�)~4�����gd&�m���u��i�kR�������hE�(m�r.�9���6:�q����p����.18���%ˆ�/�?������(+��k���wMʂZ9�W�ʤ9Zdd��i7d��f
!U���)A��w��1�⭰���#BO�J���m��
x�|�U��h��\3�9�Kudּ�QA[���<ԈQ��+W�]���#�`�J;!e�#B���=�qH����Jے������+�8��������8���׍�HH1���	 ������L@�}����ȍ�)i>�R_�_���J]�9�54�V[�D��!{��=����+90SjY�㙜eAD�E_?6�_�:����*)�2���e���A_�ʻ�U�F��ҹ0�o��V'�k/���Q̞���?T��+$;�},��4�j�ٻv����Vz��J>>N[�d��[��&[a��qS��"�fd�eRzb�\��ƚ/O�Z?-BH.��qq\��N)I�<���+de�p*���}�Ivɼ0<��v:��x՞!�kb���:����v�cV
$a�� �< ��-�zr|�X�։F����sX�ԿuŊț�w�ٮ���#��N\� �7g�^�� tE �!�8�v�m�L������ ����Ȗ�\$3W���'����E>w�Y<�b��*��u�����\st��=�>A?�+������U��a�=t�����,���K�`����	;H�6�=��|�x9Mф��c�n/������r̚�[���AQf�IҴ�B�
���<w��!�tݝ�6�@�lH���2!Z�ļ�3ZT]r�MSqg|�A�&�5�<��[#Ï�C �5%/
��{"#Ul�o^UA_XJk�-7gZ_�e����	N�a������ϡ���ۜ5��+oIu۔�V9���T� ǭ暈�It�O��?�"Y�9r�)�j�L�k���gc���R��:�0p����q���������R���聓��@VFh�|?dtj��KHH�.��)=,Y��{�1�U�/w�Q�zRڌ���e8To�n=�/sn�~��s�)�`/վ�4��>a��yp�J��q�Q.�Y��=׼H�TK]�$���3ƅS��U������ĭv�{_�aQ��I΀��Q��$���%U��v��&�����񟦞�y�ϲScX`0sM�]�Mq~�Վ쿺��_%>�C���������ѩT�t ��]U���S�j��SV<%_�{��n� ���k@¥z�=ͳ�Hu��c=+%�y�p-s���I*ڪ��sx���,�v�!9>{a�><���.�W[��Bp8�`O��ǹ-�ℶ��G��P#{.�F@m���y�"	�!p	����}\Sݓy�yh�k�����B���,��Q̎qЧ�FN����0I�)��1^l�j�Ս�Kf@%F�wx���S����D*3X
5��6�M���Ϭ�]���(G\g�#�mO���vJ{�Ƶ�|�/oU)]�m=��V�4���_�M���s��ِ3Ta�M���2+��u1��ď��}׊�T���%��.̊�|41X��a5e,jw�{���t�K:6z.�|��  ":j�2��0��3���u�kď-�`a~1�}L�M#w�zȪ�}O��v�D8h���η�~���m-M;\�&qi��Ʈk�^Ӫ�:ъY}�?��C�+��W��D�f9P�I���4��3�[dQ��1b��u���5m��>�P.��i;���[O����+�'5Wue��rQ����Ń����:cM�� ���g��!|��I�����0|�w�����ͼW����f�3�.�j���<�~M��u��i�8`��q��٤�C��=���3u�U?{�k7�Tv���e��Jq�jΡ��ڎ��#/U۾H��b�<����?�$,�I��j4�Mɩ?�"b_��8.���p�^�Q�ߙ볉_A���>�te�ʐ�Uea���6����u��=����L0H�ͮÒ0��,����鞘��j�<.��=�Q8N��(�@6D��Q�Vq�^�%���u��5�w���Ĩ���i1���`x׸!q���y����Y*�<<<%��K�Ԓ��*0g�aG�3/��p�� i��#bOq�v��K��yK���.�(L��wN���7�Q����PΕ�_��p�_?lP�9�~�s�[�ѨՊγ�ۢ+5[�X��L��'�o\�f�X)S
�����$�az���q�C���ɧ�4Q�Ė��rm�+��5ߐ�=Y�Ta���-č;��u#�Dn���Sw�
! ?oPP�y0��@n��u+���̈́ &��Z)m�nEʉo�?�u�VJ��o�!��̻v�C̯�G��dKޚ���g�Ġ�@�B؅��A��*�]��6�A��W1_6�d)�J>�e�?��c~�9\�_L+t��L�tєk[�ʎY����о���4��g�('�%r�'6"[�f�F"� �RX5[t�?�I���n�B
��/?>�1�3}W�F?DM�&���8HT��:ֳ"1�"]�h9̯XAw��;9DR]ZO��r}�����E�a�|a� %M�F��
��"�� [� �Vh���>Z���m�j���<)q��h�$�T{�T-��}�j�qDԀ5���E�W����I��Y�l�x4H|2i5 l�t�2W}mҀb�
�"����^��,����.���d��I�������|&Eh$�Mr�$_za�m�{��ԝy
�-�bܺ��D��-w�|oI٢(�-!5E��Ag|pP<���ߤh+x�q��r1$t~B��3�%Ͽ=}��^�Y�п���6�=�i[N�N�t"^��J��*���d�}=n%��`�)>�ܿ8/ 2zAc�B#�G�;jw��y��1����f�;B)В�yd,�s{ fGsI	� �N:�>;� ߴPE�I�	WWk�����U�q ��VqwA(A�k�|���6��|k��]�Og���Ӂ�I�_,ҙUTt`̀P2z>�@s�)R r�SCA�ߔe�l���Le񤍵{A����#�����{�ܵc����pk��I�s�ruv�-�%c�[��L�B�������2Dl���+�N�g�zbM���Ǟ�|��%�H��T��F��޷�u/�>���4N��Qf�rW��^+Y�j紭v�S�����9�� V�=��r��[!6?��c,��A5��p!�Gߔ�c�+�h<����x�u�G�{�<��Er����w�Jߦ/����Ĵ4B���$_v\9[���N�oy�k/b~���YpS�Ǻ�`J��.�[�3�\��FkH�����w�1���|0�Q �V�$�0̸-������P߀1�]/�hқ4E�x_h�h|� �/���r�����������Uw��K.�co�r�F<|1xـ��hz������<�ؙm~�4����K}��[��]*�9���q�؁�PS��[D���#$p�;�{�)�V��R�����K�$�q~����_���U��TR֚_&���?�>�LkT?��w�v�B"�����k�����Ȝ�} 7B���:�RZ�x;(B����F3R�Ϡ��YJ�\!�E�K�;�j$�n�+t-s[�#|�]%T�}=��)�	�CE���!l�۠����Eo�����r.�0z�쒰)�v5<F����.�DD�*%	�гYB��T�-qͱB��0�%��d�5�B���Ȭ9f�/������ ���E�ԒQ����	b'P"SbtM�AE6(�9��B�T+��p�S��A9ٵ׏��SH�2l�j*[��b�j���;j��з���u^�|B��2%�؞�*�0��9G�[�+��ʀn�Y ��C�jS����){�w��`��a�����xe�se�~�e鍠�1@��\�V�vƶz^,=)�d`ѷ�v�#���۴�H9l{c�"�x��'�cC��F7�Nm	�ꓱ�wp�;�К�a��RI�V����=pC0l�.�Mil�������Z�Ƈ
��ŶF����)-"Q��Vk��e(*�S٩�k����!OV�xd����2b'�pa����ϗ$��)�ʮP;�3}b0ȋlŅf���~��F:�4�3���:��K�i���X.Cz�!�c�Y�S����̛��P�1�9@�J�wM���Qe~2��4��\M��5AX �8^�~�kX�WB��1��w�籊��W��H+����*Na�������4�1!�/V��-{�?���!���)h��7�d����Pk[����|�00��R2�L��V�?��;�a�>�S���H�]c�1Lq�� JW	 �aL��l�a f\F�@�%�Ǌ����S$��8(�I�#c=Tml� �hSG-7��~Q8�]44�f��"����m x�8���;�w/�dl�լ�ooDl�{ipYܴs��j^:�H�	��i�G��t7)���	u~Q�P}#�_�Gn@��?���ʀ8�o�D �`�C���>��/�"l��Cэ�����<�E��Ã���ܣ�x�3�?yo�����s;9� �c��z����=p¤���%;w[���"P���q#̴�p�� ES�o����@� ��#)�d6Y���Ҥ���E�`ֈK�#�F��j�̮w�6������,������@�\[�����m+ER��=p�1�FVȎ����244F������ɤʖI�Z�����w3|O�Z�mX��Ӗ��+���CΣ����<b����s_0�ڞ<(�L!�I���7Qއ�8�f��ڡ�WA�.M0�z�KT�n9�r܅�,;8h�����������i���ј��L�C���}���n���ϊ���� z^"�r8"���:�[�}�/�C��q����3I�����2�P^P3���-/���8�?%?��{��=�<�+Uo�MSz�R���*R�/�r�Y�MN�?m�0<f���X]6S�8٨��dvM��|���P��ݗ�ar��n�a�XTA%��|�����:!b+�ӏ�a{�&`��iW��ѱ��ИBn�Z����;$��oc%���Y]8��'wO�WhWն�Q�Z����W�*%#`m��4�\�֝i�f����Ѭ���W�����w���i~M>�����3%�NF��)�v���m}�A�<�["m�]������z��8�ie��e	��:�H+�D����w��̬Z*�T�y�4*��qA	����v�ށ��5����̗��S"�{-�d7���v��m�?R����#��h�ZPgp�.�]���1"��cךL� ���۶Đ��W���� �g�|���߹܊�yi�4�f���Pt_��F$Z��gd]�@��@h#+Y�NniB�Hs�(�/x]�K����J)�gIAwؑ.�����X���D?n!��5߶����fa�v`	�oF$ϸy�t�ǝ�D�0ߡ��C�ҝkM᝞{TԐ��Q~9*���T��&s�i�9����354�x ���F�Ѡ�nZ�)U:Hվ�g .��Be�S́����F��N�)��g�6�f{l�n�w����J�t�f�?�3<>XO/|�5���D�Isb�o�ua|3hJ3�����Ɗ�wBK��@��B';����KYE���p�Q�����ܬ�m@`#�.R 3�Fz��%���ͮ��E�3Sٷ6Ky���m��-��?�[n��8mƟ
��ʗ>�߱Y�N���y1M��$���g����m����quk�,�\���/(z�Y�x?�����?�v)u���������Cz�E �.� �5��M P�vZaw�*X�O�E��=5���I�+`�?�%��#�Z��9!��)X�ҋ��?qg�w�,ʖ�1���BC�!�[��b4�����@5DkR��DT�M�`�/���x�Uȳ����r-�0��DIǄ �4�����eӹ���ʘltrn�Y��m��WTW0�������(Ai�(�����4�m>���S'cG�Kil�I��樤�^�:ː~�Q�Y�~�b9}-�@�nV8�H��J0��b�;�d!�[��m��
��P�k;��Z6�M�p�X�4a��tWQ����{Q���-��-�WQr��x�p�j��g>C�iT�`	�);R��:)o��B�y�[��Z^
O:�Ow��%���:�*G_���a!\NDs�N�>�آh�*)O�b���a�Z����`�Ɩ���B�H��}�P�N>ޫ��U�4�F�q�фp/t�9�ح1z���R��a�[�����mzg�^���G�^�	�g�	��Gz�9@��BD$�Mb8�27��=�=r�(w����E��W����%��|��?3�oG�~5l�=���4��S]���A�n���b��~i̢,��罸rDy�vH�*9�#�#��N�š7��QH�Q��1Ah�6n�2�CT(�!Q�+0���L��E��Zz~?{�B.�5>Yހ�?��7٬�)��*���z�e���K��~�=�L������\�a5�Z/%��dנ^*&f�\T�A����_T
>"q}�7d�V�u*�5�Yv/x�:�RX`Z�l �SڍH咧U����f�vv�1\:T7Vwo~�� �O@��e�/���*ǹM���3ǚ�٬Kh��4]�`��Lv�-1�H��yMߦ3!���_m�~���[�$|�%��	��p�E�Y�b������Y���r�c�-v��|!m�,�v��t�;h|��|�����'��@,{�ٸ�0����/�hL�U<R�~�ȃM�i�-7��p�nl`(�AS��\����[���?H!ݺ�m�o4�����Xm'z�l�K��U���ԶV%����̀�_��R�5ʹۨʖy��[�P��0��#m��؛fv�:�80��/���_��jɑ-�s��$͙�T�ŘO��{r�r��_E8���{CO���zi��v��2Up�:.�e�Rm/)i�t'	xRU8s�΍�[��#�+{��k�p�}3܀�&����Ƞ��<��Fer���>T��}s�_C��)LQ�%1�lz��&�O��ET$�kB-�Z��R�s��v���5e9:5Z�s��ղD�0��Al!/s8��P��2)k)��{��G�E"���<'�nbFI�����'Tps	+k�ODV�TGؓ��mm�.b�^jQl�t_����`O��A��=2�uQA�C�;ժ��+ƥQ��g����d�pO�FnBղ����U!��U���P�p(���Jx��k���&������jB��qm�JJ�Z �/mB
�=�JtkS�:Mq�Wv<�>0�v'�����>A��q��{Ɯ=8~7�jM�Y�����DŔ(.Sr�Ƭw��J&���vz�'�I�ŗ��K�����P^��+��^3�����]����m�T�ǟ���,�ë�g�t��RN8�f�9|��� ���ӵ7����z�(!sY5���}%X���Zt��6��?{�Nq�C��ަ��y��4!��%	X���@Uj�(��\d�̞�@ǉ�YЇ<] �ʤ����&))�W��{�GX1}}��"�Y|�82+=9�#��Q��s�Rs7����B<W��kjH�<�G$˨>�f�F�Kx�p/KMT�4D���W�{��7���_vo�B�`a�P��r��_��d��ءv�f̍b��=ů����>- e_��/���۳��*�\r��젨�}�=T-����)YH$4	E�o��75��}����#�\=m�U[����x�L~�����h�`C�+`�k���;���XӓF(�d�ͦM�͟>��g�Fw��ۨ@�}���u��/N����3�,�oX��n��1P��	ɚ4��Ws�f��"�}8į;�L:p*��F���L����.��a 
4�5�~�u8�[�ҋ���/�08�'���L\���'��˴h?�4�u�@mf�!��&#�?��RS�Q�-1����&%���~E��>no�)kA������~���C�ߙ�N�ѱ�������=f|œ�bM��㻅�QI�@�ϑK� �m ��>!��V3�%��Z��4�_�e3
���^�Eyf�
���BE���"�������3� �Y@�D��E)���V�wʃ�IT���`X���}��B1����ԥb��y0�j�Y=���RPBp<f:�7ն��o}�X����Gd����#�������+��2.��&��v�w=
D́l#�����T)���*)�!�%�rs���ޜ��_
55��\)_�H���_Y���V�k�u�D��v:��W=�G�[>lC�������@��ڡ�OZԬ�Yzr�t���]� SG"�?G�kR���T�9t�R����r����䶯m�E�V���K@m�g�4�i0-�H󟜸���^X�$�
IK�dv��~�>3�b0�s#��}���Z3HCnFw�}d��	��i7��N���{�d%▔�p#t�"�T�� �mGQ�5�񡦁R��Y�3�[U��!g�E��+�QY�ʲ_�
�������.�!�>�К�fX}�5ď�����$���a����b�s�x�uC��,) �����=/%�7�q"w�?Gګ�Ǝԟ�/�D[U~o��ꖌ�o����#����?e��0�K�(�|~�*�#0��Ғ�tˠK���/�ntL}G��E�C���x��L"���U<��̾�"���J���Ra�-O%�Bi ���B�ۥ�'��rk>�uzG0��J3�ɠ�uSxG}z�L����'�[iW����o�t,�F�,[�v�{���q! �����K��.����R%{�n�1S�I!�.�O�X�v��<����7��@T�O�.@����8���Bw-�e#���P�E���|��?,�q��τzN�ho/r�R֨7H~uu�ȥr_R?�4�b�R�Vć��2�X.��'D��a�ߤ�=$��;-�E��J���ذ.��H �SF  �.}���S�U;�b%�v6CVl��]�	�� {䱘6	����t�ƽFy�j�=.�J�T�eJ�8l�d2�Q�М+���#��~�>�ugRJ�ͯ�ad	��<H��/����	 
 �ꅸRXt��Q���!�?U�w��Ò�MM��:]�y�'`�q�dY�LT��X��o|�-�L����=��.9�4��C����a���]�w H>��@�0��������|�z��خ�/�p�A��;:���|	��$qiGAS�'eO��;��m@ʨ�%����I�w�"�¥� ggں��,U���3u8�K\� �&�N~�(,d~HI�����F��F�~/�Fj�N:�'��S���f�.�8����B��SU�{c��
�y�q�y>�^���f����l���9u�Ap��g�̰�<QR����;��v�^$�644�ŇҬZ?��s�]�gņ�L��n�[���<�Bfv5�4[F6)��uȥ���}]2/xP%p[�C{�4���t�$�Ba��C�d�Y\���M �`xd"\���:9�ط<����X:�t�ż�CU(�m^�,�M@/�9_�!�%���o�q����aAZ�_�]�ʙ�P�/����(h?s2�'�,����f�h��`�1�8��l�^���E�n%]H��dK��nc	��OLq
~�:�۽TuN�yS�^e�^��6�@G��<K� �������gD}HU^��$�#É��L����V;�/tB�S�]T���jG�C�U�/sZ(�/�H7�|������D,�'����Mh�GA:�S��춫������|�>0���PG�% +�2t�?�&i_�Js�디���W.��z�V�=��9 ����u��L�v!���ܐ�o^ɡ�\J�R�m�3r�~�Fu=-�� ��2dK	+ ��K嘼q/���Y��Q���ѣ���7���-!G;$�N��d� �Tn��!$^"!��f:�N
P׎ɺzx�T�� ٶ��N䄩������1�����A#�c�����֩]����?If���JV��·��,�&?h�����vv6B�)��=��2:�K�޻ ��魏2 �P׻��y�-K�Z�@����5C�O� ����ڣI�a�4�����v}g��{�π`�[�J��7Ϩ���d#�Ę�y�$��kx b��6����y�|��?��,H�a���W��j�lճrf<��&�.4Ғ4���^�qW���>~�(�9@A��������w�uRz�25�3��16�����krc�Tܤ<���~.e"q��?r�5Ц7��u�i�X4A2]d�] �Ԫ�3���tRC]�U�y�C������$R���:\A/]����I�<>2��P �}E�������#r`'�&�z��^��-v����a$b\Jه�YsWC� o4�;��\ �!�S�|a2�D�E�Mmr+���+},�jl�g���ESP�0�\ *�����̈�8��a���B�B�.��X��g���r
�@�9��d�$��B`1� �;=��Ӑ}���`z����[01�sDOy���L�RXQjz��$<`8 ུl�)q�#o�HFj$���\eGu���u3��7�6pY���HeI ��F��#���ܙ,�=_�0^nW	�;�T���aI�%Q�HS-����t
���Lo�/�,ƑC\�ݎ4Nނ��D2�6ȑ�CzkE�w	�@�JW�/�Y]�t�H=*m v�bR�IE����~VZ��6���q<��r�s�_ >{�q(��^`1X&?/�B{��D�\�3j�����i� �O�]���4�����ǰ��g���h����ou�=��c�+��ܩ�4m������&��TK��ܖ�"�a���9�j���9j �� Q�k�U�k�)��$�W�a*���!Ҝٔ������Y?"$��6b9��bɝ$��B�˖��afvP�Qt�H�ˇb*�!qw�'{f�O�M/��2�qX�}�	�m x/��Ov����#M�k��w��r�p�R�;������TF���t�3�Gx��^L-�Ϝh��6:�ע�`ϻX�;bn�M�r�ghsؐ�s�޵wT3�E-D5�R���	��Lی N�h��!s���:W�@gQ!±֝`�=uwhi�@Kj}�6������S���i�ɳ�s�2@�Y0ɧ^��L���7���v�7ŏa������y�dt+l��C���W��w�Re�mf	�b�1����t?�� шyg�^_T��tn1_��~��4�O�a��'M�u�H`��|>��L#�� t������H�ĩ-�,��j�c�g�����6EH/�� +��_�<�}��R,��}6���'�v׬GzcH��:�X���3����tM�C��d$�̹�v�F>p�z�.-#���Ͽݾ=yAv\��Eȧ�V$
�����U�H#QG���dru����+��m��ǿ��?9�2�0X~�æ�?���8+�w&|kB5�䎄�[r"�m*X�*ͰKپ��/i>��F��R���j-��n��ޅC��a������2�G���xliB��Z�g*1��M�`'gI=���};Fb�����7�������u4��йL�%��
�a#��6
�*��7;��W�.U�H'����f|�to�q�"в�jϺUY&>ge%�n��䷲��1c��7��VB�{�]��ӄ��ӺI�
�2�v��m-m���:�X�������&�j�%��׼P����f&OE���������E��h��?Ѹ+a��2��W:k�\5�6�ƘҷXpN?o���?���@ƶ3~��y�ލ��w���J�����~3m&��jw�
���`Ӡ�ȱV�����w��Z����� D.nq�ςf+v]"�,J�;��[5�'`�[�CP�5�y����ϩ�b�X�J����QG�ź0)������"t"��܂�R^3��B�K�Sp���;�$�=�-�)%�fO+:��N�Z(�2�4YZ�q���OE�Z/�_ƿ��װ\�?gB�!�!#Ѿ�x@<��8e�{�%����pjgҋ�g��GN�z�����G���v~��;"�l����|�I��h��,F��\+i�R��K�0�����ë�+��O�:�#
~Jl!�
Bw�O�Nfzw��w�7|�zতhbu���i����G�
��i�lv��9eZ�w�F���0F~��^0o@QqGشrf�����+�{��*� �)�K�B^����1�:���P�~�7_"�>]�8;���3��{����2cd���Eɞ�\U��C�٢G��#�*�N�|�ppY
U�`�(�������)��`�X%]��d6}r��bg���?`4F��J�V0�0e=�v���ZW��dGQ�(r�.��r�H`Լ-�1b4e�<����*.j�g/(#��륋x.�V�y����z@Tt��U[���l��L���YXˏ4�h���
i^����Gu0�U�<>���ɴ�J�b�|�E����bp�5�B?�0"5�1eFd�2��=G\_&��Y�Bd�U���=�cǸ����BC.�Xs�C4c��X��qjS؁Kv��U%jݫ&�8��0��6�d��ٯX���;�;���s�LH�75��z���:�Jl�Fۍ�!�GM�NTsqt,������f�Ù�O�
��apc/;R*�Rh֒2�����&�++��+���3Ȝx�֛���TL������{��y�~�3��2X����u���| w��r8Q8�p@�d�E(��f�'�#�m�X�����u�f��Q=� �r.�ۄ�Sh�)!�KT��iOu����mQ6�������p��c�{{)���&�m��>��1s��𫈖�Gtd� l;+�f���y�3�=�nL��^�����I�h�g�_�&����yj�B��C�� q��6�������ؑ���AcyE8�o�@.��)ھ��A�j����Wz>	�z�Fs�zaз����i%����~e?��E�� .e�Y����
����y8���XP��2X����80���e��L�{P��O\��A�����.�Lh�8��Q�[� ��:�)�+{����4np��t��x�W�hv��T��w�A�w?��B�/m�V�f��'ޟ�j�ʆ�K�u���\G��u�mZS���+ю����`��(Q�j�~����䍤+	Y[C�@v���q8S�`2�+0��r'[��ٕ�'�s���,����Z��n��Fr���oҺ�I�E���eJ�����&4�Y�xT����a���53����]�2Eg�����K�q{���Ų��c�?+/��U���{��s�l�9Z+�"�1��҉qn�v;oN=7�k��nh�S+*AB�fM0g|�+2�,m2��L���Ă}�3�o��@n?I�ڕE���ퟻ1.7�[C:v�0=rd4�	rۦ���ZBOob�|�3��Ѥ���?�YC�zv�x�>�F�IY�w|6����ɣ��/�j�F�WkǴ2�,R��1y���Ǫ���Г��~ON�sJb�pk���9uFX�߻���>�M��Tljؐ/�r����]���;�fu�sF!��9ɷ<S`�LJ W�Tf�+�&�k�{f-�\�j^�3�̟C8x�M)o��#�:�IU��������?�y��ѐ�>�*�z^h�����[Y�7�9ໃ�k�S�J#�ǐ�h�m���ho����
ے�1�*����
������ ��2�F��C�-��0z��.F��a9&�O�����3�MK���U��襒���S�2?�b�����򷍑$$� X� �
�4''�!jV�c�A"�r7O�2���j�·_2g��Js���Ɨ���) ��$�Se�}�vvμ���	����au9��2��r��3N�Q;�R<E_w�U�N��[���t��f�Ռ��T���x��;5[lz�̀r�L�[R��p���7���Mu�B�j��_�"ɣT������h���ebcӄ0.��bywN���?�lx���>�����>;ÑC�`�3Y�������O���Z:��b�3��8ɼ-�F.1���(*e)���n�w檯��M�Ii��\O�Sh�ێp�f N#�:{[�nG"x8ؕ2!��y5H��'���G���J_W��)l