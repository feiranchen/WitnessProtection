��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]Q�F��t�K�j�;�:i�)8	�7�n�8e�}�*�6���ծ�p�	'(�Rt�Y%�"�6x�]o��ݤЌe�V�l���i#����/Ks�c��<��J��ś@$�w��z�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i �DH�[��U -�����1�)�+q(FW�#;��Ϣ���g���l�<�a�K�Y�^�y�Ijĸ*����6;�3e��@_g6�Ω~a�iI�-���Oy�Fׂ�����Zj�S��p>�J�/�Zt8���y�!NX$ .2@x�5�m�<9�M��N�H�3c��U�y���o�ͽ�s����`T=�U?�P|�Ѹd|wH���[�o��TtB��p�;,=R7�H
��+ϵ�Q�,&@���q�Ѡ�- �_��2]d��pEc���{}����;�X������}�,�۳�L�Dtu�[,�D�DaV��$;G��K�w<c�,��X{IG�;�׳���7��էQ�7+�@�A�
d&t������Z��SP9��%趢����I��3�� /�A�]��?lJ�ݠ�Tk���s�(�v�O���GJ��rV����Ś��qG
�BN�f��w-*\�LtB`�>_,�����C���E��u�E ��D���H��IY%Qs���Og�L��g'��p��I��=L�/[D%]����\��%������ ���]r!M;9V,8�x�ݰ1�7{g��1��Ŭ:��j��M��Y�����:���+�О��@y���P/�^�n���^�NOD��S�|<�ջ��ۜѫa$s��L����{D����*«u�}C����Y��~��M��dݷ��:2�T
��}n)m�7��q��=�b�OӒ��b
ot�.@̙��)�y�*�0+��dʮ�]�?�i*LY[����掂C��t:��sC�^Yߣ��C������Ȭy��%3��z�A�L�A�D���@���^��OWz<��
�]G����[�U�+c��4��b�RZ�Pb�]͉Kj�4�5��S�E���\I�O���"R˂��՛Mu� mH�'s���4��?Q6,�?X�i�*q@��;`�H��0
�PY�-%Md+�^[���xX�&��Z��YN $�yܕ`��$L�����z��9�u =u�хw�֥W���@�.N���Ҹ*m���p�Ԣh�off�aSݾf�o�ظ����A��v�3��+���>�K�3Rey�	��{��[��U��
�z�03��}�j�d��y�T���K�X"JY`q&uz�%��*�0�Q�jL�/�t��]����uw��d�.Vo7d�b���`N�f!����rZd���1f��������mj=\ǟ�� ~���Dy�Q@�!�I���V �+TCŐ��)Q'��)��˶�pImb`�/��L�? �[�?�&s}z�^�e~&`J��5��&ɐ!	DŴ��D�8���0�5�	�#�}?ْ��m&������l�nӦ[��3��3���̲w�ܓ���3����<9��<�Fל�����Tw�K��~	7y���8˫�oܬ��l��1��ۣ)����p�S`D����r��})ڏ�N�p5|���^lZ��g���j�:�C]\�u��N�X�.�ry�U�B���Q������$8�W�eC�&���F��ё^M[��l��O�V�`rjJ��ƊC��߿z����?U����9�Q^F�^X��{P�U�P�Rj����1�M�b�]���32���$�6T6�E�[�T��o�ֳ�����Q��g{��=�6�ގ�:�N�y-�y�磨���͎�r�\���W����#��Q�4�K�}+���)^m�9"_M��лO�.��aO�-;5W��X��̫{���G� �E��>i)Y^Ď�ʥ`y̥?��H,Ӗ�`�~�{ȃƠ����g����Z�/-��g%-���W^v�R�9�{3���E�]��bP�>���-	��s�T�AS�����Q�nD`����N*��.��\aiu�1�T�� ��,bE�Xj{.���rC�s�(�X��V������u�����3�u.���\� f�9&�?��%T�y�j�_�l�`��"U�[��yc*=�vsƌ��˸���Ջ��<P�~u��Ǎ��N��X�]�����,Pg��W"��^�����z�5��!|���{U*�����?~����͵[���~t���Hݜ�M�9�uS��H���R7������z�՜��X,t���`v��x�X:=���5�'v�Ϣ�x�H>O9}е���
f��w�PP���$�2�$���/8��~�U��?�kF'@�w�y`�����G�<tuO�7���2>���3���˺[����uYPR�I/ȝVK8�8}��#�8�a�d�YF:����FM�/���3#�j4$媅�-j$�t=7���Aa�h4D4�MI	�
��i�����0���A�6� �+�eXt��?4���� �Is|�ėo�!uII��k����(��n�1�=��f���i�iF*������ɰ7���g�C�-���`6����EYCWǒ�@�ӬU>$�V�'9r(�t�N/��F�
/�;�W3��[~6�ω�v8̸�*X��k�!��PEo*�ͦ�y�O
��^lR���� t��Jd��Lw|��oA��O<�۾�V
���4��;�F\̇�#�y�+H��������1+�T��u��9!N!& �����j���
���n��S�N��Z�3�%|������o�����p���MӔ_X��Ri�G��=W#N�IeU�KR�
�Q��-r��Ud�#޵1�7vJ?��o)�= �.:R�p�Q������o�d�t�o!ƦE<b�[��2���hB1����ɹ�ʶ�~ܧF���b�f�ن�{���.����ˢѿ�� �h}٠S>�ܬB�j��Bb�V͙~����q�z{mG�=�!�d��y�n���op܌�����b��9$�>�%y�������v[ˁXX��d`T�ԧj�ӺȁG����s)z��D3#�2�����Jqڱ\%�H���(6�D�z[��!y���/@~}!r4��Q�͠y󨋋Ա)�r����u|��z����B��Q�2|����:;�!L�+x�K��b�